(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h8d9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire3;
  input wire signed [(4'hf):(1'h0)] wire2;
  input wire signed [(4'ha):(1'h0)] wire1;
  input wire signed [(3'h6):(1'h0)] wire0;
  wire signed [(3'h6):(1'h0)] wire2310;
  wire [(3'h6):(1'h0)] wire2292;
  wire [(4'he):(1'h0)] wire2291;
  wire [(4'h9):(1'h0)] wire2234;
  wire [(3'h4):(1'h0)] wire2103;
  wire [(3'h7):(1'h0)] wire2101;
  wire signed [(4'h9):(1'h0)] wire2284;
  wire [(4'hd):(1'h0)] wire2287;
  wire signed [(3'h7):(1'h0)] wire2289;
  reg signed [(2'h2):(1'h0)] reg2307 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2305 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2301 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2300 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2299 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2297 = (1'h0);
  reg [(4'hc):(1'h0)] reg2295 = (1'h0);
  reg [(3'h5):(1'h0)] reg2293 = (1'h0);
  reg [(2'h2):(1'h0)] reg2233 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2228 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2226 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2225 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2220 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2217 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2216 = (1'h0);
  reg [(3'h5):(1'h0)] reg2214 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2211 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2208 = (1'h0);
  reg [(4'hb):(1'h0)] reg2205 = (1'h0);
  reg [(4'h9):(1'h0)] reg2203 = (1'h0);
  reg [(2'h3):(1'h0)] reg2199 = (1'h0);
  reg [(4'h8):(1'h0)] reg2194 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2187 = (1'h0);
  reg [(3'h6):(1'h0)] reg2183 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2182 = (1'h0);
  reg [(3'h4):(1'h0)] reg2181 = (1'h0);
  reg [(4'he):(1'h0)] reg2179 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2176 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2172 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2158 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2168 = (1'h0);
  reg [(4'hd):(1'h0)] reg2167 = (1'h0);
  reg [(4'hb):(1'h0)] reg2164 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2161 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2160 = (1'h0);
  reg [(4'hd):(1'h0)] reg2159 = (1'h0);
  reg [(4'hd):(1'h0)] reg2136 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2131 = (1'h0);
  reg [(3'h6):(1'h0)] reg2150 = (1'h0);
  reg [(4'ha):(1'h0)] reg2145 = (1'h0);
  reg [(4'ha):(1'h0)] reg2138 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2137 = (1'h0);
  reg [(4'hd):(1'h0)] reg2133 = (1'h0);
  reg [(4'hc):(1'h0)] reg2132 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2126 = (1'h0);
  reg [(4'hb):(1'h0)] reg2124 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2122 = (1'h0);
  reg [(2'h3):(1'h0)] reg2118 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2116 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2115 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2114 = (1'h0);
  reg [(4'h9):(1'h0)] reg2109 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2105 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2107 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2104 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2237 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2241 = (1'h0);
  reg [(4'h9):(1'h0)] reg2243 = (1'h0);
  reg [(4'ha):(1'h0)] reg2247 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2253 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2256 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2258 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2259 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2261 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2263 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2264 = (1'h0);
  reg [(4'ha):(1'h0)] reg2269 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2270 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2271 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2272 = (1'h0);
  reg [(4'hc):(1'h0)] reg2277 = (1'h0);
  reg [(4'ha):(1'h0)] reg2285 = (1'h0);
  reg [(4'hd):(1'h0)] reg2309 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2308 = (1'h0);
  reg [(3'h4):(1'h0)] reg2306 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2299 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2304 = (1'h0);
  reg [(4'hc):(1'h0)] reg2303 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2302 = (1'h0);
  reg [(2'h3):(1'h0)] reg2298 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2294 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2293 = (1'h0);
  reg [(3'h6):(1'h0)] reg2296 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2294 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2286 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2283 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2267 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2265 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2264 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2282 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2281 = (1'h0);
  reg [(4'hd):(1'h0)] reg2280 = (1'h0);
  reg [(4'h9):(1'h0)] reg2279 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2278 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2274 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2273 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2269 = (1'h0);
  reg [(3'h4):(1'h0)] reg2268 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2278 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2276 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2275 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2274 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2273 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2268 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2267 = (1'h0);
  reg [(4'hd):(1'h0)] reg2266 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2265 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2262 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2260 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2256 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2251 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2250 = (1'h0);
  reg [(4'ha):(1'h0)] reg2249 = (1'h0);
  reg [(3'h6):(1'h0)] reg2248 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2245 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2242 = (1'h0);
  reg [(4'he):(1'h0)] forvar2240 = (1'h0);
  reg [(4'he):(1'h0)] reg2257 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2255 = (1'h0);
  reg [(4'hf):(1'h0)] reg2254 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2252 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2251 = (1'h0);
  reg [(3'h5):(1'h0)] reg2250 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2249 = (1'h0);
  reg [(4'he):(1'h0)] forvar2248 = (1'h0);
  reg [(3'h6):(1'h0)] reg2246 = (1'h0);
  reg [(4'hd):(1'h0)] reg2245 = (1'h0);
  reg [(4'h8):(1'h0)] reg2244 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2242 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2240 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2239 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2238 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2236 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2232 = (1'h0);
  reg [(4'hc):(1'h0)] reg2231 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2230 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2229 = (1'h0);
  reg [(4'hf):(1'h0)] reg2227 = (1'h0);
  reg [(4'hd):(1'h0)] reg2224 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2223 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2222 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2221 = (1'h0);
  reg [(5'h10):(1'h0)] reg2219 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2218 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2215 = (1'h0);
  reg [(4'hd):(1'h0)] reg2213 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2212 = (1'h0);
  reg [(3'h6):(1'h0)] reg2212 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2210 = (1'h0);
  reg [(4'hb):(1'h0)] reg2209 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2207 = (1'h0);
  reg [(2'h2):(1'h0)] reg2206 = (1'h0);
  reg [(4'h9):(1'h0)] reg2204 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2202 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2201 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2200 = (1'h0);
  reg [(4'hd):(1'h0)] reg2198 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2197 = (1'h0);
  reg [(4'hd):(1'h0)] reg2196 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2195 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2193 = (1'h0);
  reg [(5'h10):(1'h0)] reg2192 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2191 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2190 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2189 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2188 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2180 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2175 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2174 = (1'h0);
  reg [(3'h5):(1'h0)] reg2186 = (1'h0);
  reg [(3'h5):(1'h0)] reg2185 = (1'h0);
  reg [(4'hb):(1'h0)] reg2184 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2180 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2178 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2177 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2175 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2174 = (1'h0);
  reg [(3'h4):(1'h0)] reg2173 = (1'h0);
  reg [(4'hd):(1'h0)] reg2171 = (1'h0);
  reg [(2'h2):(1'h0)] reg2170 = (1'h0);
  reg [(4'he):(1'h0)] reg2169 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2166 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2163 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2159 = (1'h0);
  reg [(2'h3):(1'h0)] reg2156 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2155 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2153 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2166 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2165 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2163 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2162 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2158 = (1'h0);
  reg [(2'h3):(1'h0)] reg2157 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2156 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2155 = (1'h0);
  reg [(3'h5):(1'h0)] reg2154 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2153 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2152 = (1'h0);
  reg [(4'h9):(1'h0)] reg2148 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2145 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2137 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2121 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2119 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2108 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2104 = (1'h0);
  reg [(3'h5):(1'h0)] reg2151 = (1'h0);
  reg [(3'h7):(1'h0)] reg2149 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2148 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2147 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2146 = (1'h0);
  reg [(2'h3):(1'h0)] reg2144 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2143 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2142 = (1'h0);
  reg [(2'h2):(1'h0)] reg2141 = (1'h0);
  reg [(4'hd):(1'h0)] reg2140 = (1'h0);
  reg [(4'hf):(1'h0)] reg2139 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2136 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2135 = (1'h0);
  reg [(4'h9):(1'h0)] reg2134 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2131 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2130 = (1'h0);
  reg [(4'hc):(1'h0)] reg2129 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2128 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2127 = (1'h0);
  reg [(3'h6):(1'h0)] reg2125 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2123 = (1'h0);
  reg [(4'hc):(1'h0)] reg2121 = (1'h0);
  reg [(3'h5):(1'h0)] reg2120 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2119 = (1'h0);
  reg [(4'hb):(1'h0)] reg2117 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2107 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2113 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2112 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2111 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2110 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2109 = (1'h0);
  reg [(4'h8):(1'h0)] reg2108 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2106 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2105 = (1'h0);
  assign y = {wire2289,
                 reg2307,
                 reg2301,
                 reg2233,
                 reg2216,
                 reg2211,
                 reg2187,
                 reg2183,
                 reg2176,
                 reg2172,
                 reg2161,
                 reg2150,
                 reg2145,
                 reg2133,
                 reg2114,
                 reg2241,
                 reg2259,
                 reg2261,
                 reg2264,
                 reg2304,
                 reg2302,
                 reg2298,
                 reg2294,
                 forvar2293,
                 forvar2294,
                 reg2286,
                 reg2283,
                 reg2265,
                 forvar2264,
                 forvar2278,
                 reg2275,
                 forvar2273,
                 forvar2265,
                 forvar2251,
                 forvar2250,
                 reg2249,
                 reg2242,
                 reg2254,
                 forvar2249,
                 forvar2248,
                 reg2245,
                 reg2239,
                 reg2238,
                 reg2236,
                 reg2232,
                 reg2231,
                 reg2222,
                 forvar2218,
                 forvar2215,
                 reg2212,
                 reg2204,
                 reg2202,
                 forvar2200,
                 forvar2197,
                 reg2192,
                 forvar2189,
                 reg2188,
                 reg2185,
                 reg2184,
                 forvar2180,
                 forvar2174,
                 reg2171,
                 forvar2159,
                 forvar2166,
                 reg2163,
                 forvar2158,
                 reg2157,
                 forvar2155,
                 reg2119,
                 forvar2148,
                 forvar2143,
                 reg2142,
                 reg2134,
                 reg2130,
                 reg2128,
                 reg2127,
                 reg2125,
                 reg2123,
                 reg2121,
                 reg2120,
                 forvar2119,
                 reg2113,
                 reg2112,
                 reg2111,
                 reg2106,
                 (1'h0)};
  module4 #() modinst2102 (.wire5(wire0), .clk(clk), .y(wire2101), .wire7(wire3), .wire6(wire2), .wire8(wire1));
  assign wire2103 = "5A9aDaLoub4J";
  always
    @(posedge clk) begin
      if ($signed((8'ha2)))
        begin
          reg2104 <= $unsigned($signed(wire0));
          if ($signed(wire1))
            begin
              if ((+(8'hb8)))
                begin
                  for (forvar2105 = (1'h0); (forvar2105 < (1'h1)); forvar2105 = (forvar2105 + (1'h1)))
                    begin
                      reg2106 = {$signed($unsigned("BAVg"))};
                      reg2107 <= $unsigned($unsigned(((forvar2105 >= wire1) == (wire2101 >>> wire2103))));
                      reg2108 = $unsigned(wire3[(5'h10):(4'hc)]);
                    end
                  for (forvar2109 = (1'h0); (forvar2109 < (1'h0)); forvar2109 = (forvar2109 + (1'h1)))
                    begin
                      reg2110 = {$unsigned(wire2101[(2'h2):(1'h0)])};
                      reg2111 = reg2108;
                      reg2112 = (reg2110[(1'h1):(1'h0)] ?
                          {$unsigned({(8'hb3)})} : ("8IU9F" ?
                              wire2101 : wire2101));
                    end
                  reg2113 = $signed("lzrAbgHS8s");
                end
              else
                begin
                  if (reg2110)
                    begin
                      reg2105 <= (wire0[(2'h3):(1'h1)] ?
                          $unsigned($unsigned($signed(reg2108))) : (&reg2107));
                      reg2106 = ($unsigned(reg2105[(3'h5):(1'h1)]) ?
                          {"6LTSWCuYL"} : "3UkNQn52r");
                    end
                  else
                    begin
                      reg2105 <= {$unsigned(((wire0 >> reg2113) >> wire2))};
                    end
                  for (forvar2107 = (1'h0); (forvar2107 < (1'h0)); forvar2107 = (forvar2107 + (1'h1)))
                    begin
                      reg2109 <= ($unsigned(($unsigned(wire2103) <<< (^~wire1))) & ($unsigned(reg2106[(3'h6):(3'h5)]) ^~ $unsigned(reg2106[(3'h7):(3'h5)])));
                      reg2110 = ($unsigned($unsigned($signed(reg2107))) + $unsigned(((+wire1) >= (|wire2101))));
                      reg2111 = ((+wire3) ? reg2104 : reg2109);
                    end
                  if (($signed((reg2111[(3'h4):(2'h2)] ^~ $unsigned(wire1))) >> reg2113[(2'h3):(1'h0)]))
                    begin
                      reg2114 <= $signed("SQeVC7s");
                      reg2115 <= reg2106[(1'h1):(1'h0)];
                      reg2116 <= reg2113;
                    end
                  else
                    begin
                      reg2112 = reg2109[(4'h8):(3'h7)];
                      reg2114 <= (({((8'hac) ? forvar2105 : wire2)} ?
                              reg2105[(2'h2):(1'h1)] : reg2114) ?
                          $signed($unsigned({wire2103})) : ((!(wire2 ~^ forvar2109)) ?
                              $unsigned(reg2110) : {{forvar2109}}));
                      reg2115 <= (8'hb0);
                      reg2117 = $unsigned($signed(reg2110[(2'h2):(1'h1)]));
                    end
                end
              reg2118 <= (&reg2116[(3'h5):(2'h2)]);
              for (forvar2119 = (1'h0); (forvar2119 < (2'h2)); forvar2119 = (forvar2119 + (1'h1)))
                begin
                  if (reg2116)
                    begin
                      reg2120 = (reg2117 ?
                          ({(reg2108 ?
                                  reg2115 : reg2109)} * $unsigned((reg2118 ?
                              reg2108 : reg2114))) : reg2112[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg2120 = $unsigned({"bkIb1iMAeD"});
                      reg2121 = reg2120;
                      reg2122 <= $signed(($signed("6Z") ?
                          "5dWCpll5C" : ($signed(reg2112) == $unsigned(forvar2109))));
                    end
                  if (({(-wire0)} - $unsigned(($unsigned((8'ha3)) >>> (reg2106 < (8'haa))))))
                    begin
                      reg2123 = {$unsigned(("WoUXpMW5yUJ" ?
                              (reg2107 ?
                                  forvar2105 : reg2120) : $signed(reg2116)))};
                      reg2124 <= $signed((~|$signed({wire2})));
                      reg2125 = ("" ?
                          forvar2107[(2'h2):(2'h2)] : ({reg2112[(4'ha):(2'h3)]} >= (&{wire3})));
                    end
                  else
                    begin
                      reg2124 <= wire0;
                      reg2126 <= reg2112;
                      reg2127 = (!{{$signed((8'h9c))}});
                      reg2128 = reg2125;
                    end
                  reg2129 = reg2125;
                end
              reg2130 = wire2103[(2'h3):(2'h2)];
            end
          else
            begin
              reg2106 = ((^~$unsigned({(8'haa)})) == reg2128);
              reg2108 = "pQVxdgz1SamT";
            end
          for (forvar2131 = (1'h0); (forvar2131 < (1'h1)); forvar2131 = (forvar2131 + (1'h1)))
            begin
              reg2132 <= (8'ha7);
              reg2133 <= ((|(reg2128 ? wire1 : (|forvar2119))) >>> (8'h9d));
              reg2134 = ((^reg2127) ^ reg2133[(2'h2):(2'h2)]);
              for (forvar2135 = (1'h0); (forvar2135 < (2'h2)); forvar2135 = (forvar2135 + (1'h1)))
                begin
                  for (forvar2136 = (1'h0); (forvar2136 < (2'h3)); forvar2136 = (forvar2136 + (1'h1)))
                    begin
                      reg2137 <= $signed({(~&$signed(reg2110))});
                    end
                  if (forvar2135[(1'h0):(1'h0)])
                    begin
                      reg2138 <= (8'ha1);
                    end
                  else
                    begin
                      reg2139 = (($unsigned($unsigned(forvar2107)) > ($unsigned(reg2130) ?
                              (reg2108 ? reg2112 : wire0) : {reg2129})) ?
                          (wire0 ?
                              reg2114[(1'h1):(1'h0)] : ($unsigned(forvar2109) ?
                                  $unsigned(wire2101) : (forvar2107 == forvar2135))) : $unsigned(forvar2105));
                      reg2140 = ($signed($signed(reg2109)) ~^ $signed(($unsigned(forvar2119) <= reg2128[(4'hb):(3'h5)])));
                      reg2141 = (&reg2106[(2'h3):(2'h3)]);
                      reg2142 = $signed({$signed((wire2103 ?
                              reg2137 : (8'ha8)))});
                    end
                  for (forvar2143 = (1'h0); (forvar2143 < (2'h2)); forvar2143 = (forvar2143 + (1'h1)))
                    begin
                      reg2144 = ((reg2129 ?
                          ($unsigned(forvar2107) ?
                              (!(8'had)) : (!reg2141)) : {(~^reg2122)}) - $signed(reg2115[(4'he):(4'h8)]));
                      reg2145 <= reg2114;
                      reg2146 = (forvar2143 ?
                          ((forvar2131 ?
                              (~^reg2140) : forvar2109) > $signed((reg2130 > reg2111))) : "MDhN");
                      reg2147 = (^$unsigned(($unsigned(reg2117) ?
                          $unsigned(reg2115) : reg2144)));
                    end
                  for (forvar2148 = (1'h0); (forvar2148 < (2'h3)); forvar2148 = (forvar2148 + (1'h1)))
                    begin
                      reg2149 = reg2107[(1'h1):(1'h1)];
                      reg2150 <= $signed($signed(reg2141[(1'h1):(1'h1)]));
                      reg2151 = $unsigned({((reg2118 ? reg2111 : (8'hb1)) ?
                              $unsigned(reg2107) : $unsigned(reg2108))});
                    end
                end
            end
        end
      else
        begin
          for (forvar2104 = (1'h0); (forvar2104 < (1'h1)); forvar2104 = (forvar2104 + (1'h1)))
            begin
              for (forvar2105 = (1'h0); (forvar2105 < (1'h1)); forvar2105 = (forvar2105 + (1'h1)))
                begin
                  reg2107 <= "HIM3m";
                  for (forvar2108 = (1'h0); (forvar2108 < (2'h3)); forvar2108 = (forvar2108 + (1'h1)))
                    begin
                      reg2110 = $unsigned(($signed($signed((8'haf))) ?
                          ({reg2111} | (reg2117 ?
                              reg2144 : forvar2135)) : reg2132[(1'h1):(1'h0)]));
                      reg2114 <= $unsigned($unsigned((8'ha9)));
                    end
                  reg2117 = reg2127[(4'h8):(1'h0)];
                  if ("JHbLV4")
                    begin
                      reg2118 <= reg2146;
                      reg2119 = (reg2132 <<< (((reg2129 ^ forvar2136) || (wire0 && (8'hb5))) <<< reg2124[(4'ha):(3'h5)]));
                      reg2120 = $signed((reg2129 ?
                          $signed(forvar2119) : reg2122[(5'h10):(3'h4)]));
                    end
                  else
                    begin
                      reg2119 = $unsigned($signed((forvar2108 == forvar2135[(3'h4):(2'h2)])));
                    end
                end
              if (reg2125)
                begin
                  for (forvar2121 = (1'h0); (forvar2121 < (2'h3)); forvar2121 = (forvar2121 + (1'h1)))
                    begin
                      reg2122 <= {$unsigned($signed("eSKvisWakGO3"))};
                      reg2123 = $signed((((~|reg2129) || ((8'ha1) < reg2150)) ^~ ((~(8'hb1)) << "kZiWXmmgg")));
                    end
                end
              else
                begin
                  reg2121 = $signed((~((forvar2136 ? reg2130 : forvar2148) ?
                      (-(8'ha1)) : forvar2109[(3'h4):(3'h4)])));
                end
              if ($signed({$signed(reg2119[(3'h5):(2'h3)])}))
                begin
                  reg2125 = {(((reg2104 * forvar2108) ?
                              $signed(reg2109) : $unsigned(forvar2121)) ?
                          ($signed(reg2107) - reg2117) : wire3[(3'h4):(3'h4)])};
                end
              else
                begin
                  if ($unsigned(reg2150))
                    begin
                      reg2124 <= (8'ha5);
                      reg2125 = $signed(((-(reg2150 ?
                          reg2110 : reg2123)) || $unsigned((reg2139 && wire2101))));
                    end
                  else
                    begin
                      reg2125 = reg2144;
                      reg2126 <= reg2151[(3'h5):(2'h2)];
                      reg2131 <= wire2103;
                    end
                  reg2134 = (({(reg2145 ? reg2120 : wire0)} ^~ reg2140) ?
                      reg2115[(4'hd):(4'hc)] : (reg2139 ^~ {{reg2112}}));
                end
              for (forvar2135 = (1'h0); (forvar2135 < (2'h2)); forvar2135 = (forvar2135 + (1'h1)))
                begin
                  reg2136 <= forvar2136[(3'h4):(2'h2)];
                  for (forvar2137 = (1'h0); (forvar2137 < (1'h1)); forvar2137 = (forvar2137 + (1'h1)))
                    begin
                      reg2139 = (reg2147[(2'h2):(2'h2)] == $unsigned(((!(8'hac)) || (^~forvar2136))));
                      reg2140 = reg2146[(4'h9):(3'h7)];
                      reg2141 = ($unsigned($signed($unsigned(forvar2121))) ?
                          (^($unsigned(forvar2105) * (8'hb1))) : $unsigned($unsigned((&reg2108))));
                      reg2142 = $signed((($unsigned(reg2131) ?
                              (-reg2149) : reg2118) ?
                          $unsigned(forvar2108) : ($unsigned(reg2147) << $unsigned(reg2125))));
                    end
                  for (forvar2143 = (1'h0); (forvar2143 < (1'h1)); forvar2143 = (forvar2143 + (1'h1)))
                    begin
                      reg2144 = ((8'hb6) != reg2136[(3'h4):(1'h1)]);
                    end
                  for (forvar2145 = (1'h0); (forvar2145 < (2'h3)); forvar2145 = (forvar2145 + (1'h1)))
                    begin
                      reg2146 = {reg2128[(3'h4):(2'h3)]};
                      reg2147 = $signed(reg2140);
                    end
                end
            end
          reg2148 = forvar2119;
          reg2150 <= {(~&(|(reg2126 ? reg2147 : (8'ha9))))};
        end
      for (forvar2152 = (1'h0); (forvar2152 < (1'h1)); forvar2152 = (forvar2152 + (1'h1)))
        begin
          if (wire2[(4'h9):(1'h0)])
            begin
              reg2153 = $signed(reg2147);
              reg2154 = reg2114[(2'h2):(1'h0)];
              for (forvar2155 = (1'h0); (forvar2155 < (2'h3)); forvar2155 = (forvar2155 + (1'h1)))
                begin
                  for (forvar2156 = (1'h0); (forvar2156 < (2'h3)); forvar2156 = (forvar2156 + (1'h1)))
                    begin
                      reg2157 = reg2129[(3'h7):(3'h4)];
                    end
                  for (forvar2158 = (1'h0); (forvar2158 < (1'h1)); forvar2158 = (forvar2158 + (1'h1)))
                    begin
                      reg2159 <= $signed((!$unsigned(reg2117)));
                      reg2160 <= reg2123;
                    end
                  if ({(($signed(reg2150) ?
                              $unsigned(reg2137) : (forvar2131 >>> reg2110)) ?
                          $unsigned($signed(reg2126)) : forvar2104)})
                    begin
                      reg2161 <= $signed(reg2133[(4'h8):(1'h0)]);
                      reg2162 = $unsigned(reg2136);
                    end
                  else
                    begin
                      reg2162 = $unsigned(($signed($signed(forvar2155)) ?
                          ($signed((8'hb7)) >> reg2133[(2'h2):(1'h1)]) : $signed($unsigned(forvar2107))));
                      reg2163 = reg2138;
                      reg2164 <= ((~^($unsigned(forvar2136) ?
                          (^~reg2105) : {reg2110})) || ($signed($signed(reg2160)) ~^ reg2153[(3'h4):(3'h4)]));
                    end
                  reg2165 = "4UrpVG5ZmREwVV";
                end
              for (forvar2166 = (1'h0); (forvar2166 < (2'h3)); forvar2166 = (forvar2166 + (1'h1)))
                begin
                  reg2167 <= forvar2107;
                  reg2168 <= {$signed("eo2")};
                end
            end
          else
            begin
              for (forvar2153 = (1'h0); (forvar2153 < (2'h2)); forvar2153 = (forvar2153 + (1'h1)))
                begin
                  reg2154 = "ZfMXn6S2R";
                  reg2155 = reg2138;
                  reg2156 = $signed((~&"YUOmeegJ"));
                end
              reg2157 = $unsigned($signed("Ahd9frcVSZ5y"));
              reg2158 <= reg2108[(3'h7):(3'h7)];
              for (forvar2159 = (1'h0); (forvar2159 < (1'h0)); forvar2159 = (forvar2159 + (1'h1)))
                begin
                  reg2162 = ((reg2160 > {(8'hb0)}) != reg2131);
                  for (forvar2163 = (1'h0); (forvar2163 < (2'h2)); forvar2163 = (forvar2163 + (1'h1)))
                    begin
                      reg2165 = {reg2155[(2'h2):(1'h0)]};
                      reg2166 = $signed(("aCtx7185GnPBz" ?
                          $unsigned({reg2167}) : $unsigned($unsigned(reg2125))));
                      reg2169 = {$unsigned((~(8'ha4)))};
                    end
                  if ("kBLQU")
                    begin
                      reg2170 = (reg2142[(3'h5):(1'h1)] && $unsigned(("lA6gTwp" > {(8'hb6)})));
                      reg2171 = reg2133;
                      reg2172 <= reg2147[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg2170 = "atiH9QKKb47";
                      reg2172 <= $unsigned(({forvar2121} ?
                          forvar2155[(1'h1):(1'h1)] : ("lwU3" ?
                              (forvar2156 ^ reg2142) : $signed(wire0))));
                      reg2173 = (forvar2152 ?
                          {$signed((reg2149 && reg2145))} : $signed(($signed(reg2121) ?
                              (reg2114 <= (8'h9d)) : reg2126[(4'hc):(2'h3)])));
                    end
                end
            end
          if ($signed("T"))
            begin
              for (forvar2174 = (1'h0); (forvar2174 < (2'h2)); forvar2174 = (forvar2174 + (1'h1)))
                begin
                  if ($unsigned((wire3[(4'h9):(3'h5)] ?
                      $unsigned($signed(reg2123)) : forvar2152[(1'h0):(1'h0)])))
                    begin
                      reg2175 = ($signed((reg2145[(4'ha):(1'h0)] ?
                          reg2165 : $unsigned((8'had)))) != (^((forvar2143 | reg2137) ?
                          {reg2146} : reg2127[(4'h9):(4'h8)])));
                      reg2176 <= {$signed((|(reg2128 != reg2156)))};
                      reg2177 = $signed($signed(reg2133));
                    end
                  else
                    begin
                      reg2176 <= (8'hb0);
                      reg2177 = (forvar2104 >>> wire0);
                      reg2178 = reg2157[(2'h2):(1'h1)];
                    end
                end
              reg2179 <= (^~$signed(("yctCzvgndc" ?
                  ((8'hb4) == reg2175) : ((8'hb2) - reg2130))));
              for (forvar2180 = (1'h0); (forvar2180 < (1'h1)); forvar2180 = (forvar2180 + (1'h1)))
                begin
                  reg2181 <= {(^reg2139[(4'hc):(1'h1)])};
                  if ($signed(reg2147))
                    begin
                      reg2182 <= reg2141[(1'h1):(1'h1)];
                      reg2183 <= $unsigned((($unsigned((8'h9d)) == (-reg2112)) ?
                          (reg2158 << {reg2164}) : (~^$unsigned(reg2140))));
                      reg2184 = (8'hba);
                      reg2185 = (reg2160[(4'h9):(3'h5)] ?
                          ({$signed(reg2124)} ?
                              (^((8'ha1) << reg2146)) : (~&(^reg2164))) : reg2128);
                    end
                  else
                    begin
                      reg2184 = (^(^reg2111[(4'he):(2'h2)]));
                      reg2185 = $unsigned($unsigned((~|reg2122)));
                      reg2186 = (+reg2124);
                    end
                end
            end
          else
            begin
              reg2174 = {(-$signed((forvar2108 ? forvar2156 : reg2138)))};
              for (forvar2175 = (1'h0); (forvar2175 < (1'h1)); forvar2175 = (forvar2175 + (1'h1)))
                begin
                  if (reg2106[(3'h7):(3'h7)])
                    begin
                      reg2176 <= (+{(!$signed(reg2183))});
                      reg2177 = (&"3goZKnH3zF");
                      reg2179 <= ((reg2184[(3'h7):(2'h3)] ?
                          ((reg2140 + reg2109) ?
                              $unsigned(forvar2174) : reg2173) : $signed(forvar2166[(1'h0):(1'h0)])) * reg2171[(4'hc):(3'h5)]);
                      reg2180 = reg2170;
                    end
                  else
                    begin
                      reg2177 = ((+$signed($unsigned(reg2139))) ^~ $signed(forvar2153));
                    end
                  if (forvar2166[(4'hd):(3'h4)])
                    begin
                      reg2184 = $signed(($unsigned($signed((8'ha8))) + $unsigned(forvar2158[(4'hc):(4'hc)])));
                      reg2187 <= $signed((8'ha5));
                      reg2188 = $unsigned($unsigned(($unsigned(wire2) ?
                          $signed(reg2114) : {forvar2174})));
                    end
                  else
                    begin
                      reg2184 = "XRd";
                      reg2185 = "oZ3maP4VpPY3Dh";
                      reg2186 = $unsigned("TlNkKFeuLd6");
                    end
                  for (forvar2189 = (1'h0); (forvar2189 < (2'h2)); forvar2189 = (forvar2189 + (1'h1)))
                    begin
                      reg2190 = (~^reg2106[(4'h8):(2'h3)]);
                    end
                  if (reg2147)
                    begin
                      reg2191 = ((~"1fxOdr9YJnL") || (reg2151[(1'h0):(1'h0)] ?
                          reg2173[(3'h4):(1'h1)] : reg2141[(1'h1):(1'h0)]));
                      reg2192 = reg2171;
                      reg2193 = $unsigned(reg2181[(3'h4):(2'h2)]);
                      reg2194 <= reg2192;
                    end
                  else
                    begin
                      reg2191 = (&(8'hb6));
                    end
                end
            end
        end
      for (forvar2195 = (1'h0); (forvar2195 < (2'h2)); forvar2195 = (forvar2195 + (1'h1)))
        begin
          reg2196 = forvar2152;
          for (forvar2197 = (1'h0); (forvar2197 < (2'h2)); forvar2197 = (forvar2197 + (1'h1)))
            begin
              reg2198 = $unsigned(reg2113);
              reg2199 <= reg2115[(4'h9):(3'h7)];
              if (forvar2148)
                begin
                  for (forvar2200 = (1'h0); (forvar2200 < (2'h3)); forvar2200 = (forvar2200 + (1'h1)))
                    begin
                      reg2201 = "0uPByk";
                      reg2202 = (!$unsigned((^$unsigned(forvar2175))));
                      reg2203 <= (^"yu");
                      reg2204 = (+$signed(((reg2113 + reg2154) ?
                          $signed(forvar2136) : $signed(reg2121))));
                    end
                end
              else
                begin
                  for (forvar2200 = (1'h0); (forvar2200 < (1'h0)); forvar2200 = (forvar2200 + (1'h1)))
                    begin
                      reg2201 = {(-(reg2177[(1'h0):(1'h0)] ?
                              $unsigned(reg2192) : $signed(reg2121)))};
                      reg2202 = forvar2137;
                      reg2204 = (|(reg2151[(2'h3):(1'h1)] ^ ((reg2190 && reg2128) >= (8'ha7))));
                      reg2205 <= reg2198[(3'h4):(2'h2)];
                    end
                  reg2206 = reg2121[(4'h8):(3'h4)];
                  for (forvar2207 = (1'h0); (forvar2207 < (1'h1)); forvar2207 = (forvar2207 + (1'h1)))
                    begin
                      reg2208 <= (8'hb7);
                      reg2209 = {"W"};
                      reg2210 = ($signed((^reg2202[(1'h0):(1'h0)])) >= $unsigned(($signed(forvar2207) ?
                          $unsigned(reg2149) : (|(8'h9f)))));
                    end
                  reg2211 <= $signed("3Tt0RN04Y");
                end
            end
          if ((8'ha7))
            begin
              reg2212 = ($signed(reg2206[(1'h0):(1'h0)]) ?
                  $unsigned(((reg2199 <<< reg2147) ?
                      (&reg2128) : reg2147)) : forvar2104[(2'h3):(2'h2)]);
            end
          else
            begin
              for (forvar2212 = (1'h0); (forvar2212 < (2'h2)); forvar2212 = (forvar2212 + (1'h1)))
                begin
                  reg2213 = $signed((~^((reg2210 ? reg2194 : reg2110) ?
                      reg2193 : forvar2158)));
                  reg2214 <= {reg2140[(4'hb):(1'h1)]};
                  for (forvar2215 = (1'h0); (forvar2215 < (1'h1)); forvar2215 = (forvar2215 + (1'h1)))
                    begin
                      reg2216 <= ((~wire2103[(2'h3):(2'h2)]) ?
                          reg2115[(3'h5):(1'h0)] : $unsigned((|reg2173[(2'h3):(2'h3)])));
                    end
                  reg2217 <= reg2166;
                end
              for (forvar2218 = (1'h0); (forvar2218 < (2'h3)); forvar2218 = (forvar2218 + (1'h1)))
                begin
                  if ($signed($signed(($unsigned(reg2162) <= {reg2126}))))
                    begin
                      reg2219 = forvar2166;
                    end
                  else
                    begin
                      reg2220 <= ("gRiY5M9H5aLx" ?
                          $unsigned(forvar2166) : ((~|"ZpTuG1") == forvar2107));
                      reg2221 = "V";
                      reg2222 = ((~^$signed(reg2173)) - $signed(((|forvar2136) ?
                          ((8'hae) == (8'ha4)) : $unsigned((8'hb1)))));
                      reg2223 = "UzMmTEDS4OsSC8t";
                    end
                  reg2224 = reg2129[(2'h2):(1'h1)];
                  if ((~|reg2219))
                    begin
                      reg2225 <= reg2212[(3'h5):(1'h0)];
                      reg2226 <= $signed(($unsigned((|reg2133)) || reg2183[(3'h5):(1'h1)]));
                      reg2227 = (^$unsigned({$unsigned(reg2190)}));
                    end
                  else
                    begin
                      reg2227 = reg2154;
                      reg2228 <= {((!reg2137[(1'h0):(1'h0)]) * (^$signed(forvar2195)))};
                      reg2229 = $signed((~|reg2179[(4'h8):(3'h7)]));
                    end
                  for (forvar2230 = (1'h0); (forvar2230 < (2'h3)); forvar2230 = (forvar2230 + (1'h1)))
                    begin
                      reg2231 = reg2179;
                      reg2232 = {$unsigned(reg2127)};
                    end
                end
            end
        end
      reg2233 <= "QmF42SnzSu8AlBD";
    end
  module651 #() modinst2235 (.wire654(wire1), .wire652(reg2122), .clk(clk), .y(wire2234), .wire655(reg2136), .wire653(reg2194));
  always
    @(posedge clk) begin
      reg2236 = reg2107[(1'h0):(1'h0)];
      reg2237 <= wire1[(3'h4):(2'h3)];
      reg2238 = wire2234;
      if ((reg2199 ~^ ($unsigned((reg2109 | reg2126)) ?
          $unsigned($unsigned(reg2105)) : $unsigned((reg2226 <<< reg2205)))))
        begin
          reg2239 = $unsigned(((8'hac) & reg2104));
          reg2240 = $signed(($unsigned((~|reg2181)) && $unsigned($unsigned(reg2126))));
          reg2241 <= ((^~"7R4RIYqKcY4") >> "YPa");
          for (forvar2242 = (1'h0); (forvar2242 < (2'h3)); forvar2242 = (forvar2242 + (1'h1)))
            begin
              reg2243 <= ((|(reg2105 >= "fam49WqAWz0AEeJ")) >= ("v" >> $unsigned($unsigned(reg2138))));
              if (reg2132)
                begin
                  reg2244 = reg2225[(4'h9):(3'h4)];
                  reg2245 = $signed($signed({reg2136[(4'hb):(2'h3)]}));
                  if ($signed({$unsigned(reg2150)}))
                    begin
                      reg2246 = ((($unsigned(reg2136) != ((8'hba) ?
                          wire2103 : reg2172)) > reg2214) && $unsigned(wire3[(4'h9):(4'h9)]));
                      reg2247 <= ({$unsigned((+wire0))} ?
                          (reg2243 && ($unsigned((8'haa)) ?
                              {reg2109} : (^reg2104))) : "o4CLgRKIzJQ1");
                    end
                  else
                    begin
                      reg2246 = $unsigned("Y8dVuNH3adRecZe");
                    end
                end
              else
                begin
                  reg2244 = $unsigned(reg2168);
                end
              for (forvar2248 = (1'h0); (forvar2248 < (2'h2)); forvar2248 = (forvar2248 + (1'h1)))
                begin
                  for (forvar2249 = (1'h0); (forvar2249 < (1'h1)); forvar2249 = (forvar2249 + (1'h1)))
                    begin
                      reg2250 = $unsigned((~^(reg2187[(4'hb):(3'h5)] < ((8'hac) ?
                          reg2233 : reg2247))));
                      reg2251 = (reg2114[(4'hc):(4'ha)] <= reg2150[(3'h5):(1'h1)]);
                      reg2252 = {$signed(wire2)};
                    end
                  reg2253 <= {$unsigned(reg2220[(2'h2):(1'h0)])};
                  reg2254 = (^~((|(!reg2251)) - ($signed(reg2239) ?
                      $unsigned((8'ha5)) : wire0)));
                  if ((($signed("ALHu1r4mPUS8") ?
                          (reg2176[(2'h3):(2'h3)] ?
                              (^(8'hac)) : wire2103[(1'h1):(1'h0)]) : (+(wire2234 ?
                              reg2161 : wire0))) ?
                      (((reg2243 ?
                          reg2136 : forvar2242) <= (&forvar2249)) - reg2172[(2'h3):(1'h0)]) : reg2172[(3'h4):(2'h3)]))
                    begin
                      reg2255 = ({((reg2161 ?
                              reg2107 : reg2217) <= "")} == reg2187);
                      reg2256 <= ($signed({(reg2220 ^ reg2114)}) ?
                          (((reg2137 >= reg2208) ^ $unsigned(reg2126)) + ((reg2107 ~^ reg2246) ?
                              $unsigned(reg2187) : (-reg2236))) : $unsigned($unsigned((^~reg2247))));
                      reg2257 = (^~{$signed($signed(reg2205))});
                    end
                  else
                    begin
                      reg2256 <= reg2118[(2'h2):(1'h0)];
                    end
                end
            end
        end
      else
        begin
          if (("yoX1Pcfyl" ? $signed((8'haa)) : $signed($unsigned(reg2183))))
            begin
              reg2239 = {$signed($signed($signed(forvar2249)))};
              for (forvar2240 = (1'h0); (forvar2240 < (2'h3)); forvar2240 = (forvar2240 + (1'h1)))
                begin
                  reg2242 = reg2164[(1'h1):(1'h0)];
                end
              reg2244 = ({reg2132[(2'h2):(1'h1)]} ?
                  ($unsigned({reg2239}) ?
                      {reg2161} : forvar2240) : $signed($unsigned((+reg2236))));
              reg2245 = {(|{reg2236})};
            end
          else
            begin
              if ($unsigned("3OPI4X3uDu"))
                begin
                  reg2241 <= {{((reg2131 | reg2239) > (reg2252 >= (8'hae)))}};
                  for (forvar2242 = (1'h0); (forvar2242 < (2'h2)); forvar2242 = (forvar2242 + (1'h1)))
                    begin
                      reg2244 = $unsigned(("YM1" ?
                          "eyxKZF6DUSxoN1" : $signed($signed((8'hba)))));
                      reg2245 = (|wire3);
                      reg2247 <= $signed(reg2199);
                    end
                end
              else
                begin
                  reg2241 <= $unsigned($signed(((8'hb0) ~^ ((8'hb0) <= (8'hac)))));
                  for (forvar2242 = (1'h0); (forvar2242 < (2'h3)); forvar2242 = (forvar2242 + (1'h1)))
                    begin
                      reg2244 = {(8'hab)};
                    end
                  for (forvar2245 = (1'h0); (forvar2245 < (2'h2)); forvar2245 = (forvar2245 + (1'h1)))
                    begin
                      reg2247 <= ($signed(reg2158[(3'h7):(3'h5)]) <= reg2253[(1'h0):(1'h0)]);
                      reg2248 = $signed($signed("KxG"));
                      reg2249 = (+("UrB" | reg2252));
                    end
                end
              for (forvar2250 = (1'h0); (forvar2250 < (1'h0)); forvar2250 = (forvar2250 + (1'h1)))
                begin
                  for (forvar2251 = (1'h0); (forvar2251 < (1'h0)); forvar2251 = (forvar2251 + (1'h1)))
                    begin
                      reg2252 = $unsigned($signed(($signed(wire1) ?
                          reg2216 : "luaG")));
                      reg2254 = (reg2248[(3'h4):(1'h1)] ?
                          reg2199[(2'h2):(1'h1)] : {wire2103[(2'h2):(1'h0)]});
                      reg2255 = (reg2243 ~^ (&{wire0[(3'h4):(2'h2)]}));
                    end
                  for (forvar2256 = (1'h0); (forvar2256 < (2'h3)); forvar2256 = (forvar2256 + (1'h1)))
                    begin
                      reg2258 <= $unsigned(reg2211[(4'h9):(4'h9)]);
                      reg2259 <= $signed($signed($unsigned((^~reg2255))));
                      reg2260 = reg2105;
                      reg2261 <= $unsigned(reg2238);
                    end
                end
            end
          if ($signed(({reg2238} ? $unsigned($unsigned(reg2238)) : reg2228)))
            begin
              for (forvar2262 = (1'h0); (forvar2262 < (1'h1)); forvar2262 = (forvar2262 + (1'h1)))
                begin
                  reg2263 <= reg2132;
                  reg2264 <= wire0[(2'h3):(2'h2)];
                  for (forvar2265 = (1'h0); (forvar2265 < (1'h1)); forvar2265 = (forvar2265 + (1'h1)))
                    begin
                      reg2266 = {(reg2264[(4'ha):(2'h2)] == "o2PMXxpHtH")};
                      reg2267 = (^~reg2176[(2'h3):(1'h1)]);
                    end
                end
              if ($signed(((~(reg2203 * reg2238)) ?
                  "" : (wire2101 != reg2109))))
                begin
                  for (forvar2268 = (1'h0); (forvar2268 < (2'h2)); forvar2268 = (forvar2268 + (1'h1)))
                    begin
                      reg2269 <= (^~(((~&(8'ha4)) < reg2116) ? "i" : reg2109));
                      reg2270 <= $signed((-$signed((reg2164 > reg2239))));
                    end
                  if (reg2254)
                    begin
                      reg2271 <= $signed($unsigned((8'h9d)));
                      reg2272 <= "PNm";
                    end
                  else
                    begin
                      reg2271 <= (+{"tigOF3t9BPF"});
                    end
                  for (forvar2273 = (1'h0); (forvar2273 < (1'h0)); forvar2273 = (forvar2273 + (1'h1)))
                    begin
                      reg2274 = (|$unsigned({reg2220[(1'h0):(1'h0)]}));
                      reg2275 = (reg2208[(1'h1):(1'h0)] ?
                          "9DFP" : ($signed("v") <= "VgoLLwcE4d9d"));
                      reg2276 = ("h" ^~ {(forvar2265 ?
                              ((8'ha8) <= forvar2251) : (reg2242 ^ reg2241))});
                      reg2277 <= reg2160;
                    end
                  reg2278 = "6Cw0qJ6g";
                end
              else
                begin
                  reg2268 = reg2278[(2'h2):(1'h1)];
                  for (forvar2269 = (1'h0); (forvar2269 < (1'h0)); forvar2269 = (forvar2269 + (1'h1)))
                    begin
                      reg2273 = (("feeHXGIu" ?
                          ((|reg2246) >> ((8'ha7) > reg2182)) : (!"Ex")) && reg2245);
                    end
                  for (forvar2274 = (1'h0); (forvar2274 < (2'h2)); forvar2274 = (forvar2274 + (1'h1)))
                    begin
                      reg2275 = reg2237;
                      reg2277 <= {reg2181};
                    end
                  for (forvar2278 = (1'h0); (forvar2278 < (1'h0)); forvar2278 = (forvar2278 + (1'h1)))
                    begin
                      reg2279 = {$unsigned($signed(reg2105[(2'h2):(1'h1)]))};
                      reg2280 = $unsigned((-(^~((8'had) ? reg2272 : reg2237))));
                      reg2281 = reg2238;
                    end
                end
              reg2282 = (!(reg2260[(1'h1):(1'h0)] ?
                  (forvar2250[(4'h9):(4'h8)] ?
                      (reg2124 ? reg2263 : reg2250) : (8'hba)) : (~{reg2199})));
            end
          else
            begin
              for (forvar2262 = (1'h0); (forvar2262 < (1'h0)); forvar2262 = (forvar2262 + (1'h1)))
                begin
                  reg2263 <= (reg2158 <<< $signed($signed((reg2280 ?
                      reg2107 : reg2258))));
                  for (forvar2264 = (1'h0); (forvar2264 < (2'h2)); forvar2264 = (forvar2264 + (1'h1)))
                    begin
                      reg2265 = reg2277[(2'h3):(2'h3)];
                      reg2266 = {(+$unsigned(reg2263[(2'h2):(1'h0)]))};
                    end
                  for (forvar2267 = (1'h0); (forvar2267 < (2'h3)); forvar2267 = (forvar2267 + (1'h1)))
                    begin
                      reg2268 = $unsigned({reg2243[(1'h1):(1'h1)]});
                    end
                end
              reg2269 <= "OxzXkyHyG";
            end
          reg2283 = reg2250;
        end
    end
  assign wire2284 = reg2159[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg2285 <= $signed($unsigned({(reg2269 ? reg2115 : reg2161)}));
      reg2286 = (&($unsigned($unsigned(reg2131)) ?
          reg2176 : (&(reg2167 ? reg2136 : reg2243))));
    end
  module275 #() modinst2288 (.wire276(reg2263), .wire278(reg2132), .wire277(reg2214), .clk(clk), .wire279(reg2115), .y(wire2287));
  module651 #() modinst2290 (wire2289, clk, reg2131, reg2225, reg2237, wire2287);
  assign wire2291 = reg2116[(3'h6):(3'h6)];
  assign wire2292 = $signed($signed("GSJ3FrH1fAYDsa2"));
  always
    @(posedge clk) begin
      if ((8'haa))
        begin
          reg2293 <= reg2159;
          for (forvar2294 = (1'h0); (forvar2294 < (1'h1)); forvar2294 = (forvar2294 + (1'h1)))
            begin
              reg2295 <= "8Yi1LvhSlbhfu";
            end
          reg2296 = reg2136[(4'ha):(1'h0)];
        end
      else
        begin
          for (forvar2293 = (1'h0); (forvar2293 < (1'h1)); forvar2293 = (forvar2293 + (1'h1)))
            begin
              if (reg2261)
                begin
                  if (forvar2293[(1'h1):(1'h0)])
                    begin
                      reg2294 = (^~(8'ha0));
                    end
                  else
                    begin
                      reg2295 <= $signed($unsigned($unsigned((^~reg2183))));
                      reg2297 <= $unsigned(reg2199);
                      reg2298 = $signed((~&$unsigned(forvar2294[(2'h2):(2'h2)])));
                      reg2299 <= (-reg2107[(2'h2):(2'h2)]);
                    end
                  if ({(~^(|(-(8'hb1))))})
                    begin
                      reg2300 <= "R6FnQQXY";
                      reg2301 <= (($unsigned((8'ha1)) < (~reg2114[(4'hd):(4'h8)])) ?
                          (~^(wire3[(3'h6):(1'h0)] ?
                              reg2137 : $signed(reg2176))) : (($unsigned((8'hb5)) << (reg2194 ?
                              reg2133 : (8'hb2))) && ($unsigned(wire2103) < (^~reg2285))));
                    end
                  else
                    begin
                      reg2300 <= (~("" ^~ (|$unsigned(reg2228))));
                    end
                  if ($unsigned((((8'ha2) >> wire1[(3'h5):(1'h0)]) ?
                      {(reg2183 ? reg2256 : reg2131)} : ({reg2233} | ""))))
                    begin
                      reg2302 = (wire2289[(3'h5):(1'h0)] ?
                          reg2217 : $signed((reg2136 >= (~^reg2118))));
                      reg2303 = $unsigned(wire2289);
                    end
                  else
                    begin
                      reg2302 = (~^(8'haa));
                      reg2303 = ("negZAnyFDkq" <= ("lFoFAtosSLqrwkd" + reg2124));
                      reg2304 = {reg2241};
                    end
                end
              else
                begin
                  if (reg2225)
                    begin
                      reg2294 = $signed(reg2299);
                      reg2295 <= $unsigned(wire2291[(4'hb):(1'h1)]);
                      reg2297 <= reg2228;
                    end
                  else
                    begin
                      reg2294 = "I4Nq9gq7eETTo";
                      reg2296 = reg2228[(2'h2):(2'h2)];
                    end
                  reg2298 = $unsigned((^reg2203[(1'h0):(1'h0)]));
                  for (forvar2299 = (1'h0); (forvar2299 < (2'h3)); forvar2299 = (forvar2299 + (1'h1)))
                    begin
                      reg2302 = "H";
                    end
                  reg2305 <= (8'h9f);
                end
            end
          reg2306 = $unsigned((((reg2217 ? wire3 : reg2194) == {reg2133}) ?
              reg2137 : reg2304[(4'ha):(4'ha)]));
          reg2307 <= $signed("SuKXvKxX");
          reg2308 = reg2299;
        end
      reg2309 = ((8'hb3) ? wire1[(1'h1):(1'h1)] : reg2116);
    end
  assign wire2310 = $unsigned($signed(reg2243[(3'h6):(1'h1)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4  (y, clk, wire8, wire7, wire6, wire5);
  output wire [(32'hb62):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire8;
  input wire signed [(4'h9):(1'h0)] wire7;
  input wire [(4'hf):(1'h0)] wire6;
  input wire signed [(3'h6):(1'h0)] wire5;
  wire [(4'he):(1'h0)] wire2099;
  wire signed [(2'h2):(1'h0)] wire2025;
  wire signed [(3'h5):(1'h0)] wire2024;
  wire signed [(2'h3):(1'h0)] wire2022;
  wire [(3'h7):(1'h0)] wire10;
  wire [(4'hb):(1'h0)] wire9;
  reg signed [(4'hd):(1'h0)] reg211 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg208 = (1'h0);
  reg [(4'hd):(1'h0)] reg204 = (1'h0);
  reg [(4'hf):(1'h0)] reg199 = (1'h0);
  reg [(5'h10):(1'h0)] reg187 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg182 = (1'h0);
  reg [(4'he):(1'h0)] reg179 = (1'h0);
  reg signed [(4'he):(1'h0)] reg176 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg171 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg170 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg169 = (1'h0);
  reg [(2'h2):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg162 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg160 = (1'h0);
  reg signed [(4'he):(1'h0)] reg158 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg154 = (1'h0);
  reg [(4'hd):(1'h0)] reg148 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg147 = (1'h0);
  reg [(4'hd):(1'h0)] reg145 = (1'h0);
  reg [(4'hd):(1'h0)] reg141 = (1'h0);
  reg [(4'he):(1'h0)] reg138 = (1'h0);
  reg [(3'h6):(1'h0)] reg122 = (1'h0);
  reg [(4'h8):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg135 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg133 = (1'h0);
  reg [(2'h3):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg126 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg125 = (1'h0);
  reg [(4'he):(1'h0)] reg124 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg120 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg119 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg82 = (1'h0);
  reg [(4'ha):(1'h0)] reg108 = (1'h0);
  reg signed [(4'he):(1'h0)] reg111 = (1'h0);
  reg [(3'h4):(1'h0)] reg105 = (1'h0);
  reg [(4'he):(1'h0)] reg102 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg101 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg99 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg93 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg90 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg87 = (1'h0);
  reg [(4'hd):(1'h0)] reg97 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg96 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg95 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg94 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg83 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg76 = (1'h0);
  reg [(3'h7):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg68 = (1'h0);
  reg [(4'h8):(1'h0)] reg66 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg61 = (1'h0);
  reg [(4'hb):(1'h0)] reg45 = (1'h0);
  reg [(5'h10):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg51 = (1'h0);
  reg [(4'h8):(1'h0)] reg50 = (1'h0);
  reg [(4'h8):(1'h0)] reg48 = (1'h0);
  reg [(5'h10):(1'h0)] reg42 = (1'h0);
  reg [(2'h3):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg36 = (1'h0);
  reg signed [(4'he):(1'h0)] reg35 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg30 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg29 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg25 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg24 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg21 = (1'h0);
  reg [(4'h9):(1'h0)] reg20 = (1'h0);
  reg [(3'h6):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg14 = (1'h0);
  reg [(3'h6):(1'h0)] reg2030 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2039 = (1'h0);
  reg [(2'h2):(1'h0)] reg2042 = (1'h0);
  reg [(4'hc):(1'h0)] reg2043 = (1'h0);
  reg [(3'h5):(1'h0)] reg2051 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2054 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2056 = (1'h0);
  reg [(4'hb):(1'h0)] reg2059 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2060 = (1'h0);
  reg [(4'h9):(1'h0)] reg2065 = (1'h0);
  reg [(4'he):(1'h0)] reg2068 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2072 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2074 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2079 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2085 = (1'h0);
  reg [(4'hb):(1'h0)] reg2090 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2095 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2097 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2098 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2076 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2075 = (1'h0);
  reg [(4'hb):(1'h0)] reg2096 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2091 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2087 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2082 = (1'h0);
  reg [(2'h3):(1'h0)] reg2094 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2093 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2092 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2091 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2089 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2088 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2087 = (1'h0);
  reg [(3'h6):(1'h0)] reg2086 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2084 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2083 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2082 = (1'h0);
  reg [(4'hb):(1'h0)] reg2081 = (1'h0);
  reg [(4'he):(1'h0)] reg2080 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2078 = (1'h0);
  reg [(2'h3):(1'h0)] reg2077 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2076 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2075 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2073 = (1'h0);
  reg [(4'ha):(1'h0)] reg2071 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2063 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2062 = (1'h0);
  reg [(5'h10):(1'h0)] reg2070 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2069 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2067 = (1'h0);
  reg [(3'h5):(1'h0)] reg2066 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2064 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2063 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2062 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2061 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2058 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2057 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2055 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2053 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2052 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2050 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2049 = (1'h0);
  reg [(3'h7):(1'h0)] reg2048 = (1'h0);
  reg [(3'h7):(1'h0)] reg2047 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2046 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2045 = (1'h0);
  reg [(4'h9):(1'h0)] reg2044 = (1'h0);
  reg [(4'h8):(1'h0)] reg2041 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2040 = (1'h0);
  reg [(4'ha):(1'h0)] reg2038 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2037 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2036 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2035 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2034 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2033 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2032 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2031 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2029 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2028 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2027 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2026 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg213 = (1'h0);
  reg [(4'hf):(1'h0)] reg212 = (1'h0);
  reg [(3'h4):(1'h0)] reg210 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg209 = (1'h0);
  reg [(4'h9):(1'h0)] forvar207 = (1'h0);
  reg [(2'h3):(1'h0)] reg206 = (1'h0);
  reg [(4'h8):(1'h0)] reg205 = (1'h0);
  reg [(4'hc):(1'h0)] forvar203 = (1'h0);
  reg [(3'h6):(1'h0)] reg202 = (1'h0);
  reg signed [(4'he):(1'h0)] reg201 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg198 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg197 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar196 = (1'h0);
  reg [(3'h7):(1'h0)] forvar195 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg194 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg192 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg191 = (1'h0);
  reg [(4'he):(1'h0)] forvar190 = (1'h0);
  reg [(3'h6):(1'h0)] reg189 = (1'h0);
  reg [(3'h7):(1'h0)] reg184 = (1'h0);
  reg [(3'h4):(1'h0)] reg188 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg186 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg185 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar184 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar183 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg181 = (1'h0);
  reg [(4'he):(1'h0)] forvar178 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg177 = (1'h0);
  reg [(4'he):(1'h0)] forvar175 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar173 = (1'h0);
  reg [(4'h8):(1'h0)] reg172 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg167 = (1'h0);
  reg [(3'h7):(1'h0)] reg180 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg178 = (1'h0);
  reg [(3'h5):(1'h0)] forvar177 = (1'h0);
  reg [(4'h8):(1'h0)] reg175 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg174 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg173 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar172 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg168 = (1'h0);
  reg [(4'hc):(1'h0)] forvar167 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg166 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar165 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg164 = (1'h0);
  reg [(3'h4):(1'h0)] reg163 = (1'h0);
  reg [(3'h4):(1'h0)] forvar161 = (1'h0);
  reg [(4'hf):(1'h0)] reg159 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar157 = (1'h0);
  reg [(3'h6):(1'h0)] reg156 = (1'h0);
  reg [(3'h5):(1'h0)] forvar155 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg153 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg152 = (1'h0);
  reg [(4'hb):(1'h0)] reg151 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar150 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar149 = (1'h0);
  reg [(2'h2):(1'h0)] reg146 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg144 = (1'h0);
  reg [(3'h6):(1'h0)] forvar143 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar142 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar140 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar139 = (1'h0);
  reg [(3'h6):(1'h0)] forvar119 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg127 = (1'h0);
  reg [(3'h7):(1'h0)] reg137 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg136 = (1'h0);
  reg [(4'hf):(1'h0)] reg134 = (1'h0);
  reg [(2'h2):(1'h0)] reg132 = (1'h0);
  reg [(5'h10):(1'h0)] forvar131 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg130 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg129 = (1'h0);
  reg [(4'hf):(1'h0)] forvar127 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg123 = (1'h0);
  reg [(4'hd):(1'h0)] forvar122 = (1'h0);
  reg [(4'hf):(1'h0)] reg121 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg118 = (1'h0);
  reg [(3'h6):(1'h0)] forvar117 = (1'h0);
  reg [(4'hf):(1'h0)] forvar116 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg115 = (1'h0);
  reg [(4'hb):(1'h0)] reg114 = (1'h0);
  reg [(4'ha):(1'h0)] reg113 = (1'h0);
  reg [(3'h7):(1'h0)] forvar112 = (1'h0);
  reg [(3'h5):(1'h0)] reg104 = (1'h0);
  reg [(4'hf):(1'h0)] reg110 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg109 = (1'h0);
  reg [(4'he):(1'h0)] forvar108 = (1'h0);
  reg [(3'h5):(1'h0)] reg107 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg106 = (1'h0);
  reg [(3'h7):(1'h0)] forvar104 = (1'h0);
  reg [(3'h4):(1'h0)] reg103 = (1'h0);
  reg [(2'h3):(1'h0)] reg100 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg98 = (1'h0);
  reg [(3'h4):(1'h0)] forvar94 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar93 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg92 = (1'h0);
  reg [(5'h10):(1'h0)] reg91 = (1'h0);
  reg [(3'h5):(1'h0)] forvar90 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg89 = (1'h0);
  reg [(3'h5):(1'h0)] reg88 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar87 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg86 = (1'h0);
  reg [(2'h2):(1'h0)] reg85 = (1'h0);
  reg [(4'hf):(1'h0)] forvar84 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar82 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg81 = (1'h0);
  reg [(2'h3):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg79 = (1'h0);
  reg [(5'h10):(1'h0)] forvar77 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg72 = (1'h0);
  reg [(4'hc):(1'h0)] reg78 = (1'h0);
  reg [(4'he):(1'h0)] reg75 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg74 = (1'h0);
  reg [(4'h9):(1'h0)] forvar72 = (1'h0);
  reg [(5'h10):(1'h0)] reg71 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg70 = (1'h0);
  reg [(2'h2):(1'h0)] reg69 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar67 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg65 = (1'h0);
  reg [(3'h7):(1'h0)] reg64 = (1'h0);
  reg [(2'h2):(1'h0)] forvar63 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg62 = (1'h0);
  reg [(3'h7):(1'h0)] forvar58 = (1'h0);
  reg [(2'h3):(1'h0)] reg54 = (1'h0);
  reg [(2'h3):(1'h0)] forvar53 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg49 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg60 = (1'h0);
  reg [(3'h6):(1'h0)] reg59 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar57 = (1'h0);
  reg [(2'h2):(1'h0)] forvar56 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar54 = (1'h0);
  reg [(5'h10):(1'h0)] reg53 = (1'h0);
  reg [(2'h3):(1'h0)] reg52 = (1'h0);
  reg [(4'hc):(1'h0)] forvar49 = (1'h0);
  reg [(4'hf):(1'h0)] reg47 = (1'h0);
  reg [(4'hf):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar45 = (1'h0);
  reg [(3'h6):(1'h0)] forvar44 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg43 = (1'h0);
  reg [(4'hd):(1'h0)] forvar40 = (1'h0);
  reg [(4'hc):(1'h0)] reg39 = (1'h0);
  reg [(5'h10):(1'h0)] reg38 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg37 = (1'h0);
  reg [(3'h7):(1'h0)] reg34 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg33 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar21 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar13 = (1'h0);
  reg [(4'hd):(1'h0)] reg31 = (1'h0);
  reg [(2'h3):(1'h0)] reg28 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar27 = (1'h0);
  reg [(5'h10):(1'h0)] forvar26 = (1'h0);
  reg [(3'h7):(1'h0)] reg23 = (1'h0);
  reg [(2'h2):(1'h0)] reg22 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg18 = (1'h0);
  reg [(4'he):(1'h0)] reg17 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg15 = (1'h0);
  reg [(4'hb):(1'h0)] reg13 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar12 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg11 = (1'h0);
  assign y = {wire2024,
                 reg211,
                 reg208,
                 reg182,
                 reg171,
                 reg170,
                 reg169,
                 reg161,
                 reg162,
                 reg160,
                 reg158,
                 reg154,
                 reg148,
                 reg131,
                 reg128,
                 reg120,
                 reg108,
                 reg76,
                 reg68,
                 reg61,
                 reg50,
                 reg42,
                 reg36,
                 reg30,
                 reg29,
                 reg21,
                 reg16,
                 reg2051,
                 reg2056,
                 reg2059,
                 reg2065,
                 reg2095,
                 forvar2075,
                 reg2091,
                 reg2086,
                 forvar2082,
                 reg2081,
                 reg2080,
                 reg2077,
                 reg2076,
                 forvar2073,
                 reg2062,
                 reg2070,
                 forvar2069,
                 reg2063,
                 reg2061,
                 reg2048,
                 reg2046,
                 reg2035,
                 reg2033,
                 forvar2032,
                 forvar2026,
                 reg210,
                 reg209,
                 reg201,
                 reg200,
                 forvar195,
                 forvar190,
                 reg186,
                 reg185,
                 reg181,
                 forvar175,
                 reg172,
                 reg178,
                 forvar177,
                 forvar172,
                 reg166,
                 reg164,
                 reg163,
                 forvar157,
                 reg156,
                 reg151,
                 reg146,
                 forvar143,
                 forvar140,
                 forvar139,
                 forvar119,
                 reg134,
                 forvar131,
                 reg130,
                 forvar116,
                 reg114,
                 reg104,
                 forvar108,
                 reg84,
                 reg91,
                 forvar84,
                 reg80,
                 reg74,
                 forvar67,
                 forvar58,
                 reg54,
                 reg59,
                 reg55,
                 reg53,
                 reg47,
                 reg46,
                 forvar45,
                 reg39,
                 reg38,
                 reg37,
                 reg34,
                 forvar13,
                 reg17,
                 reg15,
                 reg13,
                 forvar12,
                 (1'h0)};
  assign wire9 = "JKQz";
  assign wire10 = ((8'hac) <<< {($signed(wire7) ?
                          wire6[(4'hb):(3'h6)] : {wire9})});
  always
    @(posedge clk) begin
      if ($signed(($unsigned("6t6u4HnC4w0m4Q") < $unsigned(wire6))))
        begin
          reg11 = wire8;
          for (forvar12 = (1'h0); (forvar12 < (2'h3)); forvar12 = (forvar12 + (1'h1)))
            begin
              if ("rW4V6guowV")
                begin
                  if (forvar12)
                    begin
                      reg13 = wire9;
                      reg14 <= $signed(($signed(forvar12[(3'h5):(1'h0)]) & "2qXiaNhHH"));
                    end
                  else
                    begin
                      reg13 = reg14;
                      reg15 = ((+reg14[(4'hf):(4'hd)]) != $unsigned(wire7));
                      reg16 <= reg14;
                    end
                  reg17 = wire8;
                end
              else
                begin
                  if (($unsigned((~{reg11})) ?
                      ((^(reg13 - reg16)) ^~ $unsigned($signed((8'ha9)))) : (~((wire6 - wire7) != (~reg16)))))
                    begin
                      reg14 <= ((reg15 == reg17) >> reg13[(3'h7):(1'h0)]);
                      reg16 <= wire9[(3'h5):(3'h4)];
                      reg17 = (~^(~&(reg17 >>> $unsigned(wire8))));
                      reg18 = wire9[(3'h7):(3'h7)];
                    end
                  else
                    begin
                      reg13 = ((8'ha4) && (|($signed((8'ha7)) == "NXoLz48iEH4PDla")));
                      reg15 = (~|(wire6[(3'h4):(1'h1)] ?
                          (^~$unsigned((8'hac))) : $unsigned(wire9)));
                      reg17 = (wire9[(4'h9):(4'h8)] ?
                          reg18[(3'h5):(2'h2)] : wire7);
                      reg19 <= reg14[(2'h2):(1'h0)];
                    end
                  reg20 <= "08KgAP9DVcN";
                  if ((~&(((!(8'hb2)) ? (^~wire7) : $unsigned(reg11)) ?
                      reg13 : (+wire6[(4'hb):(3'h4)]))))
                    begin
                      reg21 <= $unsigned(reg13[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg22 = "wZ04r";
                      reg23 = $signed(reg22);
                      reg24 <= "";
                    end
                end
            end
          reg25 <= $unsigned((&(((8'hb9) >>> reg17) ?
              ((8'hab) == (8'ha0)) : reg20)));
          for (forvar26 = (1'h0); (forvar26 < (2'h2)); forvar26 = (forvar26 + (1'h1)))
            begin
              for (forvar27 = (1'h0); (forvar27 < (1'h1)); forvar27 = (forvar27 + (1'h1)))
                begin
                  if (wire6)
                    begin
                      reg28 = {wire10};
                    end
                  else
                    begin
                      reg28 = reg19[(2'h2):(1'h0)];
                      reg29 <= forvar26;
                      reg30 <= {$unsigned((~|reg29))};
                    end
                  reg31 = forvar12;
                end
            end
        end
      else
        begin
          reg11 = reg24[(2'h2):(1'h0)];
          for (forvar12 = (1'h0); (forvar12 < (2'h3)); forvar12 = (forvar12 + (1'h1)))
            begin
              for (forvar13 = (1'h0); (forvar13 < (1'h0)); forvar13 = (forvar13 + (1'h1)))
                begin
                  if ($signed(((^"sJd9pPYf2WZxO5n") >> forvar27)))
                    begin
                      reg15 = ("KRHN" + (&(&reg30)));
                      reg16 <= "qCxnvx";
                      reg19 <= ($signed(((^reg30) * {reg22})) ?
                          $unsigned($unsigned((reg29 ?
                              reg15 : reg20))) : (~|((-reg24) ?
                              wire6[(3'h7):(2'h3)] : "")));
                    end
                  else
                    begin
                      reg14 <= $unsigned($signed(wire5));
                      reg15 = ((~&((wire8 ? (8'ha3) : reg15) ?
                              "3Mu6N" : (+reg18))) ?
                          forvar27 : reg30);
                      reg17 = reg21;
                      reg18 = "tXomRzZV";
                    end
                end
              reg20 <= reg18[(1'h0):(1'h0)];
              for (forvar21 = (1'h0); (forvar21 < (2'h2)); forvar21 = (forvar21 + (1'h1)))
                begin
                  if ($signed((wire8 >= forvar13)))
                    begin
                      reg22 = (-$unsigned(($signed(reg19) ?
                          wire10 : (reg24 ? wire8 : wire10))));
                      reg23 = (reg24 ?
                          (+{{reg21}}) : $unsigned(($unsigned(reg20) ?
                              (~|reg15) : {reg30})));
                    end
                  else
                    begin
                      reg22 = $unsigned((|wire8[(4'h8):(3'h6)]));
                      reg23 = (reg18 >>> forvar13[(3'h6):(3'h4)]);
                      reg24 <= (($unsigned((reg30 | reg15)) & reg28[(2'h3):(1'h0)]) == reg21[(2'h3):(2'h2)]);
                    end
                  if ({(($signed(reg15) != $unsigned(forvar21)) - wire7)})
                    begin
                      reg25 <= (reg21[(1'h0):(1'h0)] >= (reg28[(1'h0):(1'h0)] ?
                          $signed((forvar27 || reg30)) : "0UW349AmQSY"));
                    end
                  else
                    begin
                      reg26 = $unsigned(wire5[(3'h6):(3'h4)]);
                    end
                  for (forvar27 = (1'h0); (forvar27 < (1'h1)); forvar27 = (forvar27 + (1'h1)))
                    begin
                      reg28 = (&("mSx623VB72xXsyY" + reg23));
                      reg31 = reg31[(4'hd):(4'h9)];
                    end
                  reg32 <= reg28;
                end
              if ($unsigned(wire6[(4'h9):(2'h3)]))
                begin
                  reg33 = "79coLc7IyzZ";
                  reg34 = reg31;
                end
              else
                begin
                  if ($unsigned($unsigned("T")))
                    begin
                      reg35 <= ((~&reg18[(2'h3):(2'h2)]) ?
                          $unsigned(($unsigned(reg11) * reg25[(2'h3):(1'h0)])) : forvar26);
                    end
                  else
                    begin
                      reg35 <= (("EaXfYrtXWQE" ?
                              $unsigned(reg34) : wire8[(3'h4):(2'h3)]) ?
                          (("it3YY0y0veqeMOs" > reg31) & ($signed(wire7) + (~forvar13))) : $signed("oMAYT6DaSywQDU"));
                      reg36 <= (8'ha0);
                      reg37 = (($signed("KeFLKWVoXQANlwA") <<< (forvar26[(3'h7):(3'h7)] ?
                          (~&reg20) : (forvar27 ? reg14 : wire5))) >>> reg17);
                    end
                  if (reg29)
                    begin
                      reg38 = ($unsigned(($signed(reg17) ?
                          (&(8'hb0)) : (^~reg37))) ~^ {$signed((reg19 <= reg35))});
                      reg39 = reg36;
                    end
                  else
                    begin
                      reg38 = (^reg36);
                      reg39 = $signed((forvar26[(4'hc):(3'h6)] ?
                          (^~{reg31}) : reg34));
                    end
                  for (forvar40 = (1'h0); (forvar40 < (1'h0)); forvar40 = (forvar40 + (1'h1)))
                    begin
                      reg41 <= ($unsigned("aG") <= "MBzpO");
                      reg42 <= wire6[(4'hc):(2'h2)];
                      reg43 = $signed(reg21[(3'h4):(1'h1)]);
                    end
                end
            end
          if ($unsigned(wire9))
            begin
              for (forvar44 = (1'h0); (forvar44 < (1'h1)); forvar44 = (forvar44 + (1'h1)))
                begin
                  for (forvar45 = (1'h0); (forvar45 < (1'h0)); forvar45 = (forvar45 + (1'h1)))
                    begin
                      reg46 = (~|$signed((reg11 > (reg15 ? reg28 : (8'hb7)))));
                    end
                  if ($unsigned(forvar21))
                    begin
                      reg47 = reg34;
                    end
                  else
                    begin
                      reg47 = $signed((((forvar12 ? reg16 : reg23) ?
                          (reg17 ? (8'hb9) : reg21) : {wire8}) <= reg18));
                      reg48 <= (~&"BLYYKldofgm");
                    end
                  for (forvar49 = (1'h0); (forvar49 < (1'h0)); forvar49 = (forvar49 + (1'h1)))
                    begin
                      reg50 <= wire10[(3'h7):(1'h0)];
                      reg51 <= $unsigned(({((8'haf) & reg11)} ?
                          "O1bERJdxVyeoQ" : (~^(reg15 ? reg26 : reg21))));
                      reg52 = (|$signed(((8'hb9) & reg48[(4'h8):(4'h8)])));
                      reg53 = {$unsigned((&$signed(reg21)))};
                    end
                  for (forvar54 = (1'h0); (forvar54 < (2'h2)); forvar54 = (forvar54 + (1'h1)))
                    begin
                      reg55 = reg34[(1'h0):(1'h0)];
                    end
                end
              for (forvar56 = (1'h0); (forvar56 < (2'h3)); forvar56 = (forvar56 + (1'h1)))
                begin
                  for (forvar57 = (1'h0); (forvar57 < (2'h2)); forvar57 = (forvar57 + (1'h1)))
                    begin
                      reg58 = (8'ha4);
                      reg59 = (forvar13[(3'h5):(1'h0)] ?
                          (^~reg37) : ((forvar44[(3'h5):(1'h1)] ?
                              $unsigned((8'hb7)) : "dhfe") ^ $unsigned({(8'h9c)})));
                      reg60 = $unsigned($unsigned($unsigned((~reg22))));
                    end
                end
            end
          else
            begin
              if (({((forvar49 ? reg32 : reg16) != (forvar56 - wire7))} ?
                  (((forvar40 ^ reg17) == reg37[(4'ha):(4'h9)]) == (reg28[(1'h1):(1'h1)] ?
                      (^(8'h9e)) : (^~reg34))) : "Be6M7CVnPIhzdc"))
                begin
                  reg44 = ({(reg60 ? $signed(reg51) : $signed(reg29))} ?
                      ({$unsigned(reg41)} ?
                          "2pna" : reg25[(3'h7):(3'h6)]) : {(forvar44 << (reg48 ?
                              reg28 : reg25))});
                  for (forvar45 = (1'h0); (forvar45 < (2'h3)); forvar45 = (forvar45 + (1'h1)))
                    begin
                      reg48 <= $unsigned((reg37[(4'h9):(3'h7)] < $unsigned((reg34 ?
                          reg38 : reg41))));
                      reg49 = $unsigned(reg50);
                      reg52 = reg50[(1'h0):(1'h0)];
                    end
                  for (forvar53 = (1'h0); (forvar53 < (2'h2)); forvar53 = (forvar53 + (1'h1)))
                    begin
                      reg54 = {((~|$signed((8'hb9))) >>> $unsigned(reg25[(4'hc):(4'hb)]))};
                      reg55 = reg28[(2'h2):(1'h1)];
                      reg56 <= reg20[(4'h9):(1'h1)];
                    end
                end
              else
                begin
                  reg45 <= reg17[(3'h7):(3'h7)];
                end
              for (forvar57 = (1'h0); (forvar57 < (1'h1)); forvar57 = (forvar57 + (1'h1)))
                begin
                  for (forvar58 = (1'h0); (forvar58 < (1'h0)); forvar58 = (forvar58 + (1'h1)))
                    begin
                      reg59 = ("ixJiknkf" + $signed(reg25));
                      reg60 = wire10[(1'h0):(1'h0)];
                      reg61 <= wire8[(4'h8):(3'h5)];
                      reg62 = $unsigned(reg20);
                    end
                  for (forvar63 = (1'h0); (forvar63 < (1'h1)); forvar63 = (forvar63 + (1'h1)))
                    begin
                      reg64 = ($unsigned($signed(forvar63[(2'h2):(2'h2)])) + (($unsigned(reg50) | (8'had)) ?
                          $unsigned((&forvar40)) : "1nxtF"));
                      reg65 = ("" ? reg38 : reg51);
                      reg66 <= $unsigned(("" ? {$unsigned(reg18)} : "6n"));
                    end
                  for (forvar67 = (1'h0); (forvar67 < (1'h0)); forvar67 = (forvar67 + (1'h1)))
                    begin
                      reg68 <= reg36;
                      reg69 = reg66;
                      reg70 = $unsigned($unsigned($unsigned((reg22 * reg45))));
                      reg71 = ($unsigned("yWc5E") ? "DAi" : $signed((8'haa)));
                    end
                end
            end
        end
      if ($unsigned({{$signed(wire6)}}))
        begin
          if ({($signed(reg36) & ("Dw" >= (reg70 == reg62)))})
            begin
              for (forvar72 = (1'h0); (forvar72 < (1'h0)); forvar72 = (forvar72 + (1'h1)))
                begin
                  if ("eO3dgRQbEtvGT")
                    begin
                      reg73 <= (~$unsigned(reg50[(1'h1):(1'h0)]));
                      reg74 = {(($unsigned(wire7) + (|reg32)) ?
                              "rSwyva" : "wPALD")};
                      reg75 = $signed(reg23[(3'h6):(3'h4)]);
                    end
                  else
                    begin
                      reg73 <= $signed($signed($signed((8'haf))));
                      reg74 = forvar67;
                      reg76 <= {$unsigned(reg62[(1'h0):(1'h0)])};
                      reg77 <= {reg70};
                    end
                  reg78 = ({reg21} ~^ forvar45[(3'h4):(3'h4)]);
                end
            end
          else
            begin
              if ($unsigned(forvar53))
                begin
                  if (($unsigned((^~(wire6 <= reg34))) << "genklxYPKoJ"))
                    begin
                      reg72 = reg23;
                    end
                  else
                    begin
                      reg73 <= $signed(((-reg70) ? reg58 : forvar27));
                      reg76 <= (+"n9swpvxV");
                    end
                  for (forvar77 = (1'h0); (forvar77 < (1'h0)); forvar77 = (forvar77 + (1'h1)))
                    begin
                      reg78 = (&reg38);
                    end
                  reg79 = forvar13[(2'h2):(1'h1)];
                end
              else
                begin
                  for (forvar72 = (1'h0); (forvar72 < (1'h0)); forvar72 = (forvar72 + (1'h1)))
                    begin
                      reg74 = (((!wire6[(2'h3):(1'h0)]) ? (8'hb2) : reg34) ?
                          (reg42[(4'hc):(2'h2)] == reg21) : (|(~|$unsigned(wire9))));
                      reg75 = ($signed($unsigned((reg66 ?
                          reg43 : reg45))) < ($signed((~&forvar53)) != $unsigned((reg58 && reg50))));
                    end
                  if ($signed(($unsigned({forvar12}) ^ reg39)))
                    begin
                      reg76 <= $signed(({(~^reg51)} ?
                          reg47 : ((reg42 >>> reg60) + (forvar72 << forvar45))));
                      reg78 = (~{$unsigned(wire7[(1'h0):(1'h0)])});
                      reg79 = (("Dfu20HvHFi72t" ?
                          (-"zJeiz1NItL") : ((^reg25) ?
                              reg28 : (reg69 >= reg77))) | ($unsigned((reg64 ?
                              forvar67 : forvar54)) ?
                          reg44 : (8'hb9)));
                    end
                  else
                    begin
                      reg76 <= ((~(wire8 << $signed(forvar27))) >>> {{(reg49 <= (8'hac))}});
                      reg78 = wire7[(3'h4):(2'h2)];
                      reg79 = (wire9[(4'h9):(1'h1)] ?
                          reg58 : (reg75[(4'h8):(3'h6)] ?
                              ("TxN2wcXRDUn" ?
                                  reg31 : (reg41 != (8'h9f))) : $signed($signed(reg59))));
                      reg80 = (reg46 ?
                          (reg24[(1'h0):(1'h0)] - forvar40) : (&reg51));
                    end
                  reg81 = (~|("r0Hn" & reg58[(3'h7):(1'h0)]));
                end
            end
          for (forvar82 = (1'h0); (forvar82 < (2'h3)); forvar82 = (forvar82 + (1'h1)))
            begin
              reg83 <= reg46;
              if ((8'hb0))
                begin
                  for (forvar84 = (1'h0); (forvar84 < (1'h1)); forvar84 = (forvar84 + (1'h1)))
                    begin
                      reg85 = (^~$signed(reg74));
                      reg86 = ("EK" ?
                          (({reg60} ?
                              reg60 : reg32) << $signed($signed(reg85))) : $signed(forvar67[(2'h2):(2'h2)]));
                    end
                  for (forvar87 = (1'h0); (forvar87 < (1'h0)); forvar87 = (forvar87 + (1'h1)))
                    begin
                      reg88 = (("k0ZUHqfS7MG" ?
                              "Dua" : $signed($signed((8'hae)))) ?
                          reg24[(1'h1):(1'h1)] : $signed({reg42}));
                      reg89 = forvar57[(3'h4):(1'h0)];
                    end
                  for (forvar90 = (1'h0); (forvar90 < (1'h0)); forvar90 = (forvar90 + (1'h1)))
                    begin
                      reg91 = (!(8'ha3));
                      reg92 = reg78;
                    end
                  for (forvar93 = (1'h0); (forvar93 < (2'h3)); forvar93 = (forvar93 + (1'h1)))
                    begin
                      reg94 <= $unsigned(forvar77[(2'h2):(2'h2)]);
                      reg95 <= (!({(reg50 ? reg14 : reg13)} ?
                          reg66 : $unsigned($signed(reg75))));
                      reg96 <= (^reg11);
                      reg97 <= $signed((((reg71 ^~ reg92) >> $signed((8'ha8))) ?
                          reg20 : $unsigned((wire9 & reg83))));
                    end
                end
              else
                begin
                  if ({"4Yg6Tq"})
                    begin
                      reg84 = ($unsigned(reg45) ^~ reg95[(1'h1):(1'h0)]);
                      reg85 = reg33;
                    end
                  else
                    begin
                      reg87 <= reg31;
                      reg90 <= "fQOPr05DhQlAr";
                      reg93 <= reg87;
                    end
                  for (forvar94 = (1'h0); (forvar94 < (2'h3)); forvar94 = (forvar94 + (1'h1)))
                    begin
                      reg98 = forvar94;
                      reg99 <= (^~(|$signed((reg83 ^ reg13))));
                      reg100 = {(reg18 <= reg92[(3'h4):(2'h2)])};
                    end
                end
            end
          if (($unsigned($unsigned((reg23 ?
              wire9 : reg36))) ^~ (reg95 ~^ "UxDTgY1gbf")))
            begin
              reg101 <= ((~^"TI7") ?
                  $unsigned(reg21[(2'h3):(2'h3)]) : (~^$signed((forvar57 >>> reg38))));
              reg102 <= reg24;
            end
          else
            begin
              reg103 = $signed((reg98 < (reg75 >= "xB")));
              if (wire8)
                begin
                  for (forvar104 = (1'h0); (forvar104 < (2'h3)); forvar104 = (forvar104 + (1'h1)))
                    begin
                      reg105 <= $signed((((~|reg34) ?
                          (reg53 * forvar87) : ((8'ha2) <= forvar72)) <= ($signed(forvar12) ?
                          "krgPqg" : reg70)));
                      reg106 = reg46[(4'h8):(2'h2)];
                      reg107 = "5Rp6QTE3Q";
                    end
                  for (forvar108 = (1'h0); (forvar108 < (2'h2)); forvar108 = (forvar108 + (1'h1)))
                    begin
                      reg109 = $signed(($unsigned((^~reg19)) ?
                          wire8 : ((+forvar58) < (8'hb6))));
                      reg110 = "zXl";
                      reg111 <= {(reg83 >>> ({forvar45} ?
                              reg80 : (reg53 ? reg23 : forvar82)))};
                    end
                end
              else
                begin
                  reg104 = reg75[(4'he):(4'he)];
                  reg106 = $signed(reg46[(3'h7):(3'h6)]);
                  if ($unsigned($signed(reg54)))
                    begin
                      reg108 <= reg90[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg108 <= reg64[(2'h3):(1'h1)];
                      reg111 <= ((~reg65[(1'h1):(1'h0)]) ~^ reg102);
                    end
                  for (forvar112 = (1'h0); (forvar112 < (1'h1)); forvar112 = (forvar112 + (1'h1)))
                    begin
                      reg113 = ($unsigned((|((8'h9f) | reg14))) ?
                          wire7 : (!reg98[(4'hf):(4'he)]));
                      reg114 = $unsigned($unsigned((8'h9c)));
                    end
                end
              reg115 = ("T" ?
                  $unsigned($signed((forvar67 ^~ (8'h9f)))) : reg96[(1'h0):(1'h0)]);
            end
        end
      else
        begin
          if ($unsigned($signed($unsigned($signed(reg52)))))
            begin
              for (forvar72 = (1'h0); (forvar72 < (1'h1)); forvar72 = (forvar72 + (1'h1)))
                begin
                  if ($signed((^~(+reg23[(2'h3):(2'h3)]))))
                    begin
                      reg73 <= "7fC3dpFz3hZvOpn";
                    end
                  else
                    begin
                      reg73 <= $signed({$unsigned(reg89)});
                      reg74 = reg76[(2'h3):(2'h2)];
                      reg75 = ((^~(((8'ha2) && reg55) & forvar12[(4'ha):(3'h7)])) == "a31mxT1Us0PLE");
                    end
                  if (reg55)
                    begin
                      reg78 = reg55[(2'h3):(2'h2)];
                      reg82 <= $signed($signed(((reg102 + reg98) ?
                          reg51[(2'h3):(1'h0)] : reg98)));
                      reg83 <= $unsigned($unsigned({forvar21[(3'h4):(2'h3)]}));
                    end
                  else
                    begin
                      reg78 = forvar57[(1'h1):(1'h1)];
                      reg82 <= reg85[(2'h2):(2'h2)];
                      reg83 <= $signed((("tahvvSd0T7" ?
                          reg65[(1'h0):(1'h0)] : wire9) && forvar44));
                    end
                  for (forvar84 = (1'h0); (forvar84 < (1'h0)); forvar84 = (forvar84 + (1'h1)))
                    begin
                      reg85 = $unsigned("STi4QmT1RM");
                      reg87 <= reg111[(4'he):(4'ha)];
                    end
                end
            end
          else
            begin
              if ("fKmn00gZU2Xf5B3")
                begin
                  if ((($unsigned((^reg18)) << $unsigned((reg59 ?
                      reg48 : reg87))) <= reg96))
                    begin
                      reg72 = $unsigned($unsigned($signed((!reg72))));
                    end
                  else
                    begin
                      reg73 <= ($signed((((8'h9f) ? (8'ha0) : reg34) ?
                              $unsigned(reg75) : {reg98})) ?
                          reg42 : ({(reg30 ?
                                  reg58 : reg83)} <<< $unsigned(reg56)));
                      reg74 = (((forvar53 <= $unsigned(reg54)) <<< (8'h9d)) ?
                          "rY" : (reg30[(2'h2):(1'h0)] >>> (+(reg94 ?
                              reg111 : reg76))));
                      reg75 = (!($unsigned((reg58 ?
                          forvar84 : (8'haa))) <= forvar84));
                      reg78 = reg19[(2'h3):(2'h3)];
                    end
                  reg79 = reg83;
                end
              else
                begin
                  reg73 <= reg80[(2'h3):(1'h0)];
                  if (forvar104)
                    begin
                      reg76 <= ((reg18[(3'h4):(2'h3)] << $unsigned("qv6")) ?
                          (~|$signed((reg61 ?
                              reg104 : wire6))) : $signed(reg52[(1'h0):(1'h0)]));
                      reg78 = {reg32};
                      reg79 = (reg18 >= ($unsigned(forvar27[(1'h1):(1'h1)]) << reg31[(2'h2):(1'h1)]));
                      reg80 = $signed($signed(reg17[(3'h7):(3'h7)]));
                    end
                  else
                    begin
                      reg74 = (^$signed(reg75));
                      reg75 = "S65rtHYlQdUV";
                      reg78 = "pQeA1b2zzK8Uv";
                    end
                  reg81 = {($signed(reg19[(1'h0):(1'h0)]) >> ($signed(reg59) ?
                          reg35[(3'h7):(3'h6)] : (+reg87)))};
                  if ($signed($signed($unsigned((~reg53)))))
                    begin
                      reg84 = (&reg114[(3'h4):(3'h4)]);
                      reg85 = "8yUQILba";
                      reg87 <= $unsigned((($signed((8'hb4)) ?
                              "RAttvWllxlt3f" : (^~reg108)) ?
                          (reg81[(4'he):(1'h1)] ?
                              (forvar108 ?
                                  reg54 : reg89) : (^reg48)) : forvar57[(3'h7):(3'h4)]));
                      reg90 <= (reg91[(2'h3):(2'h2)] <= ($signed(reg25[(4'hc):(4'hc)]) && $signed("KqY3pgFrzP2")));
                    end
                  else
                    begin
                      reg84 = reg51[(4'h9):(1'h1)];
                      reg87 <= ($signed($signed($unsigned(reg11))) ~^ (~&{{reg29}}));
                      reg90 <= forvar49;
                    end
                end
            end
        end
      if ((~|forvar44[(3'h5):(2'h3)]))
        begin
          for (forvar116 = (1'h0); (forvar116 < (2'h3)); forvar116 = (forvar116 + (1'h1)))
            begin
              for (forvar117 = (1'h0); (forvar117 < (2'h2)); forvar117 = (forvar117 + (1'h1)))
                begin
                  reg118 = reg71;
                  if ((reg51[(4'hb):(2'h2)] ?
                      (("aQ1ROrCymh3qi" ^ (reg62 || reg51)) >>> ((^forvar40) ?
                          $signed(wire7) : $unsigned((8'hb0)))) : reg100))
                    begin
                      reg119 <= (~&{(forvar108 ^ $signed(reg35))});
                      reg120 <= {$unsigned((((8'ha0) ^ (8'haf)) ?
                              (+wire10) : (forvar53 != (8'ha0))))};
                    end
                  else
                    begin
                      reg121 = {$signed(reg29)};
                    end
                  for (forvar122 = (1'h0); (forvar122 < (1'h1)); forvar122 = (forvar122 + (1'h1)))
                    begin
                      reg123 = (!(8'hb6));
                      reg124 <= $unsigned((reg23 ? "X3o" : {(+reg71)}));
                      reg125 <= forvar84[(3'h4):(1'h0)];
                      reg126 <= {(!reg119)};
                    end
                end
              for (forvar127 = (1'h0); (forvar127 < (1'h1)); forvar127 = (forvar127 + (1'h1)))
                begin
                  if ({$unsigned($signed((reg76 > reg32)))})
                    begin
                      reg128 <= reg75[(4'hb):(4'ha)];
                      reg129 = $unsigned($unsigned("S50"));
                      reg130 = reg114[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg128 <= $signed($unsigned($unsigned((8'hb9))));
                    end
                end
              for (forvar131 = (1'h0); (forvar131 < (2'h2)); forvar131 = (forvar131 + (1'h1)))
                begin
                  reg132 = "aMJUWRaye";
                  reg133 <= "daez7C32P8";
                  reg134 = (~reg62[(2'h2):(2'h2)]);
                end
              reg135 <= ((~(~^"cRoVmb")) && "odphzK1nu");
            end
          reg136 = reg85;
          reg137 = (reg113[(4'h8):(3'h5)] ? "TWO9Urny6JNCb0" : "t8LJ");
        end
      else
        begin
          for (forvar116 = (1'h0); (forvar116 < (2'h2)); forvar116 = (forvar116 + (1'h1)))
            begin
              for (forvar117 = (1'h0); (forvar117 < (2'h3)); forvar117 = (forvar117 + (1'h1)))
                begin
                  reg118 = wire10;
                end
              if ($unsigned((~^$unsigned($signed((8'hac))))))
                begin
                  if (reg75[(4'h9):(4'h8)])
                    begin
                      reg121 = ($unsigned((reg25[(2'h3):(2'h3)] || (-reg22))) && $signed((forvar12 > (reg119 ?
                          forvar122 : reg43))));
                    end
                  else
                    begin
                      reg119 <= $unsigned($signed(reg13));
                      reg120 <= (((reg39[(3'h7):(1'h0)] ?
                              reg49[(1'h0):(1'h0)] : reg23[(2'h2):(2'h2)]) <= ((reg115 - forvar117) < (reg86 ?
                              reg29 : (8'hb0)))) ?
                          reg109[(3'h4):(3'h4)] : "Wf32qbRCPE25UBk");
                      reg121 = $unsigned((reg20[(3'h4):(2'h2)] ?
                          reg120 : "IRiUkqD7nTe2"));
                    end
                  for (forvar122 = (1'h0); (forvar122 < (2'h3)); forvar122 = (forvar122 + (1'h1)))
                    begin
                      reg123 = $unsigned((reg106[(1'h1):(1'h0)] && forvar82[(1'h0):(1'h0)]));
                      reg124 <= (|(!(8'h9f)));
                      reg125 <= reg115[(4'h9):(2'h3)];
                    end
                  if (forvar72[(3'h4):(1'h1)])
                    begin
                      reg127 = $unsigned(reg86[(1'h0):(1'h0)]);
                      reg129 = (($unsigned(forvar53) ?
                              reg18[(2'h3):(2'h2)] : (8'hb2)) ?
                          (((8'hac) ? "lsxU73ERIeC" : reg69) ?
                              ("5IvYkzuH" & (~^forvar108)) : $unsigned((~|(8'hb7)))) : {(&reg91[(5'h10):(1'h0)])});
                      reg131 <= reg65;
                    end
                  else
                    begin
                      reg127 = reg45[(4'h8):(3'h7)];
                      reg129 = "a6";
                      reg130 = (&$unsigned((reg106[(1'h0):(1'h0)] != $signed(reg125))));
                      reg131 <= "rl9aGv8";
                    end
                  if ((~$unsigned({$unsigned(reg80)})))
                    begin
                      reg132 = "nVS9Jaz9mg03";
                      reg133 <= "GsQW0Szg";
                      reg134 = ((~({forvar63} ?
                          "WBPQQCO" : (reg58 ?
                              reg50 : reg97))) | $signed((((8'hb2) ?
                              reg71 : (8'hae)) ?
                          $unsigned(reg36) : (forvar67 ? reg93 : (8'h9f)))));
                    end
                  else
                    begin
                      reg133 <= {reg82};
                      reg134 = $unsigned($signed(reg25));
                      reg136 = $unsigned({forvar49});
                    end
                end
              else
                begin
                  for (forvar119 = (1'h0); (forvar119 < (2'h3)); forvar119 = (forvar119 + (1'h1)))
                    begin
                      reg120 <= (reg130[(1'h0):(1'h0)] ?
                          "ICSx" : (~(^(reg15 ? reg88 : reg90))));
                      reg121 = $signed(reg73);
                      reg122 <= (forvar119[(2'h3):(1'h1)] ^ $unsigned(reg33));
                      reg123 = "sHViq";
                    end
                  if ($signed(forvar58[(3'h5):(2'h2)]))
                    begin
                      reg127 = "6";
                      reg129 = {reg92[(3'h6):(2'h2)]};
                    end
                  else
                    begin
                      reg127 = $signed(reg135[(3'h4):(2'h2)]);
                      reg129 = (~{$unsigned(reg84[(3'h5):(1'h0)])});
                    end
                  reg130 = (!(~|($unsigned(forvar57) ?
                      {reg58} : $unsigned(reg84))));
                  reg132 = $unsigned($unsigned({(~|reg94)}));
                end
              reg138 <= reg69[(1'h1):(1'h0)];
            end
        end
      for (forvar139 = (1'h0); (forvar139 < (1'h1)); forvar139 = (forvar139 + (1'h1)))
        begin
          for (forvar140 = (1'h0); (forvar140 < (1'h0)); forvar140 = (forvar140 + (1'h1)))
            begin
              reg141 <= "49nncQr";
              for (forvar142 = (1'h0); (forvar142 < (1'h0)); forvar142 = (forvar142 + (1'h1)))
                begin
                  for (forvar143 = (1'h0); (forvar143 < (1'h1)); forvar143 = (forvar143 + (1'h1)))
                    begin
                      reg144 = forvar72[(3'h4):(3'h4)];
                      reg145 <= reg35;
                    end
                  reg146 = (!reg46[(2'h3):(2'h2)]);
                  if (({"8NGESpKDHS6vBmP"} ? (8'hb2) : "q"))
                    begin
                      reg147 <= {({(reg95 ?
                                  reg49 : reg114)} && {$signed((8'hab))})};
                      reg148 <= ($unsigned($unsigned(reg30)) ?
                          (^~(8'h9e)) : reg44[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg147 <= "mmnXAL6MSSCm";
                      reg148 <= "qCppG7vv9PJx9";
                    end
                end
              for (forvar149 = (1'h0); (forvar149 < (1'h1)); forvar149 = (forvar149 + (1'h1)))
                begin
                  for (forvar150 = (1'h0); (forvar150 < (1'h0)); forvar150 = (forvar150 + (1'h1)))
                    begin
                      reg151 = "7yOV";
                    end
                  reg152 = $unsigned(("lPw" ~^ ("1LUbRySSF3I" << {forvar142})));
                  reg153 = reg26[(1'h1):(1'h1)];
                end
              reg154 <= forvar54[(4'ha):(1'h0)];
            end
          for (forvar155 = (1'h0); (forvar155 < (1'h0)); forvar155 = (forvar155 + (1'h1)))
            begin
              reg156 = forvar84;
              for (forvar157 = (1'h0); (forvar157 < (2'h2)); forvar157 = (forvar157 + (1'h1)))
                begin
                  reg158 <= (((|{reg114}) - wire9) ?
                      (((reg14 ?
                          reg36 : reg55) << reg94) ^ $signed((-forvar54))) : reg113);
                end
              if (reg70)
                begin
                  reg159 = (~&$signed(wire7));
                  reg160 <= $signed($signed({$signed(reg115)}));
                  for (forvar161 = (1'h0); (forvar161 < (2'h3)); forvar161 = (forvar161 + (1'h1)))
                    begin
                      reg162 <= forvar49[(1'h0):(1'h0)];
                      reg163 = $signed({($unsigned(reg106) || reg95[(3'h4):(3'h4)])});
                      reg164 = ($unsigned((&(~|reg35))) ^~ reg46);
                    end
                  for (forvar165 = (1'h0); (forvar165 < (1'h0)); forvar165 = (forvar165 + (1'h1)))
                    begin
                      reg166 = ({reg41} && $signed(({reg141} + "YGCZc")));
                    end
                end
              else
                begin
                  reg159 = $signed(reg160);
                  reg160 <= $unsigned(($unsigned((reg138 & (8'hb3))) ?
                      $unsigned((reg33 ? reg152 : reg105)) : $signed({reg29})));
                  reg161 <= $signed("6g2tCw");
                end
              if ((8'hb9))
                begin
                  for (forvar167 = (1'h0); (forvar167 < (2'h2)); forvar167 = (forvar167 + (1'h1)))
                    begin
                      reg168 = $signed(reg159[(3'h4):(3'h4)]);
                      reg169 <= (8'h9c);
                      reg170 <= "t4icpYcKKpGotN";
                      reg171 <= "DaAl4nf09w3c";
                    end
                  for (forvar172 = (1'h0); (forvar172 < (1'h0)); forvar172 = (forvar172 + (1'h1)))
                    begin
                      reg173 = $signed((reg128 ?
                          ($signed(reg79) < (reg132 ^~ forvar155)) : ("q6oJsUhyDyzyfD" ?
                              "3Etd" : $signed(reg20))));
                      reg174 = (~|(8'ha3));
                      reg175 = (~"mOnhmxz");
                      reg176 <= (((^~(reg168 ^~ (8'ha0))) <<< reg120) ?
                          forvar112[(1'h0):(1'h0)] : forvar87);
                    end
                  for (forvar177 = (1'h0); (forvar177 < (1'h0)); forvar177 = (forvar177 + (1'h1)))
                    begin
                      reg178 = ((((reg118 ? (8'hb6) : reg69) & reg54) ?
                          $signed($unsigned(forvar82)) : (!((8'ha7) ?
                              reg71 : reg105))) ~^ reg20[(3'h6):(1'h0)]);
                      reg179 <= ({reg90} ? wire9 : $signed(("F" < {(8'hb5)})));
                      reg180 = reg45;
                    end
                end
              else
                begin
                  if ((!reg103))
                    begin
                      reg167 = reg26[(1'h0):(1'h0)];
                      reg169 <= $signed({forvar172});
                      reg170 <= (($unsigned((8'h9c)) <= (reg38[(3'h4):(2'h3)] ?
                          ((8'hb5) ?
                              reg73 : forvar56) : $unsigned(reg37))) <<< $signed((reg22[(1'h1):(1'h0)] && $unsigned(reg77))));
                      reg172 = (~^reg152);
                    end
                  else
                    begin
                      reg167 = (^reg99);
                      reg169 <= reg64[(3'h5):(1'h0)];
                    end
                  for (forvar173 = (1'h0); (forvar173 < (1'h0)); forvar173 = (forvar173 + (1'h1)))
                    begin
                      reg174 = {reg69[(2'h2):(1'h0)]};
                    end
                  for (forvar175 = (1'h0); (forvar175 < (2'h2)); forvar175 = (forvar175 + (1'h1)))
                    begin
                      reg176 <= reg171;
                      reg177 = reg30[(4'hc):(4'h8)];
                    end
                  for (forvar178 = (1'h0); (forvar178 < (2'h2)); forvar178 = (forvar178 + (1'h1)))
                    begin
                      reg180 = wire9;
                      reg181 = ($signed(forvar26[(4'h9):(3'h6)]) <<< reg58);
                      reg182 <= $signed($unsigned($unsigned(reg39)));
                    end
                end
            end
          for (forvar183 = (1'h0); (forvar183 < (1'h1)); forvar183 = (forvar183 + (1'h1)))
            begin
              if ($signed($signed(($signed(forvar94) ~^ reg56[(3'h5):(3'h4)]))))
                begin
                  for (forvar184 = (1'h0); (forvar184 < (1'h0)); forvar184 = (forvar184 + (1'h1)))
                    begin
                      reg185 = "b";
                      reg186 = $unsigned($unsigned("IE5d8v2kf"));
                      reg187 <= $signed((reg147 != (~|$signed(reg162))));
                    end
                  reg188 = ($unsigned(reg61[(3'h6):(2'h3)]) ?
                      $signed(($signed(reg73) ?
                          (forvar72 ?
                              forvar45 : forvar26) : $unsigned(reg75))) : (^~((+wire10) ^ (reg109 ?
                          reg131 : reg95))));
                end
              else
                begin
                  if (($unsigned("oTNA41CNl") > ($signed((reg102 ?
                      (8'ha6) : reg81)) >>> $signed((reg128 != reg174)))))
                    begin
                      reg184 = reg167[(3'h7):(3'h6)];
                      reg187 <= {forvar112[(2'h3):(1'h0)]};
                    end
                  else
                    begin
                      reg187 <= reg134[(4'hb):(2'h2)];
                      reg188 = $signed(({((8'hb4) + forvar131)} ?
                          $signed((reg172 ? forvar26 : reg96)) : reg49));
                    end
                  reg189 = (&(({(8'ha3)} ? reg161[(1'h0):(1'h0)] : reg138) ?
                      "JwEZ" : forvar119));
                  for (forvar190 = (1'h0); (forvar190 < (1'h1)); forvar190 = (forvar190 + (1'h1)))
                    begin
                      reg191 = $unsigned($signed($unsigned((^(8'ha9)))));
                      reg192 = $unsigned(reg114[(2'h2):(2'h2)]);
                      reg193 = $unsigned((~&forvar142[(3'h6):(3'h6)]));
                      reg194 = reg138[(3'h7):(1'h1)];
                    end
                end
              for (forvar195 = (1'h0); (forvar195 < (1'h1)); forvar195 = (forvar195 + (1'h1)))
                begin
                  for (forvar196 = (1'h0); (forvar196 < (2'h3)); forvar196 = (forvar196 + (1'h1)))
                    begin
                      reg197 = (forvar49[(4'hb):(2'h3)] | (~|((forvar150 ?
                              reg171 : reg42) ?
                          reg137[(2'h3):(2'h2)] : $signed(reg174))));
                    end
                  reg198 = (reg197[(1'h1):(1'h1)] ?
                      (8'hab) : $signed(reg161[(1'h0):(1'h0)]));
                  if ($signed(($signed(reg175) ?
                      (reg53 ?
                          $signed((8'hb9)) : $unsigned(forvar49)) : $signed((+reg198)))))
                    begin
                      reg199 <= (("FW" ^~ (|$unsigned(reg21))) + ($unsigned((reg121 || reg79)) ?
                          {$unsigned(reg105)} : (&(~^reg77))));
                      reg200 = (~($unsigned((~&reg49)) >>> $signed((forvar167 >> wire10))));
                      reg201 = forvar117;
                      reg202 = $signed(reg77[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg199 <= "F";
                    end
                  for (forvar203 = (1'h0); (forvar203 < (1'h1)); forvar203 = (forvar203 + (1'h1)))
                    begin
                      reg204 <= $unsigned(({reg33[(3'h7):(1'h0)]} >> $signed($signed(forvar44))));
                      reg205 = (~&(($unsigned((8'hab)) == $unsigned(reg122)) >>> reg15));
                      reg206 = "HJvRivssHR7oh7";
                    end
                end
              if ((reg185[(4'hc):(2'h3)] ?
                  {(reg129 ? (8'hae) : {(8'hb3)})} : "O"))
                begin
                  for (forvar207 = (1'h0); (forvar207 < (1'h0)); forvar207 = (forvar207 + (1'h1)))
                    begin
                      reg208 <= forvar87;
                      reg209 = "D7SBe3";
                      reg210 = (~^(~^"azS4VL"));
                      reg211 <= ($unsigned("VepcJloHTPV5m") ?
                          (reg78[(1'h0):(1'h0)] > (&(^reg105))) : ($signed(wire8) >= (!(|reg88))));
                    end
                end
              else
                begin
                  for (forvar207 = (1'h0); (forvar207 < (1'h0)); forvar207 = (forvar207 + (1'h1)))
                    begin
                      reg208 <= reg158[(3'h5):(2'h2)];
                    end
                  reg209 = (~^(((reg119 >>> reg113) ?
                      $signed(reg173) : (forvar183 + reg87)) | $unsigned((reg78 ?
                      (8'h9e) : reg154))));
                  if ($unsigned({((reg84 ? forvar131 : reg130) - (reg153 ?
                          reg89 : reg22))}))
                    begin
                      reg210 = $unsigned({((forvar157 && reg126) & (~|reg34))});
                      reg211 <= ("" ?
                          ($signed((reg181 ?
                              forvar84 : reg65)) < ($unsigned(reg186) <<< $unsigned(forvar94))) : wire6);
                      reg212 = {(($signed(reg75) ?
                                  $signed((8'hb1)) : "eop3cOYh5qKXxd") ?
                              reg28[(2'h3):(1'h1)] : (~&forvar117))};
                      reg213 = (((forvar184 ?
                          (-forvar87) : $signed((8'hb7))) < $unsigned((reg31 == reg192))) >> {forvar143[(2'h2):(1'h0)]});
                    end
                  else
                    begin
                      reg210 = (~|$signed(reg101[(3'h7):(1'h0)]));
                    end
                end
            end
        end
    end
  module214 #() modinst2023 (wire2022, clk, reg124, reg126, reg14, reg102, reg141);
  assign wire2024 = $unsigned(($unsigned("W2wxZI") ?
                        reg126 : (^~(reg158 ? reg36 : reg101))));
  assign wire2025 = $signed("");
  always
    @(posedge clk) begin
      for (forvar2026 = (1'h0); (forvar2026 < (1'h1)); forvar2026 = (forvar2026 + (1'h1)))
        begin
          reg2027 = "";
          for (forvar2028 = (1'h0); (forvar2028 < (2'h2)); forvar2028 = (forvar2028 + (1'h1)))
            begin
              for (forvar2029 = (1'h0); (forvar2029 < (1'h0)); forvar2029 = (forvar2029 + (1'h1)))
                begin
                  reg2030 <= ((~$signed((reg158 << wire2024))) ?
                      (&reg147) : reg19);
                  reg2031 = ($unsigned({reg102}) >> $signed("hTlhKKwV"));
                  for (forvar2032 = (1'h0); (forvar2032 < (1'h1)); forvar2032 = (forvar2032 + (1'h1)))
                    begin
                      reg2033 = (~|$signed($signed((^wire10))));
                      reg2034 = (~|reg161);
                      reg2035 = $unsigned(((reg102[(4'hc):(4'hc)] ?
                              $signed(reg111) : (reg96 ? (8'ha4) : reg61)) ?
                          reg2030[(2'h3):(2'h2)] : reg41[(2'h2):(1'h1)]));
                    end
                  reg2036 = reg161[(1'h0):(1'h0)];
                end
              for (forvar2037 = (1'h0); (forvar2037 < (1'h1)); forvar2037 = (forvar2037 + (1'h1)))
                begin
                  reg2038 = (^~reg29[(3'h5):(3'h4)]);
                  reg2039 <= ({("iyRneKH" ?
                          "IymtLCo9WmbcaGL" : ((8'h9f) + reg179))} | {"aB2vBLOt3oKDPHv"});
                  for (forvar2040 = (1'h0); (forvar2040 < (1'h1)); forvar2040 = (forvar2040 + (1'h1)))
                    begin
                      reg2041 = reg2031[(2'h2):(1'h0)];
                      reg2042 <= ($unsigned(reg42[(3'h4):(2'h2)]) ?
                          reg42 : {(reg2039 >>> (reg42 * reg141))});
                      reg2043 <= "zIf4zVmxwMpbhr0";
                      reg2044 = $signed((($signed(reg147) ?
                          {reg51} : reg138[(4'h8):(3'h6)]) + $unsigned({reg204})));
                    end
                  for (forvar2045 = (1'h0); (forvar2045 < (1'h0)); forvar2045 = (forvar2045 + (1'h1)))
                    begin
                      reg2046 = reg102;
                      reg2047 = reg50[(2'h2):(1'h0)];
                      reg2048 = "POhya";
                    end
                end
            end
        end
      for (forvar2049 = (1'h0); (forvar2049 < (1'h1)); forvar2049 = (forvar2049 + (1'h1)))
        begin
          for (forvar2050 = (1'h0); (forvar2050 < (1'h0)); forvar2050 = (forvar2050 + (1'h1)))
            begin
              reg2051 <= {($signed(reg97) | (((8'ha3) << reg30) | (reg24 - reg171)))};
              reg2052 = reg2051[(1'h0):(1'h0)];
            end
          for (forvar2053 = (1'h0); (forvar2053 < (1'h1)); forvar2053 = (forvar2053 + (1'h1)))
            begin
              reg2054 <= {((~^$signed(forvar2053)) || (+reg21[(2'h2):(1'h1)]))};
              for (forvar2055 = (1'h0); (forvar2055 < (1'h1)); forvar2055 = (forvar2055 + (1'h1)))
                begin
                  reg2056 <= {$unsigned($signed((reg41 ? (8'ha3) : reg42)))};
                  for (forvar2057 = (1'h0); (forvar2057 < (1'h1)); forvar2057 = (forvar2057 + (1'h1)))
                    begin
                      reg2058 = "bHUZJ";
                      reg2059 <= reg2056[(3'h4):(2'h2)];
                      reg2060 <= ($signed(($signed(reg77) > ((8'hb2) ^~ reg83))) ?
                          wire10[(3'h7):(1'h0)] : (~{$unsigned(reg176)}));
                      reg2061 = (~&$unsigned((8'hb1)));
                    end
                end
              if ("2HnhW")
                begin
                  for (forvar2062 = (1'h0); (forvar2062 < (1'h1)); forvar2062 = (forvar2062 + (1'h1)))
                    begin
                      reg2063 = reg126[(3'h4):(2'h3)];
                      reg2064 = reg2041;
                      reg2065 <= $signed((~^"nnqAVOyltO"));
                      reg2066 = (~|reg125[(3'h6):(1'h0)]);
                    end
                  reg2067 = reg131[(1'h1):(1'h1)];
                  reg2068 <= (((^~reg128) ?
                      ($unsigned(reg2052) << (reg182 < forvar2028)) : (!$unsigned(reg2043))) >> (({reg122} ?
                          forvar2037 : {forvar2032}) ?
                      ($signed(reg2039) ?
                          $signed(reg128) : (reg2060 ?
                              reg77 : forvar2053)) : $unsigned($unsigned(reg2052))));
                  for (forvar2069 = (1'h0); (forvar2069 < (1'h1)); forvar2069 = (forvar2069 + (1'h1)))
                    begin
                      reg2070 = "xQNha8v";
                    end
                end
              else
                begin
                  reg2062 = $unsigned(forvar2057[(3'h4):(1'h1)]);
                  for (forvar2063 = (1'h0); (forvar2063 < (2'h2)); forvar2063 = (forvar2063 + (1'h1)))
                    begin
                      reg2064 = (($signed("hBKKDNxELH9N") ^ reg2065[(2'h3):(1'h0)]) ?
                          (((+reg2059) ?
                              (~^wire9) : $unsigned(reg73)) != ((8'hb5) ?
                              {wire2024} : $signed(reg2063))) : forvar2029[(2'h3):(2'h3)]);
                    end
                end
              reg2071 = $unsigned((~^{forvar2029}));
            end
          reg2072 <= $unsigned($signed({(~reg51)}));
        end
      for (forvar2073 = (1'h0); (forvar2073 < (1'h1)); forvar2073 = (forvar2073 + (1'h1)))
        begin
          reg2074 <= reg131;
          if (($signed((&(reg41 ? wire2024 : wire7))) ? reg48 : (8'h9c)))
            begin
              if ($signed((((reg126 <= reg2071) ?
                      (reg2059 ?
                          (8'ha5) : forvar2026) : reg2070[(4'h9):(1'h1)]) ?
                  ((~^forvar2057) >> $unsigned((8'hac))) : {reg176})))
                begin
                  reg2075 = $signed(reg32[(3'h5):(3'h5)]);
                end
              else
                begin
                  if (($signed($unsigned(reg131)) ?
                      (8'hb6) : $signed($unsigned((~^reg161)))))
                    begin
                      reg2075 = ($signed(((forvar2049 >> reg211) <<< $unsigned((8'hb3)))) ?
                          $signed("ZgwRf496EkTO") : (!reg30));
                      reg2076 = reg160[(2'h2):(1'h1)];
                      reg2077 = $signed(wire6[(4'h9):(1'h1)]);
                      reg2078 = $unsigned((-("f2odavJnfvmQBO9" ?
                          $signed(wire7) : reg2035[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg2079 <= $signed("");
                      reg2080 = reg73[(3'h4):(2'h2)];
                      reg2081 = (|reg148);
                    end
                end
              if (reg61[(1'h1):(1'h0)])
                begin
                  for (forvar2082 = (1'h0); (forvar2082 < (1'h1)); forvar2082 = (forvar2082 + (1'h1)))
                    begin
                      reg2083 = $unsigned(reg2046[(3'h7):(3'h7)]);
                      reg2084 = (($signed((wire2022 ?
                              forvar2055 : reg2068)) & $signed($signed(reg211))) ?
                          ({((8'hb5) ?
                                  reg2061 : reg171)} == reg2063[(3'h6):(1'h1)]) : (^reg2052));
                      reg2085 <= $signed((&reg95));
                      reg2086 = ($signed((^(8'ha6))) | wire6[(4'ha):(4'ha)]);
                    end
                  for (forvar2087 = (1'h0); (forvar2087 < (2'h3)); forvar2087 = (forvar2087 + (1'h1)))
                    begin
                      reg2088 = {reg2064};
                      reg2089 = $signed((~&$unsigned("XJkhycN5chI")));
                      reg2090 <= (reg2067 ?
                          forvar2062[(1'h0):(1'h0)] : (^~reg2079));
                    end
                  for (forvar2091 = (1'h0); (forvar2091 < (1'h1)); forvar2091 = (forvar2091 + (1'h1)))
                    begin
                      reg2092 = (forvar2029 ?
                          reg2066[(2'h3):(2'h2)] : $signed($signed(reg42[(4'hd):(4'hd)])));
                      reg2093 = "mqHGIuX1vnHlEq1";
                      reg2094 = forvar2069[(2'h2):(1'h0)];
                      reg2095 <= $unsigned((8'ha2));
                    end
                end
              else
                begin
                  if (forvar2040[(1'h0):(1'h0)])
                    begin
                      reg2082 = {($signed($signed(reg145)) * reg138[(4'ha):(4'ha)])};
                      reg2085 <= $signed(wire5[(2'h2):(1'h1)]);
                      reg2086 = (((reg187[(4'ha):(3'h7)] ?
                          (~&forvar2062) : reg2034[(4'hb):(4'h9)]) <= (~(^~reg2051))) | reg2031);
                      reg2087 = (8'hb7);
                    end
                  else
                    begin
                      reg2082 = $unsigned((($unsigned(reg77) ?
                              ((8'ha1) ?
                                  reg2089 : reg131) : reg2086[(3'h4):(2'h3)]) ?
                          (reg2067[(2'h3):(1'h1)] ?
                              reg102 : $signed(reg2042)) : {((8'hb0) ?
                                  reg122 : reg45)}));
                      reg2085 <= {(reg2095[(3'h7):(3'h5)] ^~ $unsigned(reg124))};
                    end
                  reg2088 = reg68[(4'hc):(2'h3)];
                  reg2089 = (!$signed(forvar2057[(2'h2):(1'h1)]));
                  reg2091 = "zq";
                end
              reg2096 = (&{(^~(8'ha8))});
            end
          else
            begin
              for (forvar2075 = (1'h0); (forvar2075 < (1'h0)); forvar2075 = (forvar2075 + (1'h1)))
                begin
                  for (forvar2076 = (1'h0); (forvar2076 < (1'h1)); forvar2076 = (forvar2076 + (1'h1)))
                    begin
                      reg2077 = $signed((|$unsigned((+reg187))));
                      reg2078 = $signed(("P9bP0v" ?
                          (reg73[(2'h2):(2'h2)] ?
                              (reg2083 >> wire2024) : $unsigned(reg135)) : reg126));
                    end
                  if ($unsigned(((^~reg2085[(1'h0):(1'h0)]) ?
                      (reg32[(3'h5):(2'h3)] == ((8'h9e) ?
                          (8'ha2) : reg2072)) : reg122[(2'h3):(2'h3)])))
                    begin
                      reg2080 = $unsigned(reg2078);
                      reg2085 <= ($signed((reg2080[(2'h3):(1'h0)] ?
                              "4T" : forvar2087[(4'ha):(4'h8)])) ?
                          $unsigned(((forvar2037 ? reg76 : forvar2063) ?
                              reg111 : reg124[(3'h6):(1'h1)])) : {({forvar2057} ?
                                  (reg95 <= reg24) : reg160[(2'h3):(2'h3)])});
                    end
                  else
                    begin
                      reg2079 <= $signed({{$unsigned(reg50)}});
                      reg2080 = ($unsigned(((reg24 < forvar2049) ^~ (reg95 != forvar2063))) ^ ("5AtRT1CqkpitW" && $signed((reg82 >> wire2024))));
                      reg2085 <= reg131[(4'h8):(4'h8)];
                    end
                  reg2086 = (^~(((~^reg169) <= reg20) ?
                      ("P02mSk" ?
                          reg111[(3'h5):(3'h4)] : (^~reg2085)) : (|(reg42 ?
                          reg20 : wire9))));
                end
              reg2090 <= ($signed(reg97[(3'h7):(2'h3)]) ?
                  $signed(reg133) : reg2063[(4'he):(2'h3)]);
            end
          reg2097 <= (("WabWUVA3S3" >= (!forvar2063[(3'h5):(3'h4)])) > reg145[(3'h4):(3'h4)]);
          reg2098 <= reg2096;
        end
    end
  module358 #() modinst2100 (.wire361(reg147), .wire359(reg102), .wire363(reg176), .wire360(reg182), .clk(clk), .wire362(reg199), .y(wire2099));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module214  (y, clk, wire215, wire216, wire217, wire218, wire219);
  output wire [(32'h40e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire215;
  input wire [(4'hc):(1'h0)] wire216;
  input wire [(4'hf):(1'h0)] wire217;
  input wire [(4'he):(1'h0)] wire218;
  input wire signed [(3'h7):(1'h0)] wire219;
  wire signed [(2'h2):(1'h0)] wire2021;
  wire [(3'h6):(1'h0)] wire2020;
  wire [(3'h4):(1'h0)] wire220;
  wire signed [(4'he):(1'h0)] wire274;
  wire [(4'ha):(1'h0)] wire1977;
  reg signed [(4'ha):(1'h0)] reg2016 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2012 = (1'h0);
  reg [(5'h10):(1'h0)] reg2006 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2004 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2003 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2002 = (1'h0);
  reg [(4'h9):(1'h0)] reg2000 = (1'h0);
  reg [(5'h10):(1'h0)] reg1996 = (1'h0);
  reg [(2'h2):(1'h0)] reg1995 = (1'h0);
  reg [(4'hf):(1'h0)] reg1986 = (1'h0);
  reg [(4'h8):(1'h0)] reg225 = (1'h0);
  reg [(4'h9):(1'h0)] reg227 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg229 = (1'h0);
  reg [(5'h10):(1'h0)] reg230 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg231 = (1'h0);
  reg [(4'ha):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg248 = (1'h0);
  reg [(4'hf):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg252 = (1'h0);
  reg [(4'hc):(1'h0)] reg254 = (1'h0);
  reg [(4'ha):(1'h0)] reg259 = (1'h0);
  reg signed [(4'he):(1'h0)] reg260 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg262 = (1'h0);
  reg [(4'hd):(1'h0)] reg263 = (1'h0);
  reg [(3'h5):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg265 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg267 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg270 = (1'h0);
  reg [(4'ha):(1'h0)] reg246 = (1'h0);
  reg [(4'h8):(1'h0)] reg257 = (1'h0);
  reg [(3'h4):(1'h0)] reg272 = (1'h0);
  reg [(4'h8):(1'h0)] reg2019 = (1'h0);
  reg [(4'hb):(1'h0)] reg2018 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2017 = (1'h0);
  reg [(3'h5):(1'h0)] reg1982 = (1'h0);
  reg [(3'h4):(1'h0)] reg1981 = (1'h0);
  reg [(4'hf):(1'h0)] reg2015 = (1'h0);
  reg [(4'h9):(1'h0)] reg2014 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2013 = (1'h0);
  reg [(2'h2):(1'h0)] reg2011 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2010 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2009 = (1'h0);
  reg [(4'hf):(1'h0)] reg2008 = (1'h0);
  reg [(5'h10):(1'h0)] reg2007 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2005 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2001 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1999 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1998 = (1'h0);
  reg [(4'hb):(1'h0)] reg1997 = (1'h0);
  reg [(4'he):(1'h0)] reg1994 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1993 = (1'h0);
  reg [(3'h6):(1'h0)] reg1992 = (1'h0);
  reg [(2'h3):(1'h0)] reg1991 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1990 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1989 = (1'h0);
  reg [(5'h10):(1'h0)] reg1988 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1987 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1985 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1984 = (1'h0);
  reg [(3'h6):(1'h0)] reg1983 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1982 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1981 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1980 = (1'h0);
  reg [(4'hc):(1'h0)] reg1979 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg273 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg269 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar268 = (1'h0);
  reg [(2'h3):(1'h0)] forvar250 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg253 = (1'h0);
  reg [(3'h5):(1'h0)] reg245 = (1'h0);
  reg [(3'h7):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg271 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar269 = (1'h0);
  reg [(5'h10):(1'h0)] reg268 = (1'h0);
  reg [(2'h3):(1'h0)] reg266 = (1'h0);
  reg [(4'he):(1'h0)] reg261 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar258 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar257 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg256 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg255 = (1'h0);
  reg [(2'h2):(1'h0)] forvar253 = (1'h0);
  reg [(3'h7):(1'h0)] reg251 = (1'h0);
  reg [(4'he):(1'h0)] reg249 = (1'h0);
  reg [(4'he):(1'h0)] reg247 = (1'h0);
  reg [(3'h4):(1'h0)] forvar246 = (1'h0);
  reg [(2'h2):(1'h0)] forvar245 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg244 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg243 = (1'h0);
  reg [(4'hf):(1'h0)] forvar242 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg241 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg240 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg239 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg238 = (1'h0);
  reg [(4'h8):(1'h0)] reg237 = (1'h0);
  reg [(4'hc):(1'h0)] forvar236 = (1'h0);
  reg signed [(4'he):(1'h0)] reg234 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar233 = (1'h0);
  reg [(4'h8):(1'h0)] forvar232 = (1'h0);
  reg [(3'h7):(1'h0)] reg228 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg226 = (1'h0);
  reg [(4'h9):(1'h0)] forvar224 = (1'h0);
  reg [(3'h6):(1'h0)] forvar223 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar222 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar221 = (1'h0);
  assign y = {wire2021,
                 reg2003,
                 reg2002,
                 reg2000,
                 reg235,
                 reg252,
                 reg263,
                 reg267,
                 reg270,
                 reg2019,
                 reg2011,
                 reg2008,
                 reg2007,
                 forvar1998,
                 reg1992,
                 forvar1989,
                 reg1988,
                 forvar1982,
                 reg245,
                 reg242,
                 reg261,
                 forvar258,
                 forvar257,
                 forvar253,
                 reg251,
                 reg249,
                 reg247,
                 forvar246,
                 reg243,
                 forvar242,
                 reg240,
                 forvar236,
                 forvar233,
                 reg228,
                 forvar224,
                 (1'h0)};
  assign wire220 = $signed(wire215);
  always
    @(posedge clk) begin
      for (forvar221 = (1'h0); (forvar221 < (2'h3)); forvar221 = (forvar221 + (1'h1)))
        begin
          for (forvar222 = (1'h0); (forvar222 < (1'h0)); forvar222 = (forvar222 + (1'h1)))
            begin
              for (forvar223 = (1'h0); (forvar223 < (2'h2)); forvar223 = (forvar223 + (1'h1)))
                begin
                  for (forvar224 = (1'h0); (forvar224 < (2'h2)); forvar224 = (forvar224 + (1'h1)))
                    begin
                      reg225 <= $unsigned((wire218 ?
                          wire219 : ((forvar221 * wire220) ?
                              (+forvar224) : (forvar224 ?
                                  wire220 : forvar221))));
                      reg226 = $unsigned(reg225);
                    end
                  if ($signed(((8'hb3) != (~wire219[(3'h6):(1'h0)]))))
                    begin
                      reg227 <= wire218[(1'h1):(1'h0)];
                      reg228 = $unsigned((("KHI" <<< (&reg225)) ?
                          $signed((forvar221 ?
                              (8'ha8) : reg226)) : wire215[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg228 = (($unsigned(wire219) <<< wire215) ?
                          wire220[(1'h1):(1'h1)] : $signed(forvar221));
                      reg229 <= reg227[(1'h0):(1'h0)];
                      reg230 <= reg227;
                      reg231 <= $unsigned(({(^~reg229)} ?
                          (~(&(8'hba))) : ((|reg227) ? reg226 : forvar222)));
                    end
                end
              for (forvar232 = (1'h0); (forvar232 < (2'h2)); forvar232 = (forvar232 + (1'h1)))
                begin
                  for (forvar233 = (1'h0); (forvar233 < (2'h3)); forvar233 = (forvar233 + (1'h1)))
                    begin
                      reg234 = ($signed($unsigned((wire217 ?
                              reg227 : reg230))) ?
                          wire215 : "oh1EYwEh");
                      reg235 <= $unsigned($unsigned({reg226[(4'hb):(3'h6)]}));
                    end
                  for (forvar236 = (1'h0); (forvar236 < (1'h1)); forvar236 = (forvar236 + (1'h1)))
                    begin
                      reg237 = wire216[(4'hb):(3'h6)];
                      reg238 = $unsigned({(reg228[(1'h0):(1'h0)] <<< (reg225 - (8'haf)))});
                      reg239 = $unsigned(reg238);
                    end
                  if (forvar232)
                    begin
                      reg240 = {reg238[(3'h7):(3'h7)]};
                    end
                  else
                    begin
                      reg240 = reg239;
                      reg241 = (~&(((forvar236 ?
                              reg235 : reg227) ^ (~|reg225)) ?
                          ("cVdqTVDm" ?
                              reg230[(4'hf):(2'h2)] : forvar232[(4'h8):(1'h1)]) : $signed({forvar233})));
                    end
                end
            end
          if (((|$signed($unsigned(wire216))) ?
              {$signed($signed(reg229))} : reg231[(3'h7):(1'h1)]))
            begin
              for (forvar242 = (1'h0); (forvar242 < (1'h0)); forvar242 = (forvar242 + (1'h1)))
                begin
                  reg243 = ("pbpaEgCXU4" ?
                      reg231[(4'hb):(1'h0)] : reg235[(3'h6):(3'h5)]);
                end
              reg244 = (&"TytVFA03eQBLiav");
              for (forvar245 = (1'h0); (forvar245 < (2'h3)); forvar245 = (forvar245 + (1'h1)))
                begin
                  for (forvar246 = (1'h0); (forvar246 < (1'h0)); forvar246 = (forvar246 + (1'h1)))
                    begin
                      reg247 = wire218[(1'h0):(1'h0)];
                    end
                  if ({$unsigned(({reg243} > "y"))})
                    begin
                      reg248 <= reg241[(4'h9):(4'h9)];
                      reg249 = (^~($unsigned($unsigned(forvar222)) < reg230));
                      reg250 <= (!reg239);
                      reg251 = $signed((!$unsigned($signed(reg241))));
                    end
                  else
                    begin
                      reg249 = forvar221;
                      reg250 <= ($signed($unsigned((wire216 >> (8'ha8)))) ?
                          $signed(reg249[(4'hb):(1'h0)]) : (($unsigned(wire216) ?
                              $signed(forvar222) : forvar224[(2'h2):(1'h0)]) ^~ $signed(forvar221)));
                      reg251 = ("CQ9raG4So1" ?
                          wire216[(4'ha):(1'h0)] : (8'haf));
                      reg252 <= {($signed(((8'hba) && forvar223)) << (~|$unsigned((8'hb7))))};
                    end
                  for (forvar253 = (1'h0); (forvar253 < (1'h1)); forvar253 = (forvar253 + (1'h1)))
                    begin
                      reg254 <= $unsigned(wire219[(1'h0):(1'h0)]);
                      reg255 = {"d0rZA9bGisf1CHn"};
                      reg256 = reg252[(1'h1):(1'h1)];
                    end
                end
              for (forvar257 = (1'h0); (forvar257 < (1'h0)); forvar257 = (forvar257 + (1'h1)))
                begin
                  for (forvar258 = (1'h0); (forvar258 < (2'h3)); forvar258 = (forvar258 + (1'h1)))
                    begin
                      reg259 <= $unsigned(reg229);
                      reg260 <= forvar246[(1'h0):(1'h0)];
                      reg261 = (forvar224[(3'h4):(2'h3)] != forvar246[(3'h4):(2'h3)]);
                    end
                  if ({"W1R6rWnhG1lV0"})
                    begin
                      reg262 <= ((~^$signed($signed(forvar223))) ?
                          forvar233[(1'h1):(1'h1)] : reg244);
                      reg263 <= forvar221;
                      reg264 <= forvar233;
                      reg265 <= ((&$unsigned($signed(wire220))) ?
                          ((|$unsigned(forvar242)) <= reg240) : "Y");
                    end
                  else
                    begin
                      reg266 = ((~&{(forvar224 ?
                              forvar242 : reg249)}) * ($signed(reg227[(3'h4):(2'h3)]) ?
                          ($signed(forvar245) == (~&reg240)) : ($signed(reg229) ?
                              $signed(reg237) : reg238)));
                      reg267 <= ((~^reg248) ?
                          ($unsigned(forvar236[(4'h9):(1'h0)]) ?
                              reg259[(3'h4):(1'h1)] : reg243) : reg230[(4'hd):(3'h7)]);
                      reg268 = reg263;
                    end
                  for (forvar269 = (1'h0); (forvar269 < (2'h2)); forvar269 = (forvar269 + (1'h1)))
                    begin
                      reg270 <= reg266;
                      reg271 = wire216[(3'h6):(1'h0)];
                    end
                end
            end
          else
            begin
              if ($signed("n9VvIqqAaQ"))
                begin
                  if ({(-("Hvz" ? reg266[(1'h1):(1'h1)] : $signed(reg265)))})
                    begin
                      reg242 = wire220[(1'h0):(1'h0)];
                      reg243 = {wire220[(1'h0):(1'h0)]};
                      reg244 = ({$unsigned(reg226)} ?
                          "dDIZu4SElq5Cz" : wire220[(1'h1):(1'h0)]);
                      reg245 = ($unsigned($unsigned(reg251[(3'h4):(1'h1)])) ^~ reg243);
                    end
                  else
                    begin
                      reg246 <= {reg259};
                    end
                  reg248 <= ((~&((reg268 ?
                          forvar232 : wire215) - (~&forvar224))) ?
                      {(!{(8'ha7)})} : $signed(reg234[(4'h8):(2'h3)]));
                  reg249 = $unsigned({$signed(reg244)});
                  if ((~(~|$signed(reg263[(1'h1):(1'h0)]))))
                    begin
                      reg251 = (($unsigned({(8'hab)}) ?
                              (((8'h9c) ? (8'hb4) : reg256) ?
                                  {forvar232} : (!reg235)) : $unsigned($signed(forvar236))) ?
                          "2lv7" : reg265[(4'h8):(4'h8)]);
                      reg253 = reg227[(4'h9):(3'h5)];
                    end
                  else
                    begin
                      reg250 <= "";
                      reg251 = "C2W";
                      reg252 <= "1M8A2LwYSePF";
                      reg253 = forvar269;
                    end
                end
              else
                begin
                  if ($signed($unsigned(reg235)))
                    begin
                      reg242 = (+(((reg242 ?
                              (8'haa) : reg251) >>> $unsigned(reg263)) ?
                          reg234 : ("YSnJ5" & $unsigned(wire220))));
                      reg246 <= ($signed((^~(reg270 ? reg256 : wire215))) ?
                          $signed($signed("")) : $signed((forvar269[(3'h7):(3'h6)] ~^ (reg234 ?
                              forvar222 : reg225))));
                      reg247 = $unsigned((~^((reg231 || (8'hb2)) - (reg270 * reg265))));
                      reg249 = reg247[(4'hd):(4'hd)];
                    end
                  else
                    begin
                      reg242 = {(8'h9c)};
                      reg243 = (!(reg245 ? {(8'hb4)} : (-{reg260})));
                      reg244 = ((-forvar269) & $signed(("NX14V3Gn5XTI" ?
                          (reg254 >>> forvar242) : wire220)));
                      reg246 <= $signed(reg229[(4'h9):(4'h8)]);
                    end
                  for (forvar250 = (1'h0); (forvar250 < (1'h0)); forvar250 = (forvar250 + (1'h1)))
                    begin
                      reg251 = {$unsigned("bQFOZv")};
                      reg253 = reg234[(1'h1):(1'h1)];
                      reg255 = reg246[(2'h3):(1'h0)];
                      reg257 <= $unsigned(reg245);
                    end
                  for (forvar258 = (1'h0); (forvar258 < (1'h1)); forvar258 = (forvar258 + (1'h1)))
                    begin
                      reg261 = reg235[(3'h5):(2'h2)];
                      reg266 = $unsigned($unsigned(($unsigned((8'haa)) ?
                          $unsigned(forvar257) : (+reg255))));
                      reg267 <= (8'h9c);
                    end
                end
              if (wire217)
                begin
                  for (forvar268 = (1'h0); (forvar268 < (1'h0)); forvar268 = (forvar268 + (1'h1)))
                    begin
                      reg269 = $signed(reg267[(2'h2):(1'h1)]);
                      reg270 <= reg253;
                      reg271 = $signed($signed((reg249[(4'h9):(4'h8)] ?
                          ((8'hb3) ^ reg259) : $unsigned((8'ha7)))));
                    end
                end
              else
                begin
                  for (forvar268 = (1'h0); (forvar268 < (2'h3)); forvar268 = (forvar268 + (1'h1)))
                    begin
                      reg269 = reg255[(1'h1):(1'h1)];
                      reg271 = "LMAmfuOaD";
                      reg272 <= (({(~|forvar224)} ?
                          (!(~&wire215)) : $unsigned((reg235 ?
                              reg263 : reg268))) ^~ $signed(((reg231 | forvar221) ?
                          (~reg246) : reg264[(2'h2):(1'h1)])));
                      reg273 = reg264;
                    end
                end
            end
        end
    end
  assign wire274 = wire219[(2'h3):(1'h1)];
  module275 #() modinst1978 (wire1977, clk, reg252, reg267, wire274, reg263);
  always
    @(posedge clk) begin
      reg1979 = reg250[(4'h8):(2'h2)];
      reg1980 = {reg270};
      if ((^~$unsigned({reg262})))
        begin
          for (forvar1981 = (1'h0); (forvar1981 < (2'h3)); forvar1981 = (forvar1981 + (1'h1)))
            begin
              for (forvar1982 = (1'h0); (forvar1982 < (2'h2)); forvar1982 = (forvar1982 + (1'h1)))
                begin
                  if (($unsigned(reg254[(2'h3):(1'h0)]) ?
                      {reg252[(5'h10):(3'h7)]} : $unsigned((~|(reg254 ?
                          reg262 : reg257)))))
                    begin
                      reg1983 = $unsigned((reg248 == ($signed(reg265) ?
                          reg231 : (|reg1980))));
                      reg1984 = reg250[(4'ha):(3'h7)];
                      reg1985 = (8'h9c);
                    end
                  else
                    begin
                      reg1983 = $unsigned("PZMt84Okir");
                      reg1984 = {{$unsigned(wire1977[(3'h5):(3'h4)])}};
                      reg1985 = (((wire216[(3'h6):(2'h3)] ?
                              (reg262 | reg235) : "msJ6oh") - (((8'ha6) ?
                              reg227 : wire216) << $signed(reg252))) ?
                          reg265 : (((wire217 >= reg262) ?
                              (reg252 > wire216) : "DE7IBrKUNCM") ^~ {reg263}));
                      reg1986 <= (~^($unsigned(forvar1981[(1'h0):(1'h0)]) * $signed(((8'ha5) ?
                          reg272 : reg264))));
                    end
                  for (forvar1987 = (1'h0); (forvar1987 < (1'h0)); forvar1987 = (forvar1987 + (1'h1)))
                    begin
                      reg1988 = $unsigned(reg1984);
                    end
                  for (forvar1989 = (1'h0); (forvar1989 < (1'h1)); forvar1989 = (forvar1989 + (1'h1)))
                    begin
                      reg1990 = (reg267 ?
                          (("UQ4Mnco49IN" << (reg227 ?
                              (8'h9c) : reg1988)) << forvar1982) : (~|$unsigned(forvar1987[(1'h0):(1'h0)])));
                      reg1991 = ((wire1977[(4'h8):(3'h4)] & (reg254[(4'h9):(4'h8)] ?
                          reg272 : {(8'hac)})) << {(8'hb7)});
                      reg1992 = reg1988;
                    end
                  for (forvar1993 = (1'h0); (forvar1993 < (2'h2)); forvar1993 = (forvar1993 + (1'h1)))
                    begin
                      reg1994 = ((reg1991 ?
                          $signed($unsigned(reg1984)) : (&(8'ha6))) >> "ON");
                      reg1995 <= $unsigned($unsigned({$signed(wire274)}));
                      reg1996 <= ("pELoW9BXF072c0G" ?
                          $unsigned($unsigned((!reg264))) : "M");
                    end
                end
              reg1997 = reg230;
              for (forvar1998 = (1'h0); (forvar1998 < (2'h3)); forvar1998 = (forvar1998 + (1'h1)))
                begin
                  for (forvar1999 = (1'h0); (forvar1999 < (1'h0)); forvar1999 = (forvar1999 + (1'h1)))
                    begin
                      reg2000 <= ((~$unsigned({(8'ha5)})) ?
                          (((^forvar1987) ?
                                  ((8'hb3) ?
                                      reg250 : reg1994) : $unsigned(reg1984)) ?
                              wire1977[(3'h7):(2'h2)] : (reg225 ?
                                  reg272 : (~^reg229))) : (&(^reg1986)));
                      reg2001 = (~$signed(reg229));
                      reg2002 <= reg250;
                      reg2003 <= (reg1979[(4'ha):(4'ha)] ?
                          (((reg2000 ?
                              forvar1981 : (8'ha7)) >>> (^~reg1986)) <<< $unsigned(reg231[(4'h8):(4'h8)])) : (("Ms8aHxZtB03Ia5" || $unsigned(reg1986)) ?
                              (+reg225[(1'h1):(1'h0)]) : ({(8'hb3)} > reg1988[(4'he):(4'he)])));
                    end
                  reg2004 <= $signed($unsigned((^~(~&reg246))));
                end
              if (reg1992[(3'h5):(1'h1)])
                begin
                  if (reg270[(3'h5):(1'h0)])
                    begin
                      reg2005 = (^~(&(wire218[(4'h8):(1'h0)] ?
                          $unsigned(wire274) : (reg2002 > reg259))));
                    end
                  else
                    begin
                      reg2006 <= reg2002[(3'h6):(1'h0)];
                      reg2007 = reg231;
                      reg2008 = $signed({$signed($unsigned(reg2006))});
                    end
                  reg2009 = (reg250 ?
                      (((wire215 != reg1979) != reg2008[(4'hb):(4'ha)]) ?
                          $signed($signed(reg2007)) : (|reg1992[(2'h3):(2'h3)])) : ({(reg1979 == reg246)} ?
                          ($unsigned(reg259) ?
                              {reg1990} : reg272[(1'h0):(1'h0)]) : "NaRY6izQOOxtz"));
                  if (("" - reg2009))
                    begin
                      reg2010 = {(~reg1992)};
                      reg2011 = reg260;
                    end
                  else
                    begin
                      reg2012 <= ($signed($signed(((8'hba) < (8'ha2)))) >>> reg263);
                      reg2013 = $unsigned($signed((((8'ha2) ?
                              forvar1989 : reg248) ?
                          $unsigned(reg1980) : (wire274 + reg1990))));
                      reg2014 = (reg1983 ?
                          ((^~(forvar1989 < (8'ha9))) >>> $unsigned("")) : reg1992);
                      reg2015 = (^reg1980);
                    end
                  reg2016 <= "w";
                end
              else
                begin
                  reg2006 <= $signed((((forvar1993 == forvar1998) ~^ (reg252 ?
                      reg2003 : wire215)) <= $unsigned((forvar1993 == reg1979))));
                end
            end
        end
      else
        begin
          reg1981 = reg248;
          reg1982 = $signed($unsigned($unsigned(reg2010[(2'h3):(2'h2)])));
        end
      reg2017 = $signed(reg1991[(1'h1):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg2018 = (~|(8'haa));
      reg2019 = "1XGdwWHMlJwoTBX";
    end
  assign wire2020 = (wire1977 ? (8'h9d) : reg248);
  assign wire2021 = reg235[(2'h2):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module275
#(parameter param1976 = ((({(8'ha1)} | ((8'hb9) ? (8'had) : (8'haa))) ? (((8'ha7) ? (8'hb3) : (8'h9c)) >>> (!(8'hb1))) : ((-(8'h9f)) + ((8'h9c) ? (8'hae) : (8'ha2)))) <= ((((8'h9c) ? (8'h9d) : (8'ha2)) != {(8'hb4)}) ? {((8'h9f) == (8'hb2))} : ((!(8'h9e)) < (-(8'hab))))))
(y, clk, wire279, wire278, wire277, wire276);
  output wire [(32'h7a8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire279;
  input wire [(4'hc):(1'h0)] wire278;
  input wire signed [(3'h5):(1'h0)] wire277;
  input wire signed [(4'hd):(1'h0)] wire276;
  wire [(4'he):(1'h0)] wire1975;
  wire signed [(4'hf):(1'h0)] wire1974;
  wire signed [(3'h4):(1'h0)] wire1973;
  wire signed [(4'ha):(1'h0)] wire1972;
  wire [(4'h9):(1'h0)] wire1971;
  wire signed [(2'h3):(1'h0)] wire1232;
  wire [(4'hf):(1'h0)] wire323;
  wire signed [(4'he):(1'h0)] wire1234;
  wire signed [(4'he):(1'h0)] wire1874;
  wire [(4'hf):(1'h0)] wire1876;
  wire [(3'h6):(1'h0)] wire1877;
  wire signed [(3'h6):(1'h0)] wire1878;
  wire signed [(5'h10):(1'h0)] wire1968;
  wire [(4'hb):(1'h0)] wire1969;
  reg [(4'h9):(1'h0)] reg1966 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1963 = (1'h0);
  reg [(5'h10):(1'h0)] reg1960 = (1'h0);
  reg [(4'hf):(1'h0)] reg1951 = (1'h0);
  reg [(2'h3):(1'h0)] reg1949 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1938 = (1'h0);
  reg [(2'h2):(1'h0)] reg1953 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1952 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1948 = (1'h0);
  reg [(3'h7):(1'h0)] reg1945 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1942 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1941 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1940 = (1'h0);
  reg [(4'h9):(1'h0)] reg1939 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1935 = (1'h0);
  reg [(4'ha):(1'h0)] reg1932 = (1'h0);
  reg [(3'h6):(1'h0)] reg1927 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1926 = (1'h0);
  reg [(2'h3):(1'h0)] reg1915 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1913 = (1'h0);
  reg [(2'h3):(1'h0)] reg1910 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1907 = (1'h0);
  reg [(4'hb):(1'h0)] reg1905 = (1'h0);
  reg [(2'h2):(1'h0)] reg1898 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1892 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1890 = (1'h0);
  reg [(4'h9):(1'h0)] reg1889 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1888 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1880 = (1'h0);
  reg [(4'ha):(1'h0)] reg357 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg354 = (1'h0);
  reg [(4'hc):(1'h0)] reg350 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg349 = (1'h0);
  reg [(3'h5):(1'h0)] reg347 = (1'h0);
  reg [(4'ha):(1'h0)] reg345 = (1'h0);
  reg [(4'h8):(1'h0)] reg335 = (1'h0);
  reg [(3'h6):(1'h0)] reg339 = (1'h0);
  reg [(4'hf):(1'h0)] reg336 = (1'h0);
  reg signed [(4'he):(1'h0)] reg331 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg322 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg320 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg319 = (1'h0);
  reg [(5'h10):(1'h0)] reg318 = (1'h0);
  reg [(2'h2):(1'h0)] reg313 = (1'h0);
  reg [(3'h7):(1'h0)] reg311 = (1'h0);
  reg [(4'he):(1'h0)] reg309 = (1'h0);
  reg [(4'hd):(1'h0)] reg308 = (1'h0);
  reg [(5'h10):(1'h0)] reg307 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg302 = (1'h0);
  reg [(4'he):(1'h0)] reg303 = (1'h0);
  reg [(3'h7):(1'h0)] reg300 = (1'h0);
  reg [(4'hd):(1'h0)] reg297 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg293 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg290 = (1'h0);
  reg [(4'h8):(1'h0)] reg289 = (1'h0);
  reg [(2'h3):(1'h0)] reg286 = (1'h0);
  reg [(4'h8):(1'h0)] reg284 = (1'h0);
  reg [(4'hc):(1'h0)] reg280 = (1'h0);
  reg [(4'hd):(1'h0)] reg1967 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1965 = (1'h0);
  reg [(3'h7):(1'h0)] reg1964 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1962 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1961 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1959 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1958 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1957 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1956 = (1'h0);
  reg [(4'hb):(1'h0)] reg1955 = (1'h0);
  reg [(4'hc):(1'h0)] reg1954 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1935 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1934 = (1'h0);
  reg [(4'hd):(1'h0)] reg1933 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1951 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1950 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1949 = (1'h0);
  reg [(4'he):(1'h0)] reg1947 = (1'h0);
  reg [(4'hd):(1'h0)] reg1946 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1944 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1943 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1938 = (1'h0);
  reg [(4'hf):(1'h0)] reg1937 = (1'h0);
  reg [(4'hf):(1'h0)] reg1936 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1934 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1933 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1931 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1930 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1929 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1928 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1925 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1924 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1923 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1922 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1921 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1920 = (1'h0);
  reg [(5'h10):(1'h0)] reg1919 = (1'h0);
  reg [(4'he):(1'h0)] reg1918 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1917 = (1'h0);
  reg [(4'h8):(1'h0)] reg1916 = (1'h0);
  reg [(3'h6):(1'h0)] reg1914 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1912 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1911 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1909 = (1'h0);
  reg [(4'h9):(1'h0)] reg1908 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1906 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1904 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1903 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1902 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1901 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1900 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1895 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1900 = (1'h0);
  reg [(4'hf):(1'h0)] reg1899 = (1'h0);
  reg [(5'h10):(1'h0)] reg1897 = (1'h0);
  reg [(4'he):(1'h0)] reg1896 = (1'h0);
  reg [(3'h6):(1'h0)] reg1895 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1894 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1893 = (1'h0);
  reg [(3'h4):(1'h0)] reg1891 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1887 = (1'h0);
  reg [(4'hd):(1'h0)] reg1886 = (1'h0);
  reg [(4'hf):(1'h0)] reg1885 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1884 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1883 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1882 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1881 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1879 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg356 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg355 = (1'h0);
  reg signed [(4'he):(1'h0)] reg353 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar352 = (1'h0);
  reg [(4'h8):(1'h0)] reg351 = (1'h0);
  reg [(3'h4):(1'h0)] reg348 = (1'h0);
  reg [(3'h5):(1'h0)] forvar346 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg344 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg343 = (1'h0);
  reg [(5'h10):(1'h0)] forvar342 = (1'h0);
  reg [(4'hd):(1'h0)] forvar341 = (1'h0);
  reg [(5'h10):(1'h0)] reg340 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar338 = (1'h0);
  reg [(4'h8):(1'h0)] reg338 = (1'h0);
  reg [(4'h8):(1'h0)] reg337 = (1'h0);
  reg [(4'ha):(1'h0)] forvar335 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg334 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg333 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg332 = (1'h0);
  reg [(4'hd):(1'h0)] reg330 = (1'h0);
  reg [(4'h9):(1'h0)] reg329 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg328 = (1'h0);
  reg [(4'h9):(1'h0)] reg327 = (1'h0);
  reg [(4'hb):(1'h0)] reg326 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg325 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar324 = (1'h0);
  reg [(2'h3):(1'h0)] reg324 = (1'h0);
  reg [(4'he):(1'h0)] forvar321 = (1'h0);
  reg [(4'hd):(1'h0)] reg317 = (1'h0);
  reg [(4'h9):(1'h0)] forvar316 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg315 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg314 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg312 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg310 = (1'h0);
  reg [(3'h4):(1'h0)] forvar307 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar296 = (1'h0);
  reg [(4'hb):(1'h0)] reg294 = (1'h0);
  reg [(4'hd):(1'h0)] forvar290 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar288 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar285 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar283 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar282 = (1'h0);
  reg [(4'h9):(1'h0)] reg281 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar303 = (1'h0);
  reg [(4'ha):(1'h0)] forvar299 = (1'h0);
  reg [(4'hd):(1'h0)] reg306 = (1'h0);
  reg [(4'ha):(1'h0)] reg305 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg304 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar302 = (1'h0);
  reg [(4'h9):(1'h0)] reg301 = (1'h0);
  reg signed [(4'he):(1'h0)] reg299 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar298 = (1'h0);
  reg [(3'h7):(1'h0)] reg298 = (1'h0);
  reg [(4'he):(1'h0)] reg296 = (1'h0);
  reg [(2'h2):(1'h0)] reg295 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar294 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg292 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg291 = (1'h0);
  reg [(2'h3):(1'h0)] reg288 = (1'h0);
  reg [(3'h4):(1'h0)] reg287 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg285 = (1'h0);
  reg [(4'ha):(1'h0)] reg283 = (1'h0);
  reg [(4'hd):(1'h0)] reg282 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar281 = (1'h0);
  reg [(4'h9):(1'h0)] forvar280 = (1'h0);
  assign y = {wire1974,
                 wire1232,
                 wire323,
                 wire1878,
                 wire1968,
                 reg1966,
                 reg1941,
                 reg1939,
                 reg1926,
                 reg1905,
                 reg354,
                 reg347,
                 reg336,
                 reg322,
                 reg320,
                 reg319,
                 reg313,
                 reg309,
                 reg308,
                 reg300,
                 reg290,
                 reg289,
                 reg286,
                 reg280,
                 reg1964,
                 forvar1962,
                 reg1959,
                 forvar1958,
                 reg1956,
                 forvar1935,
                 reg1933,
                 forvar1949,
                 reg1947,
                 reg1946,
                 forvar1944,
                 reg1936,
                 reg1934,
                 forvar1933,
                 reg1931,
                 reg1919,
                 reg1918,
                 reg1916,
                 forvar1912,
                 forvar1911,
                 reg1908,
                 reg1906,
                 reg1901,
                 forvar1895,
                 reg1894,
                 reg1886,
                 reg1884,
                 reg356,
                 reg355,
                 reg353,
                 forvar352,
                 forvar338,
                 reg337,
                 forvar324,
                 reg324,
                 reg317,
                 forvar316,
                 reg315,
                 reg314,
                 forvar296,
                 reg294,
                 forvar282,
                 reg281,
                 reg306,
                 reg304,
                 reg299,
                 forvar298,
                 reg298,
                 reg296,
                 reg288,
                 reg285,
                 reg282,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (("H" ? (8'h9d) : wire279))
        begin
          if (({$signed((|wire276))} <<< wire276))
            begin
              reg280 <= $unsigned(wire279);
            end
          else
            begin
              for (forvar280 = (1'h0); (forvar280 < (1'h0)); forvar280 = (forvar280 + (1'h1)))
                begin
                  for (forvar281 = (1'h0); (forvar281 < (2'h3)); forvar281 = (forvar281 + (1'h1)))
                    begin
                      reg282 = ((8'hba) ?
                          ({""} ? $signed({wire276}) : forvar281) : "zIQAI");
                      reg283 = ($signed("9bdn1bBW") ?
                          (8'hb3) : ("2swriMQA3EOb0uB" >>> (~^(^~(8'hb3)))));
                      reg284 <= {(~^forvar281)};
                      reg285 = {(^$unsigned(reg284))};
                    end
                  if ((^~(&(!(forvar280 ? wire279 : wire278)))))
                    begin
                      reg286 <= $signed($unsigned(reg280));
                      reg287 = $unsigned(reg280[(4'hb):(1'h0)]);
                      reg288 = $signed(($signed(reg285[(2'h3):(1'h1)]) == $signed($unsigned(forvar281))));
                      reg289 <= wire277;
                    end
                  else
                    begin
                      reg286 <= (~&($signed({reg287}) && wire277));
                      reg287 = wire279[(3'h5):(3'h5)];
                      reg289 <= $unsigned((~|reg280[(4'h9):(1'h1)]));
                      reg290 <= $signed($unsigned($signed((~wire277))));
                    end
                  reg291 = $unsigned(($unsigned($signed(forvar281)) ~^ reg289[(3'h6):(1'h1)]));
                end
              reg292 = reg290[(4'h9):(3'h6)];
              reg293 <= ({$signed(reg290[(4'hb):(3'h6)])} << (~|((~&reg284) ^~ (wire277 ?
                  reg290 : reg287))));
              for (forvar294 = (1'h0); (forvar294 < (2'h3)); forvar294 = (forvar294 + (1'h1)))
                begin
                  reg295 = ($unsigned("nl6sdoq") <<< reg282[(3'h5):(1'h0)]);
                  reg296 = "vWber0";
                  reg297 <= "U46";
                end
            end
          if ((+(~|"")))
            begin
              if ($signed((8'hb9)))
                begin
                  reg298 = ($unsigned($signed(reg296)) == {$signed((reg284 ?
                          wire278 : (8'h9e)))});
                end
              else
                begin
                  for (forvar298 = (1'h0); (forvar298 < (1'h1)); forvar298 = (forvar298 + (1'h1)))
                    begin
                      reg299 = (~|($unsigned({reg286}) ^ {$unsigned((8'ha5))}));
                      reg300 <= $signed((8'ha1));
                    end
                  reg301 = ({((reg293 ?
                          (8'hae) : forvar294) && wire277)} & $unsigned(wire277));
                  for (forvar302 = (1'h0); (forvar302 < (2'h3)); forvar302 = (forvar302 + (1'h1)))
                    begin
                      reg303 <= wire276;
                      reg304 = reg295;
                      reg305 = {"YR9Z5GaTKuzoa"};
                      reg306 = {{(^~(reg288 ? reg287 : reg289))}};
                    end
                end
            end
          else
            begin
              if ($signed((reg286 >= reg297)))
                begin
                  reg298 = "NnE0YmqD";
                  for (forvar299 = (1'h0); (forvar299 < (1'h1)); forvar299 = (forvar299 + (1'h1)))
                    begin
                      reg300 <= $unsigned("TbuV4IM7Y8RO");
                      reg302 <= wire276[(1'h0):(1'h0)];
                    end
                  for (forvar303 = (1'h0); (forvar303 < (1'h1)); forvar303 = (forvar303 + (1'h1)))
                    begin
                      reg304 = $signed(reg302);
                      reg305 = $signed(forvar281);
                      reg307 <= reg295;
                      reg308 <= ((8'ha3) <= (((8'h9e) ^~ "hzuxk") < (reg280 && (forvar294 ?
                          reg302 : (8'haf)))));
                    end
                end
              else
                begin
                  reg298 = ((~&"vvD1BfqbkgJq") > (wire277 ?
                      forvar299 : "P9zNyYiudslqsmP"));
                end
            end
        end
      else
        begin
          if ($unsigned($signed($signed((~reg301)))))
            begin
              reg280 <= reg283;
            end
          else
            begin
              reg281 = $signed(reg280[(2'h2):(1'h0)]);
              for (forvar282 = (1'h0); (forvar282 < (2'h2)); forvar282 = (forvar282 + (1'h1)))
                begin
                  for (forvar283 = (1'h0); (forvar283 < (2'h3)); forvar283 = (forvar283 + (1'h1)))
                    begin
                      reg284 <= $unsigned($unsigned(reg281[(1'h0):(1'h0)]));
                    end
                end
            end
          for (forvar285 = (1'h0); (forvar285 < (2'h2)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg287 = $unsigned($signed(reg295[(1'h0):(1'h0)]));
              for (forvar288 = (1'h0); (forvar288 < (1'h0)); forvar288 = (forvar288 + (1'h1)))
                begin
                  reg289 <= $unsigned(({(reg301 ? reg286 : reg286)} ?
                      (^~$signed((8'ha6))) : $signed(reg306)));
                  for (forvar290 = (1'h0); (forvar290 < (1'h1)); forvar290 = (forvar290 + (1'h1)))
                    begin
                      reg291 = ((reg298[(3'h6):(1'h0)] | ((^~reg298) ?
                              ((8'haf) ? reg287 : reg304) : (reg284 ?
                                  forvar290 : forvar290))) ?
                          (~$signed($signed(reg281))) : ($unsigned((forvar285 ?
                                  reg299 : (8'h9c))) ?
                              reg306[(3'h7):(1'h1)] : $signed((forvar302 ?
                                  (8'haf) : forvar294))));
                      reg293 <= $unsigned((^reg301[(3'h5):(2'h2)]));
                      reg294 = (8'ha9);
                      reg295 = {((forvar281 ?
                              (reg285 <<< reg303) : (reg281 ?
                                  forvar282 : reg301)) >> "hPHttXtp4xy")};
                    end
                end
              for (forvar296 = (1'h0); (forvar296 < (2'h2)); forvar296 = (forvar296 + (1'h1)))
                begin
                  reg298 = (reg292[(4'h9):(3'h4)] ?
                      ((~(reg297 ~^ forvar302)) ?
                          ($unsigned(forvar298) - reg292[(4'h9):(4'h8)]) : $signed(forvar294[(2'h3):(1'h0)])) : (((forvar303 >= reg281) ?
                          ((8'hba) ^~ reg282) : (~forvar299)) > $signed(((8'ha0) | (8'hb8)))));
                  reg300 <= (^~(reg281 ?
                      $unsigned(reg302[(1'h0):(1'h0)]) : reg288[(2'h3):(1'h1)]));
                  reg301 = $signed(reg294);
                  for (forvar302 = (1'h0); (forvar302 < (1'h0)); forvar302 = (forvar302 + (1'h1)))
                    begin
                      reg304 = forvar302[(3'h6):(2'h2)];
                      reg305 = $signed(forvar282[(2'h2):(1'h1)]);
                      reg306 = reg302[(2'h3):(2'h2)];
                    end
                end
              for (forvar307 = (1'h0); (forvar307 < (1'h1)); forvar307 = (forvar307 + (1'h1)))
                begin
                  if (forvar290[(3'h6):(1'h1)])
                    begin
                      reg308 <= (|{reg290});
                      reg309 <= reg285[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg310 = $unsigned(((~^$unsigned(reg293)) ?
                          $signed(((8'ha3) ?
                              wire278 : wire278)) : ("f" - reg309[(4'h9):(3'h4)])));
                      reg311 <= ($unsigned(((wire278 ?
                              (8'ha1) : reg306) != "zNvQzi")) ?
                          $unsigned("1IO6kcQ8n") : reg284);
                    end
                  if (((|(reg283 >>> (reg286 && forvar294))) <<< reg290[(3'h4):(2'h3)]))
                    begin
                      reg312 = reg291;
                    end
                  else
                    begin
                      reg312 = (8'ha3);
                      reg313 <= reg299;
                      reg314 = reg313[(2'h2):(2'h2)];
                      reg315 = $unsigned($unsigned(({reg295} ?
                          (forvar298 ?
                              forvar290 : reg308) : $unsigned(forvar281))));
                    end
                  for (forvar316 = (1'h0); (forvar316 < (1'h0)); forvar316 = (forvar316 + (1'h1)))
                    begin
                      reg317 = (reg301[(2'h3):(1'h1)] < $signed(({reg288} ?
                          (reg305 ?
                              reg307 : reg299) : wire276[(3'h6):(3'h6)])));
                      reg318 <= "5hmwtg";
                      reg319 <= "P5kfhghgqT";
                      reg320 <= $signed(((8'hae) ? reg280 : "UfXF2J"));
                    end
                  for (forvar321 = (1'h0); (forvar321 < (2'h2)); forvar321 = (forvar321 + (1'h1)))
                    begin
                      reg322 <= ($signed({$unsigned(forvar298)}) ?
                          (&((forvar282 * reg308) ?
                              (reg286 ?
                                  reg314 : forvar282) : (^~(8'hb7)))) : (|(reg280[(4'hc):(3'h6)] | (forvar307 < wire279))));
                    end
                end
            end
        end
    end
  assign wire323 = reg322;
  always
    @(posedge clk) begin
      if ($unsigned((reg320[(2'h2):(2'h2)] ?
          $signed("TWW9GPL") : $signed({(8'haa)}))))
        begin
          reg324 = (("KOGiyGnuTyw" > ($unsigned((8'h9d)) - {reg302})) >= ($unsigned($unsigned((8'hb4))) ?
              (8'hb5) : $unsigned((^~reg297))));
        end
      else
        begin
          if ((reg318[(3'h7):(2'h3)] ?
              $unsigned($unsigned("ibK")) : $signed(wire323)))
            begin
              if ($unsigned(reg307))
                begin
                  for (forvar324 = (1'h0); (forvar324 < (1'h0)); forvar324 = (forvar324 + (1'h1)))
                    begin
                      reg325 = (&(reg280 << (^~{(8'h9e)})));
                      reg326 = $signed($signed(((~^reg290) ?
                          reg325[(1'h1):(1'h0)] : (~^reg293))));
                      reg327 = $signed(reg307);
                    end
                  if ($signed(($signed((^~wire276)) ?
                      reg318[(3'h5):(1'h1)] : forvar324[(1'h0):(1'h0)])))
                    begin
                      reg328 = reg326[(1'h1):(1'h1)];
                      reg329 = (wire276[(4'ha):(4'ha)] ?
                          $unsigned(((reg320 ? forvar324 : wire277) ?
                              (reg319 ?
                                  reg303 : reg322) : $unsigned(reg328))) : (^$unsigned((reg326 < reg319))));
                      reg330 = "rXVF07";
                    end
                  else
                    begin
                      reg331 <= (reg297[(4'ha):(1'h1)] || reg313);
                      reg332 = (reg324[(2'h2):(1'h0)] ?
                          ("" ?
                              $unsigned($unsigned(reg329)) : $unsigned({reg328})) : (($signed(reg331) << reg330) ?
                              reg328 : reg330));
                      reg333 = $unsigned((!(reg322 ^ "")));
                    end
                end
              else
                begin
                  if ((($signed({reg313}) ?
                      ($signed(reg293) ?
                          (reg332 ?
                              reg327 : reg318) : $signed(reg302)) : wire277[(1'h0):(1'h0)]) <<< "iqVQclz9A"))
                    begin
                      reg324 = reg330;
                      reg325 = $signed(reg280);
                      reg326 = (+$unsigned($unsigned($unsigned(reg320))));
                    end
                  else
                    begin
                      reg324 = ((!"xST3A") ?
                          ({reg311[(3'h7):(2'h3)]} ?
                              reg329[(1'h0):(1'h0)] : ((8'hb3) ?
                                  reg302[(3'h4):(1'h1)] : wire279[(3'h4):(1'h1)])) : $unsigned("ZDe"));
                      reg331 <= reg308[(1'h1):(1'h1)];
                    end
                end
              if (($unsigned((^~(wire323 == reg303))) > reg319[(3'h4):(2'h2)]))
                begin
                  reg334 = {(reg280 << (reg300[(1'h0):(1'h0)] > (8'hb3)))};
                  for (forvar335 = (1'h0); (forvar335 < (2'h3)); forvar335 = (forvar335 + (1'h1)))
                    begin
                      reg336 <= "OZd9YBhoJ";
                    end
                  reg337 = $signed("Qhxupe");
                  reg338 = (+("7P" ?
                      ((!reg322) >= $unsigned((8'hb3))) : $signed($signed(reg313))));
                end
              else
                begin
                  reg334 = reg337;
                end
              reg339 <= (reg327[(1'h1):(1'h0)] ?
                  ("" ?
                      reg290[(3'h7):(3'h7)] : (|reg303[(3'h7):(3'h7)])) : {$unsigned($unsigned(reg302))});
            end
          else
            begin
              for (forvar324 = (1'h0); (forvar324 < (1'h1)); forvar324 = (forvar324 + (1'h1)))
                begin
                  if (reg290)
                    begin
                      reg325 = $unsigned((+(reg311 ?
                          $signed(reg289) : $signed(reg289))));
                    end
                  else
                    begin
                      reg325 = ("M0467" == wire323[(3'h7):(2'h3)]);
                      reg331 <= $signed(forvar324[(3'h4):(1'h1)]);
                      reg332 = reg320;
                      reg333 = {(8'ha0)};
                    end
                  reg335 <= $unsigned($unsigned(((reg289 <= wire276) ?
                      (-reg337) : wire279[(3'h5):(3'h4)])));
                  reg337 = reg303[(1'h1):(1'h0)];
                  for (forvar338 = (1'h0); (forvar338 < (2'h3)); forvar338 = (forvar338 + (1'h1)))
                    begin
                      reg340 = ($signed(reg318) != ({$unsigned(reg332)} - $unsigned((~&reg322))));
                    end
                end
              for (forvar341 = (1'h0); (forvar341 < (2'h2)); forvar341 = (forvar341 + (1'h1)))
                begin
                  for (forvar342 = (1'h0); (forvar342 < (1'h1)); forvar342 = (forvar342 + (1'h1)))
                    begin
                      reg343 = ((~|$unsigned((reg309 ? reg302 : wire276))) ?
                          (reg327 ^ forvar342) : $signed(((reg340 ?
                                  reg293 : forvar342) ?
                              "aKsHcgFvGo5i2Rh" : reg290)));
                      reg344 = $signed($unsigned("RmObC426"));
                      reg345 <= (~&(&{(reg325 ? (8'ha5) : reg308)}));
                    end
                  for (forvar346 = (1'h0); (forvar346 < (1'h0)); forvar346 = (forvar346 + (1'h1)))
                    begin
                      reg347 <= $signed(("78Z" ?
                          ($unsigned((8'ha8)) - $unsigned(reg340)) : (8'ha4)));
                      reg348 = {((!(reg337 ? forvar335 : (8'ha7))) ?
                              reg313 : $signed(forvar324))};
                      reg349 <= reg280;
                      reg350 <= ({(~&(forvar346 << reg329))} <= ($signed((reg348 == reg328)) <<< ((reg297 >> reg331) ?
                          reg286[(1'h1):(1'h0)] : reg334)));
                    end
                  reg351 = "Hq9n";
                  for (forvar352 = (1'h0); (forvar352 < (1'h0)); forvar352 = (forvar352 + (1'h1)))
                    begin
                      reg353 = forvar341;
                      reg354 <= {$signed((((8'hb4) ? forvar352 : reg340) ?
                              (reg340 & reg353) : (reg328 || forvar338)))};
                      reg355 = $signed(((reg353 <<< $signed(reg340)) != {{reg319}}));
                      reg356 = (((~^(reg348 <<< reg313)) ?
                              "WgW" : ({reg327} ~^ (-reg336))) ?
                          (((reg336 ? forvar341 : reg319) ?
                              (~wire277) : reg338[(2'h2):(1'h1)]) - forvar346) : $unsigned($unsigned("P")));
                    end
                end
            end
        end
      reg357 <= $unsigned(("4GxQ1u4E1cFg" ^ (!((8'hb6) * forvar341))));
    end
  module358 #() modinst1233 (wire1232, clk, reg303, reg336, reg320, reg302, wire279);
  assign wire1234 = ((reg319 ?
                        (+(wire278 - reg357)) : (wire278 >> reg302[(4'he):(3'h7)])) + ("cUcJ8" > (wire278 << (reg345 >> reg280))));
  module1235 #() modinst1875 (.wire1238(reg308), .clk(clk), .wire1237(reg350), .wire1239(reg319), .y(wire1874), .wire1236(reg300));
  assign wire1876 = (reg335 | ((((8'hb3) ?
                        (8'haa) : wire1234) || reg345[(3'h5):(1'h0)]) == (8'hb8)));
  assign wire1877 = reg302;
  assign wire1878 = "oPCoRVc";
  always
    @(posedge clk) begin
      reg1879 = (reg302[(3'h4):(1'h1)] + wire278[(3'h5):(2'h3)]);
      reg1880 <= (|($unsigned((reg313 << reg349)) >> ($signed((8'ha9)) ~^ {reg320})));
      for (forvar1881 = (1'h0); (forvar1881 < (1'h0)); forvar1881 = (forvar1881 + (1'h1)))
        begin
          for (forvar1882 = (1'h0); (forvar1882 < (2'h2)); forvar1882 = (forvar1882 + (1'h1)))
            begin
              for (forvar1883 = (1'h0); (forvar1883 < (2'h3)); forvar1883 = (forvar1883 + (1'h1)))
                begin
                  if (wire277)
                    begin
                      reg1884 = (($unsigned($signed(forvar1881)) || ($unsigned(wire323) >>> reg286[(2'h3):(1'h1)])) <= (+($signed(wire276) <= {wire323})));
                      reg1885 = reg331;
                    end
                  else
                    begin
                      reg1884 = (~&(^~(reg318 | reg345[(3'h7):(1'h0)])));
                      reg1885 = {{(wire1234 && (8'h9d))}};
                      reg1886 = reg357[(3'h7):(3'h5)];
                    end
                  for (forvar1887 = (1'h0); (forvar1887 < (2'h3)); forvar1887 = (forvar1887 + (1'h1)))
                    begin
                      reg1888 <= (~|$unsigned(reg303[(4'ha):(4'ha)]));
                      reg1889 <= (reg1879[(1'h0):(1'h0)] >>> $unsigned($unsigned($unsigned(wire278))));
                      reg1890 <= $unsigned((~^$signed($unsigned(wire1877))));
                      reg1891 = (^reg307);
                    end
                  reg1892 <= "CdSAgdXarYR";
                  for (forvar1893 = (1'h0); (forvar1893 < (1'h1)); forvar1893 = (forvar1893 + (1'h1)))
                    begin
                      reg1894 = wire1877[(1'h0):(1'h0)];
                    end
                end
              if (reg335)
                begin
                  reg1895 = {{(~$signed(reg336))}};
                  if ((((forvar1887 ? ((8'hac) - reg350) : reg1894) ^~ reg307) ?
                      $signed($unsigned({reg1890})) : (((reg1884 ^ reg1885) | (reg286 * forvar1893)) <<< (8'had))))
                    begin
                      reg1896 = reg284;
                      reg1897 = ("3q5vBegNCEOJ1" ?
                          $signed($unsigned($unsigned(reg313))) : (~^reg1888[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1898 <= (&$signed((~(reg335 || reg318))));
                      reg1899 = wire276[(2'h3):(2'h3)];
                    end
                  reg1900 = {forvar1882[(1'h0):(1'h0)]};
                end
              else
                begin
                  for (forvar1895 = (1'h0); (forvar1895 < (2'h3)); forvar1895 = (forvar1895 + (1'h1)))
                    begin
                      reg1898 <= $unsigned((($unsigned(wire1878) ?
                              $signed(wire1878) : (wire323 < forvar1887)) ?
                          wire277 : $unsigned({(8'ha9)})));
                      reg1899 = "478Bqe69zV";
                    end
                  for (forvar1900 = (1'h0); (forvar1900 < (1'h1)); forvar1900 = (forvar1900 + (1'h1)))
                    begin
                      reg1901 = $signed($unsigned($signed((8'hac))));
                      reg1902 = {reg302[(4'hf):(1'h1)]};
                      reg1903 = forvar1900[(2'h2):(1'h0)];
                    end
                  for (forvar1904 = (1'h0); (forvar1904 < (1'h0)); forvar1904 = (forvar1904 + (1'h1)))
                    begin
                      reg1905 <= ((~^(+$signed(reg354))) == (($signed(reg1894) >>> $unsigned(wire1876)) ^ wire1877));
                      reg1906 = {$unsigned((^$unsigned(reg1894)))};
                      reg1907 <= $unsigned({reg345[(4'h9):(1'h1)]});
                      reg1908 = $unsigned((reg1896[(2'h3):(2'h3)] ?
                          $signed((reg309 ? (8'hb0) : reg309)) : reg331));
                    end
                end
            end
          for (forvar1909 = (1'h0); (forvar1909 < (2'h2)); forvar1909 = (forvar1909 + (1'h1)))
            begin
              reg1910 <= (^~(reg313[(2'h2):(2'h2)] ?
                  "w" : reg300[(2'h3):(1'h0)]));
            end
          for (forvar1911 = (1'h0); (forvar1911 < (1'h0)); forvar1911 = (forvar1911 + (1'h1)))
            begin
              for (forvar1912 = (1'h0); (forvar1912 < (1'h0)); forvar1912 = (forvar1912 + (1'h1)))
                begin
                  if (forvar1883)
                    begin
                      reg1913 <= $unsigned((&$unsigned($signed(forvar1881))));
                      reg1914 = (("I0XvfUfxg7" ?
                          wire1232[(1'h0):(1'h0)] : ((forvar1904 ^ reg286) ?
                              (reg1913 >> reg1908) : (^reg1906))) | wire1874[(4'h9):(3'h4)]);
                      reg1915 <= (8'hab);
                      reg1916 = ($unsigned("aigToRGPCmbyft3") <<< (forvar1881[(2'h2):(2'h2)] >> $signed(((8'ha6) >= forvar1904))));
                    end
                  else
                    begin
                      reg1913 <= reg1890[(3'h6):(3'h5)];
                      reg1914 = $unsigned(((reg297 ?
                          wire277 : (+(8'hb7))) ^~ forvar1887[(4'hb):(1'h1)]));
                      reg1916 = $unsigned($unsigned((((8'ha7) - forvar1904) ?
                          forvar1900[(1'h0):(1'h0)] : (^~reg297))));
                    end
                  for (forvar1917 = (1'h0); (forvar1917 < (2'h2)); forvar1917 = (forvar1917 + (1'h1)))
                    begin
                      reg1918 = $unsigned(wire323[(3'h4):(1'h0)]);
                      reg1919 = ((|$signed(reg1889)) ? reg1913 : "Sg");
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1920 = (1'h0); (forvar1920 < (1'h1)); forvar1920 = (forvar1920 + (1'h1)))
        begin
          for (forvar1921 = (1'h0); (forvar1921 < (2'h3)); forvar1921 = (forvar1921 + (1'h1)))
            begin
              for (forvar1922 = (1'h0); (forvar1922 < (1'h1)); forvar1922 = (forvar1922 + (1'h1)))
                begin
                  for (forvar1923 = (1'h0); (forvar1923 < (1'h1)); forvar1923 = (forvar1923 + (1'h1)))
                    begin
                      reg1924 = (reg290[(4'hd):(4'ha)] ?
                          {(~|reg320[(3'h7):(3'h4)])} : reg297[(3'h7):(3'h7)]);
                      reg1925 = $unsigned(($unsigned(wire1878) ^ {reg284}));
                      reg1926 <= (~|$signed(reg336[(3'h6):(1'h0)]));
                      reg1927 <= "NrHM9KXnql";
                    end
                  for (forvar1928 = (1'h0); (forvar1928 < (2'h2)); forvar1928 = (forvar1928 + (1'h1)))
                    begin
                      reg1929 = {forvar1922[(2'h3):(1'h0)]};
                      reg1930 = (wire276 ?
                          $signed($unsigned(wire276[(3'h7):(2'h3)])) : reg1929[(3'h6):(1'h0)]);
                      reg1931 = reg280;
                    end
                  reg1932 <= reg1930[(3'h4):(2'h3)];
                end
            end
          if ({$unsigned($unsigned($signed(reg286)))})
            begin
              if ($signed((+((&(8'ha8)) ?
                  reg354[(4'h9):(3'h6)] : (reg1924 & reg303)))))
                begin
                  for (forvar1933 = (1'h0); (forvar1933 < (1'h1)); forvar1933 = (forvar1933 + (1'h1)))
                    begin
                      reg1934 = (wire1877[(3'h5):(3'h4)] >= (~reg313[(1'h0):(1'h0)]));
                      reg1935 <= (^~$unsigned(wire1877));
                      reg1936 = (!reg1898[(1'h1):(1'h1)]);
                      reg1937 = reg307;
                    end
                end
              else
                begin
                  for (forvar1933 = (1'h0); (forvar1933 < (1'h1)); forvar1933 = (forvar1933 + (1'h1)))
                    begin
                      reg1934 = reg302;
                      reg1936 = reg290[(4'hb):(3'h5)];
                    end
                end
              for (forvar1938 = (1'h0); (forvar1938 < (2'h2)); forvar1938 = (forvar1938 + (1'h1)))
                begin
                  reg1939 <= (~^(|((~wire278) == (&wire279))));
                  if (forvar1921[(4'he):(1'h1)])
                    begin
                      reg1940 <= $signed((reg339 ?
                          $unsigned($signed(reg1939)) : reg350[(2'h3):(2'h2)]));
                      reg1941 <= $signed(reg318[(5'h10):(4'h9)]);
                      reg1942 <= {$signed(((reg311 << reg300) ?
                              reg1935 : $unsigned(wire278)))};
                    end
                  else
                    begin
                      reg1940 <= "S1CdDoulStPCfnX";
                      reg1941 <= ($signed(reg347) >= reg335);
                      reg1942 <= $signed((&(!"A")));
                    end
                  reg1943 = $unsigned((!forvar1920));
                end
              if ($signed(wire276[(2'h2):(1'h0)]))
                begin
                  for (forvar1944 = (1'h0); (forvar1944 < (1'h1)); forvar1944 = (forvar1944 + (1'h1)))
                    begin
                      reg1945 <= ($unsigned($signed({reg1889})) == ((8'hab) < reg300[(3'h4):(2'h3)]));
                      reg1946 = reg336;
                      reg1947 = ({(reg1932 ? $unsigned(reg1890) : (^~reg336))} ?
                          "38QZGue63XAX" : (^"WQpQProbEF"));
                      reg1948 <= (|$unsigned($signed(reg290[(2'h3):(2'h2)])));
                    end
                  for (forvar1949 = (1'h0); (forvar1949 < (2'h2)); forvar1949 = (forvar1949 + (1'h1)))
                    begin
                      reg1950 = $signed((~&(|(reg322 ? reg1939 : wire277))));
                    end
                  for (forvar1951 = (1'h0); (forvar1951 < (1'h1)); forvar1951 = (forvar1951 + (1'h1)))
                    begin
                      reg1952 <= $signed($unsigned($unsigned((reg347 ?
                          reg1932 : (8'ha6)))));
                      reg1953 <= $unsigned(reg357[(3'h7):(2'h3)]);
                    end
                end
              else
                begin
                  for (forvar1944 = (1'h0); (forvar1944 < (2'h2)); forvar1944 = (forvar1944 + (1'h1)))
                    begin
                      reg1946 = {(forvar1933 <= {$unsigned(reg331)})};
                    end
                end
            end
          else
            begin
              reg1933 = $signed((reg1936 ?
                  (((8'ha0) & reg1926) <= $signed(reg1889)) : wire1877));
              for (forvar1934 = (1'h0); (forvar1934 < (1'h1)); forvar1934 = (forvar1934 + (1'h1)))
                begin
                  for (forvar1935 = (1'h0); (forvar1935 < (1'h0)); forvar1935 = (forvar1935 + (1'h1)))
                    begin
                      reg1938 <= {($signed($signed((8'haf))) | {(+wire323)})};
                    end
                  reg1943 = (forvar1920 < $unsigned({wire276}));
                  for (forvar1944 = (1'h0); (forvar1944 < (2'h3)); forvar1944 = (forvar1944 + (1'h1)))
                    begin
                      reg1946 = ((~&reg309[(4'hb):(4'h9)]) >= $signed(reg1889));
                      reg1947 = (~^(-(8'h9c)));
                    end
                  if (($unsigned((^"gh5Op7pVZSGRGp1")) ?
                      reg1927 : ($unsigned(reg1948) ^~ ((forvar1921 ?
                          reg1953 : wire277) << reg1942))))
                    begin
                      reg1948 <= reg1939[(3'h7):(3'h4)];
                      reg1949 <= {forvar1935};
                      reg1950 = ((~|(((8'h9c) ? reg322 : wire276) ?
                              reg1933[(4'h9):(1'h0)] : (forvar1951 || reg1943))) ?
                          "g" : $signed(reg1905));
                      reg1951 <= wire1234;
                    end
                  else
                    begin
                      reg1950 = $signed($unsigned((^~(^~(8'ha2)))));
                      reg1951 <= $signed((reg1934[(3'h6):(2'h3)] || reg1947));
                      reg1954 = $signed((^~$signed({reg1929})));
                      reg1955 = (8'hba);
                    end
                end
              reg1956 = $signed(reg302);
              for (forvar1957 = (1'h0); (forvar1957 < (1'h1)); forvar1957 = (forvar1957 + (1'h1)))
                begin
                  for (forvar1958 = (1'h0); (forvar1958 < (2'h3)); forvar1958 = (forvar1958 + (1'h1)))
                    begin
                      reg1959 = "u5J0";
                      reg1960 <= reg1907[(4'he):(3'h4)];
                      reg1961 = {($unsigned(forvar1949) ?
                              ("ft" >>> forvar1922[(1'h0):(1'h0)]) : (&"fWdyGyHX8JT7T"))};
                    end
                  for (forvar1962 = (1'h0); (forvar1962 < (1'h1)); forvar1962 = (forvar1962 + (1'h1)))
                    begin
                      reg1963 <= reg347[(3'h4):(2'h2)];
                      reg1964 = $unsigned((reg320[(3'h5):(1'h0)] >>> $unsigned("Tyd8rAy")));
                      reg1965 = (&reg1952);
                      reg1966 <= wire1878;
                    end
                end
            end
        end
      reg1967 = reg307[(4'ha):(4'h9)];
    end
  assign wire1968 = reg357;
  module358 #() modinst1970 (.wire360(wire1876), .y(wire1969), .wire363(wire1234), .wire359(wire1874), .clk(clk), .wire362(reg322), .wire361(reg1945));
  assign wire1971 = (reg1963 ?
                        (+"ebF5d") : (~^((reg320 ?
                            wire1968 : reg1939) != (wire1878 ?
                            reg286 : reg1940))));
  assign wire1972 = reg1880;
  assign wire1973 = $signed(((|"p0mJ") ?
                        reg1905 : $signed($unsigned(reg1963))));
  assign wire1974 = reg1966;
  assign wire1975 = "UEsEfnbC";
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1235
#(parameter param1873 = (^((((8'h9f) >> (8'hb3)) ? (^~(8'hba)) : {(8'hb9)}) != (((8'hb9) << (8'hb1)) ? (^(8'ha0)) : ((8'hab) > (8'ha4))))))
(y, clk, wire1236, wire1237, wire1238, wire1239);
  output wire [(32'h2c9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire1236;
  input wire signed [(3'h6):(1'h0)] wire1237;
  input wire signed [(4'hd):(1'h0)] wire1238;
  input wire [(3'h5):(1'h0)] wire1239;
  wire signed [(4'h8):(1'h0)] wire1851;
  wire [(4'h9):(1'h0)] wire1240;
  wire [(4'h9):(1'h0)] wire1241;
  wire signed [(4'hd):(1'h0)] wire1245;
  wire signed [(5'h10):(1'h0)] wire1246;
  wire signed [(3'h5):(1'h0)] wire1290;
  wire [(4'h9):(1'h0)] wire1849;
  reg [(2'h3):(1'h0)] reg1870 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1868 = (1'h0);
  reg [(3'h7):(1'h0)] reg1854 = (1'h0);
  reg [(2'h2):(1'h0)] reg1283 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1282 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1278 = (1'h0);
  reg [(4'hf):(1'h0)] reg1275 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1274 = (1'h0);
  reg [(4'ha):(1'h0)] reg1271 = (1'h0);
  reg [(2'h3):(1'h0)] reg1270 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1264 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1261 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1260 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1251 = (1'h0);
  reg [(4'hf):(1'h0)] reg1256 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1247 = (1'h0);
  reg [(4'he):(1'h0)] reg1243 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1872 = (1'h0);
  reg [(4'hc):(1'h0)] reg1871 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1869 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1867 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1866 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1865 = (1'h0);
  reg [(3'h6):(1'h0)] reg1864 = (1'h0);
  reg [(2'h2):(1'h0)] reg1863 = (1'h0);
  reg [(3'h4):(1'h0)] reg1862 = (1'h0);
  reg [(4'he):(1'h0)] forvar1861 = (1'h0);
  reg [(4'h8):(1'h0)] reg1860 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1859 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1858 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1857 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1856 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1855 = (1'h0);
  reg [(4'hf):(1'h0)] reg1853 = (1'h0);
  reg [(4'hd):(1'h0)] reg1852 = (1'h0);
  reg [(4'hd):(1'h0)] reg1289 = (1'h0);
  reg [(4'he):(1'h0)] reg1288 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1287 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1286 = (1'h0);
  reg [(4'hd):(1'h0)] reg1285 = (1'h0);
  reg [(3'h5):(1'h0)] reg1284 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1281 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1280 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1279 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1277 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1276 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1273 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1272 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1269 = (1'h0);
  reg [(2'h2):(1'h0)] reg1268 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1267 = (1'h0);
  reg [(3'h4):(1'h0)] reg1266 = (1'h0);
  reg [(4'h9):(1'h0)] reg1265 = (1'h0);
  reg [(4'hc):(1'h0)] reg1263 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1262 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1259 = (1'h0);
  reg [(4'hc):(1'h0)] reg1258 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1257 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1252 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1249 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1253 = (1'h0);
  reg [(5'h10):(1'h0)] reg1255 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1254 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1253 = (1'h0);
  reg [(4'he):(1'h0)] reg1252 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1251 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1250 = (1'h0);
  reg [(4'hd):(1'h0)] reg1249 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1248 = (1'h0);
  reg [(4'hc):(1'h0)] reg1244 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1242 = (1'h0);
  assign y = {wire1851,
                 wire1849,
                 reg1854,
                 reg1282,
                 reg1278,
                 reg1260,
                 reg1256,
                 reg1247,
                 reg1863,
                 reg1862,
                 reg1860,
                 reg1859,
                 forvar1858,
                 forvar1855,
                 reg1852,
                 reg1289,
                 forvar1287,
                 forvar1281,
                 forvar1277,
                 forvar1269,
                 reg1268,
                 reg1266,
                 reg1265,
                 reg1257,
                 forvar1252,
                 forvar1249,
                 reg1254,
                 reg1253,
                 forvar1251,
                 (1'h0)};
  assign wire1240 = wire1239[(1'h0):(1'h0)];
  assign wire1241 = "PhQWViM2";
  always
    @(posedge clk) begin
      reg1242 = (^($unsigned((~^(8'ha8))) ?
          {$unsigned(wire1239)} : wire1241[(3'h5):(3'h4)]));
    end
  always
    @(posedge clk) begin
      reg1243 <= ($unsigned(wire1240[(4'h8):(2'h3)]) + $signed($unsigned((~^wire1237))));
      reg1244 = wire1241;
    end
  assign wire1245 = wire1237;
  assign wire1246 = "DPV";
  always
    @(posedge clk) begin
      reg1247 <= wire1239;
      if ("QqLvl")
        begin
          for (forvar1248 = (1'h0); (forvar1248 < (1'h1)); forvar1248 = (forvar1248 + (1'h1)))
            begin
              if ("i3z")
                begin
                  reg1249 = {(8'hb3)};
                end
              else
                begin
                  reg1249 = $signed(("r2Cm55dENY" ~^ ""));
                  reg1250 = $signed(reg1247[(3'h7):(2'h2)]);
                end
            end
          for (forvar1251 = (1'h0); (forvar1251 < (2'h3)); forvar1251 = (forvar1251 + (1'h1)))
            begin
              reg1252 = $unsigned((8'hb9));
              if (reg1252[(4'h9):(2'h2)])
                begin
                  reg1253 = (wire1239 ^ $unsigned(((wire1239 ?
                      reg1247 : reg1250) * "40lCcZEgWgvt")));
                  reg1254 = $unsigned($signed(forvar1248));
                  reg1255 = wire1245[(4'hc):(1'h0)];
                end
              else
                begin
                  for (forvar1253 = (1'h0); (forvar1253 < (1'h0)); forvar1253 = (forvar1253 + (1'h1)))
                    begin
                      reg1254 = (^({(^~forvar1253)} - $signed(wire1237[(2'h3):(2'h3)])));
                      reg1255 = wire1236[(3'h5):(3'h4)];
                      reg1256 <= ($unsigned({(forvar1251 ?
                              wire1239 : (8'hb4))}) != $signed(wire1237));
                    end
                end
            end
        end
      else
        begin
          for (forvar1248 = (1'h0); (forvar1248 < (1'h0)); forvar1248 = (forvar1248 + (1'h1)))
            begin
              for (forvar1249 = (1'h0); (forvar1249 < (1'h1)); forvar1249 = (forvar1249 + (1'h1)))
                begin
                  reg1251 <= (reg1247 + $unsigned({wire1236}));
                end
              for (forvar1252 = (1'h0); (forvar1252 < (1'h0)); forvar1252 = (forvar1252 + (1'h1)))
                begin
                  reg1253 = (8'ha2);
                end
              if (forvar1253[(1'h1):(1'h1)])
                begin
                  reg1256 <= (!(8'ha0));
                end
              else
                begin
                  if ((|({$unsigned(forvar1249)} ~^ wire1241)))
                    begin
                      reg1256 <= "JMCKCRP7cstQ1";
                      reg1257 = {(wire1245 << "7vMD3X")};
                      reg1258 = wire1239[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1254 = {(^~$signed(wire1241))};
                      reg1256 <= (wire1239 << "Jl8rUZldEeNi4eP");
                    end
                  for (forvar1259 = (1'h0); (forvar1259 < (1'h0)); forvar1259 = (forvar1259 + (1'h1)))
                    begin
                      reg1260 <= $unsigned($unsigned(forvar1253));
                      reg1261 <= (($unsigned((-forvar1248)) ?
                              $unsigned(reg1254[(3'h4):(2'h3)]) : wire1240) ?
                          ((wire1241 ?
                                  reg1247 : (reg1260 ? wire1236 : forvar1252)) ?
                              ($signed((8'hb6)) ?
                                  $unsigned(reg1243) : "8wS3p") : (reg1243[(4'hb):(2'h2)] ?
                                  reg1247 : (wire1240 ?
                                      (8'hb5) : wire1240))) : (8'ha2));
                    end
                  for (forvar1262 = (1'h0); (forvar1262 < (1'h1)); forvar1262 = (forvar1262 + (1'h1)))
                    begin
                      reg1263 = (forvar1248[(1'h1):(1'h1)] ^~ (reg1247 ?
                          ((~^(8'hb6)) + (reg1249 >= forvar1251)) : reg1257[(4'h9):(1'h0)]));
                      reg1264 <= reg1255;
                      reg1265 = {$unsigned(($signed(reg1243) ?
                              (forvar1259 <= (8'hba)) : (&reg1257)))};
                    end
                end
            end
          reg1266 = (^reg1249[(3'h5):(3'h4)]);
          for (forvar1267 = (1'h0); (forvar1267 < (2'h3)); forvar1267 = (forvar1267 + (1'h1)))
            begin
              reg1268 = forvar1252;
              for (forvar1269 = (1'h0); (forvar1269 < (1'h1)); forvar1269 = (forvar1269 + (1'h1)))
                begin
                  if ($signed({({wire1240} ? (^reg1250) : (+wire1236))}))
                    begin
                      reg1270 <= $unsigned(($signed($unsigned(reg1255)) ?
                          forvar1248[(1'h0):(1'h0)] : forvar1248));
                    end
                  else
                    begin
                      reg1270 <= $unsigned(reg1263[(4'hb):(3'h6)]);
                      reg1271 <= forvar1259;
                      reg1272 = "3creRxNJmEU3OX";
                    end
                  for (forvar1273 = (1'h0); (forvar1273 < (2'h3)); forvar1273 = (forvar1273 + (1'h1)))
                    begin
                      reg1274 <= (reg1250[(3'h4):(1'h1)] <= (!reg1265));
                      reg1275 <= $unsigned($signed(((|reg1272) == wire1239[(2'h2):(2'h2)])));
                    end
                  reg1276 = reg1252[(2'h3):(2'h2)];
                end
              for (forvar1277 = (1'h0); (forvar1277 < (1'h0)); forvar1277 = (forvar1277 + (1'h1)))
                begin
                  reg1278 <= reg1257;
                end
            end
        end
      for (forvar1279 = (1'h0); (forvar1279 < (1'h0)); forvar1279 = (forvar1279 + (1'h1)))
        begin
          for (forvar1280 = (1'h0); (forvar1280 < (2'h2)); forvar1280 = (forvar1280 + (1'h1)))
            begin
              for (forvar1281 = (1'h0); (forvar1281 < (2'h3)); forvar1281 = (forvar1281 + (1'h1)))
                begin
                  if (reg1266)
                    begin
                      reg1282 <= ({{"Jos"}} >= {(-(reg1265 >> forvar1251))});
                      reg1283 <= ("4sC" ? (~^(^$unsigned(wire1246))) : "VlRP1");
                      reg1284 = (|($signed($signed(reg1251)) ^ (reg1256 ?
                          (wire1237 ?
                              reg1260 : wire1240) : ((8'hb9) & reg1271))));
                    end
                  else
                    begin
                      reg1284 = {((~^{reg1265}) ?
                              (reg1249 ^ wire1237[(1'h1):(1'h1)]) : "55")};
                      reg1285 = reg1263[(4'hc):(3'h4)];
                    end
                end
            end
          for (forvar1286 = (1'h0); (forvar1286 < (2'h3)); forvar1286 = (forvar1286 + (1'h1)))
            begin
              for (forvar1287 = (1'h0); (forvar1287 < (1'h1)); forvar1287 = (forvar1287 + (1'h1)))
                begin
                  reg1288 = wire1239[(3'h5):(3'h4)];
                end
            end
          reg1289 = (8'hb6);
        end
    end
  assign wire1290 = wire1239[(3'h5):(1'h1)];
  module1291 #() modinst1850 (.wire1293(reg1260), .wire1296(reg1261), .wire1295(reg1256), .wire1294(wire1238), .wire1292(reg1247), .clk(clk), .y(wire1849));
  assign wire1851 = reg1274;
  always
    @(posedge clk) begin
      reg1852 = $unsigned((~^(~&(wire1237 ? (8'hae) : (8'hab)))));
      if ($unsigned($signed(reg1260)))
        begin
          reg1853 = "X";
        end
      else
        begin
          reg1854 <= (|$signed($unsigned(((8'hb2) ? reg1251 : reg1282))));
          for (forvar1855 = (1'h0); (forvar1855 < (1'h1)); forvar1855 = (forvar1855 + (1'h1)))
            begin
              for (forvar1856 = (1'h0); (forvar1856 < (2'h2)); forvar1856 = (forvar1856 + (1'h1)))
                begin
                  reg1857 = (~^($signed($unsigned(reg1270)) ?
                      $unsigned($unsigned(reg1270)) : reg1271));
                end
              for (forvar1858 = (1'h0); (forvar1858 < (1'h1)); forvar1858 = (forvar1858 + (1'h1)))
                begin
                  reg1859 = $unsigned(wire1246[(4'h8):(2'h2)]);
                  reg1860 = ($signed(({reg1270} == (forvar1858 ?
                      wire1241 : reg1275))) ~^ ((&{reg1278}) + $unsigned({(8'h9e)})));
                  for (forvar1861 = (1'h0); (forvar1861 < (2'h3)); forvar1861 = (forvar1861 + (1'h1)))
                    begin
                      reg1862 = "YZtJrW7NLGqv5";
                      reg1863 = ((((wire1236 ^ reg1270) ?
                              ((8'h9d) ?
                                  reg1862 : reg1251) : {wire1849}) - $signed(wire1238)) ?
                          reg1862 : $unsigned($unsigned($unsigned(wire1239))));
                      reg1864 = $signed(forvar1858[(3'h5):(3'h4)]);
                    end
                end
              for (forvar1865 = (1'h0); (forvar1865 < (1'h1)); forvar1865 = (forvar1865 + (1'h1)))
                begin
                  for (forvar1866 = (1'h0); (forvar1866 < (2'h2)); forvar1866 = (forvar1866 + (1'h1)))
                    begin
                      reg1867 = $unsigned(((wire1245 ?
                          $signed((8'hb5)) : {forvar1861}) >= ((reg1264 ?
                              (8'haf) : reg1854) ?
                          (+reg1247) : (&reg1270))));
                      reg1868 <= (reg1852[(3'h5):(1'h0)] * wire1237);
                    end
                  for (forvar1869 = (1'h0); (forvar1869 < (2'h3)); forvar1869 = (forvar1869 + (1'h1)))
                    begin
                      reg1870 <= "H7VQlS3VH";
                      reg1871 = (-"IlH8qTNnKtOCet");
                    end
                end
            end
          reg1872 = $signed(((reg1261 ? reg1282 : $unsigned(reg1261)) ?
              $unsigned((reg1857 ?
                  wire1290 : reg1256)) : (wire1240 ^~ (reg1862 * reg1867))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module358
#(parameter param1231 = ((8'hac) & (^(^((8'hb8) - (8'ha7))))))
(y, clk, wire359, wire360, wire361, wire362, wire363);
  output wire [(32'h5b7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire359;
  input wire signed [(4'hf):(1'h0)] wire360;
  input wire signed [(2'h2):(1'h0)] wire361;
  input wire signed [(4'hf):(1'h0)] wire362;
  input wire [(4'he):(1'h0)] wire363;
  wire [(3'h5):(1'h0)] wire1136;
  wire signed [(4'hb):(1'h0)] wire364;
  wire signed [(4'ha):(1'h0)] wire498;
  wire signed [(4'he):(1'h0)] wire543;
  wire [(4'ha):(1'h0)] wire1134;
  reg signed [(5'h10):(1'h0)] reg1215 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1227 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1220 = (1'h0);
  reg [(3'h5):(1'h0)] reg1218 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1217 = (1'h0);
  reg [(4'h9):(1'h0)] reg1212 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1210 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1209 = (1'h0);
  reg [(3'h6):(1'h0)] reg1207 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1202 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1203 = (1'h0);
  reg [(3'h4):(1'h0)] reg1200 = (1'h0);
  reg [(3'h4):(1'h0)] reg1199 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1194 = (1'h0);
  reg [(2'h3):(1'h0)] reg1193 = (1'h0);
  reg [(3'h5):(1'h0)] reg1190 = (1'h0);
  reg [(3'h7):(1'h0)] reg1186 = (1'h0);
  reg [(4'h9):(1'h0)] reg1184 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1182 = (1'h0);
  reg [(3'h7):(1'h0)] reg1181 = (1'h0);
  reg [(4'hc):(1'h0)] reg1179 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1175 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1174 = (1'h0);
  reg [(3'h6):(1'h0)] reg1173 = (1'h0);
  reg [(3'h5):(1'h0)] reg1168 = (1'h0);
  reg [(2'h3):(1'h0)] reg1161 = (1'h0);
  reg [(4'hc):(1'h0)] reg1160 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1159 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1147 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1158 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1154 = (1'h0);
  reg [(4'hf):(1'h0)] reg1152 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1149 = (1'h0);
  reg [(4'hc):(1'h0)] reg1140 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1142 = (1'h0);
  reg [(5'h10):(1'h0)] reg1145 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1143 = (1'h0);
  reg [(4'h8):(1'h0)] reg502 = (1'h0);
  reg [(4'hd):(1'h0)] reg503 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg515 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg520 = (1'h0);
  reg [(4'hd):(1'h0)] reg523 = (1'h0);
  reg [(4'hf):(1'h0)] reg525 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg526 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg527 = (1'h0);
  reg [(2'h3):(1'h0)] reg528 = (1'h0);
  reg signed [(4'he):(1'h0)] reg529 = (1'h0);
  reg signed [(4'he):(1'h0)] reg530 = (1'h0);
  reg [(3'h4):(1'h0)] reg534 = (1'h0);
  reg [(4'ha):(1'h0)] reg539 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1217 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1216 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1230 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1229 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1229 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1228 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1226 = (1'h0);
  reg [(3'h7):(1'h0)] reg1225 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1224 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1223 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1222 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1221 = (1'h0);
  reg [(4'hb):(1'h0)] reg1219 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1216 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1215 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1214 = (1'h0);
  reg [(4'h9):(1'h0)] reg1213 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1211 = (1'h0);
  reg [(4'hb):(1'h0)] reg1208 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1201 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1199 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1196 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1188 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1187 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1208 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1206 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1200 = (1'h0);
  reg [(2'h3):(1'h0)] reg1195 = (1'h0);
  reg [(2'h3):(1'h0)] reg1205 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1204 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1202 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1201 = (1'h0);
  reg [(3'h7):(1'h0)] reg1198 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1197 = (1'h0);
  reg [(2'h2):(1'h0)] reg1196 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1195 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1192 = (1'h0);
  reg [(4'ha):(1'h0)] reg1191 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1189 = (1'h0);
  reg [(2'h3):(1'h0)] reg1188 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1187 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1185 = (1'h0);
  reg [(4'h9):(1'h0)] reg1183 = (1'h0);
  reg [(4'h8):(1'h0)] reg1180 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1179 = (1'h0);
  reg [(3'h4):(1'h0)] reg1178 = (1'h0);
  reg [(2'h2):(1'h0)] reg1177 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1176 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1175 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1172 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1171 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1170 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1169 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1159 = (1'h0);
  reg [(4'ha):(1'h0)] reg1167 = (1'h0);
  reg [(4'hd):(1'h0)] reg1166 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1165 = (1'h0);
  reg [(2'h3):(1'h0)] reg1164 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1163 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1162 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1148 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1145 = (1'h0);
  reg [(3'h7):(1'h0)] reg1157 = (1'h0);
  reg [(4'hd):(1'h0)] reg1156 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1155 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1153 = (1'h0);
  reg [(4'hc):(1'h0)] reg1151 = (1'h0);
  reg [(3'h4):(1'h0)] reg1150 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1148 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1147 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1141 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1146 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1144 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1142 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1141 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1140 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1139 = (1'h0);
  reg [(3'h5):(1'h0)] reg1138 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1137 = (1'h0);
  reg [(4'h9):(1'h0)] reg542 = (1'h0);
  reg [(4'hd):(1'h0)] reg541 = (1'h0);
  reg signed [(4'he):(1'h0)] reg540 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar538 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg537 = (1'h0);
  reg [(4'hd):(1'h0)] reg536 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg535 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg533 = (1'h0);
  reg [(4'hb):(1'h0)] forvar532 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg531 = (1'h0);
  reg [(4'hf):(1'h0)] forvar524 = (1'h0);
  reg [(3'h7):(1'h0)] reg517 = (1'h0);
  reg [(5'h10):(1'h0)] forvar513 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg522 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg521 = (1'h0);
  reg [(4'hd):(1'h0)] reg519 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg518 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar517 = (1'h0);
  reg [(3'h4):(1'h0)] reg516 = (1'h0);
  reg [(4'h8):(1'h0)] forvar514 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg513 = (1'h0);
  reg [(3'h4):(1'h0)] reg512 = (1'h0);
  reg [(4'hb):(1'h0)] reg511 = (1'h0);
  reg [(3'h7):(1'h0)] reg510 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar509 = (1'h0);
  reg [(4'ha):(1'h0)] reg508 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg507 = (1'h0);
  reg [(4'hc):(1'h0)] reg506 = (1'h0);
  reg [(2'h3):(1'h0)] reg505 = (1'h0);
  reg [(4'ha):(1'h0)] forvar504 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar501 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar500 = (1'h0);
  assign y = {wire364,
                 wire498,
                 reg1215,
                 reg1220,
                 reg1218,
                 reg1207,
                 reg1203,
                 reg1200,
                 reg1199,
                 reg1193,
                 reg1190,
                 reg1179,
                 reg1175,
                 reg1173,
                 reg1160,
                 reg1147,
                 reg1152,
                 reg1145,
                 reg1143,
                 reg502,
                 reg515,
                 reg526,
                 reg534,
                 reg1230,
                 reg1229,
                 reg1226,
                 forvar1221,
                 reg1214,
                 reg1213,
                 reg1201,
                 forvar1199,
                 forvar1196,
                 forvar1188,
                 reg1187,
                 forvar1208,
                 reg1206,
                 reg1205,
                 reg1204,
                 reg1198,
                 reg1196,
                 forvar1195,
                 reg1192,
                 reg1191,
                 reg1185,
                 reg1180,
                 forvar1179,
                 reg1178,
                 reg1177,
                 reg1176,
                 forvar1175,
                 reg1172,
                 reg1169,
                 forvar1159,
                 reg1162,
                 forvar1148,
                 reg1157,
                 reg1153,
                 reg1148,
                 forvar1147,
                 reg1139,
                 reg542,
                 reg541,
                 reg540,
                 reg533,
                 forvar532,
                 reg517,
                 reg522,
                 forvar517,
                 reg507,
                 reg506,
                 forvar501,
                 (1'h0)};
  assign wire364 = wire360;
  module365 #() modinst499 (wire498, clk, wire364, wire359, wire362, wire360);
  always
    @(posedge clk) begin
      for (forvar500 = (1'h0); (forvar500 < (2'h3)); forvar500 = (forvar500 + (1'h1)))
        begin
          for (forvar501 = (1'h0); (forvar501 < (2'h3)); forvar501 = (forvar501 + (1'h1)))
            begin
              reg502 <= $unsigned($unsigned("r4CTNFu880"));
              reg503 <= wire362[(4'hb):(1'h0)];
              for (forvar504 = (1'h0); (forvar504 < (1'h1)); forvar504 = (forvar504 + (1'h1)))
                begin
                  if ($unsigned(((wire360[(4'h9):(2'h3)] ?
                          reg503 : (+forvar501)) ?
                      (wire498[(4'ha):(1'h1)] - (~^wire362)) : reg502[(1'h1):(1'h1)])))
                    begin
                      reg505 = (^$unsigned((|$signed(wire498))));
                      reg506 = (|(((wire498 >= wire362) ?
                          $signed(wire361) : $unsigned((8'ha6))) ~^ $signed((-(8'ha7)))));
                      reg507 = wire363[(3'h7):(2'h3)];
                      reg508 = ({(8'ha4)} + reg502);
                    end
                  else
                    begin
                      reg505 = ((+reg507) ?
                          wire364 : $unsigned($unsigned(((8'hb8) ?
                              wire361 : reg505))));
                      reg506 = wire359;
                    end
                end
            end
          for (forvar509 = (1'h0); (forvar509 < (2'h2)); forvar509 = (forvar509 + (1'h1)))
            begin
              reg510 = (^wire361);
              reg511 = wire363;
            end
          reg512 = (+($unsigned((~&(8'hb9))) > $signed((reg506 >>> wire359))));
          if (((wire498 ? reg502 : forvar509[(1'h1):(1'h0)]) ?
              wire364 : {((^reg506) & $signed(wire361))}))
            begin
              if (((wire364[(3'h6):(1'h1)] ?
                      reg510[(3'h7):(2'h2)] : ($unsigned((8'hb7)) & (reg505 ?
                          wire362 : reg508))) ?
                  (~&forvar500) : wire363[(2'h3):(2'h2)]))
                begin
                  reg513 = $unsigned((~|$unsigned({forvar509})));
                end
              else
                begin
                  reg513 = forvar504;
                  for (forvar514 = (1'h0); (forvar514 < (1'h1)); forvar514 = (forvar514 + (1'h1)))
                    begin
                      reg515 <= reg508;
                      reg516 = wire360;
                    end
                  for (forvar517 = (1'h0); (forvar517 < (1'h0)); forvar517 = (forvar517 + (1'h1)))
                    begin
                      reg518 = ($unsigned(($unsigned(reg513) >>> $unsigned(reg508))) ?
                          "lffvTGy2h" : $unsigned(($unsigned(wire363) ^~ {(8'hb1)})));
                    end
                  if ((({"398LguZa"} ?
                          ((forvar501 ? wire360 : reg515) ?
                              (reg516 && reg503) : (~&reg503)) : wire359[(3'h5):(1'h0)]) ?
                      (wire361 | ((~&forvar504) ?
                          (reg515 ?
                              wire364 : wire498) : reg503[(4'hc):(3'h5)])) : ($unsigned(reg516) + (^~$signed(wire363)))))
                    begin
                      reg519 = (($unsigned(reg505) ~^ reg513[(3'h5):(2'h3)]) - ((^(reg508 != reg515)) << "VJv2O"));
                      reg520 <= "ittc";
                    end
                  else
                    begin
                      reg519 = (($unsigned($signed((8'hb0))) ?
                              wire363 : reg512[(1'h1):(1'h1)]) ?
                          ($unsigned((^~reg505)) ?
                              reg519[(4'hd):(3'h5)] : $signed({reg520})) : "X");
                      reg521 = $unsigned("WshSybrdFM");
                    end
                end
              reg522 = forvar514;
            end
          else
            begin
              for (forvar513 = (1'h0); (forvar513 < (1'h1)); forvar513 = (forvar513 + (1'h1)))
                begin
                  for (forvar514 = (1'h0); (forvar514 < (2'h2)); forvar514 = (forvar514 + (1'h1)))
                    begin
                      reg515 <= reg503;
                      reg516 = "d8fELx6CDv";
                      reg517 = (&wire498[(4'h8):(1'h0)]);
                    end
                end
              reg520 <= $signed({("Zdn3mbvNQdmMSaI" ?
                      $signed(forvar514) : wire360[(4'h9):(1'h1)])});
              reg523 <= forvar504;
              if (forvar514)
                begin
                  for (forvar524 = (1'h0); (forvar524 < (2'h3)); forvar524 = (forvar524 + (1'h1)))
                    begin
                      reg525 <= ($unsigned(reg511[(1'h1):(1'h1)]) && reg517);
                      reg526 <= $unsigned($unsigned({{wire498}}));
                      reg527 <= (~&(((reg526 ? forvar514 : (8'haf)) ?
                              (forvar504 ?
                                  reg511 : (8'hac)) : (wire363 ~^ reg513)) ?
                          $unsigned("3OyWMeG") : (~^$signed(reg522))));
                    end
                  reg528 <= wire364[(1'h0):(1'h0)];
                  if ((~("uIYIwHWRlH6Qwb" ?
                      ($unsigned(reg516) > (&wire498)) : wire360)))
                    begin
                      reg529 <= (&(wire360 ? reg519 : wire362[(4'hc):(3'h7)]));
                      reg530 <= (-reg517);
                    end
                  else
                    begin
                      reg529 <= reg507;
                      reg531 = (forvar513[(3'h5):(1'h0)] ^ (wire360 ?
                          (((8'had) >>> reg507) ?
                              (reg525 >= forvar509) : "6k") : (+reg515)));
                    end
                end
              else
                begin
                  for (forvar524 = (1'h0); (forvar524 < (1'h1)); forvar524 = (forvar524 + (1'h1)))
                    begin
                      reg531 = (((~&$unsigned(reg525)) ~^ (+((8'hab) <= wire360))) ?
                          $unsigned(forvar517) : ((8'hac) ?
                              $signed({reg505}) : ((reg527 ?
                                  reg502 : reg517) && (!wire361))));
                    end
                  for (forvar532 = (1'h0); (forvar532 < (1'h0)); forvar532 = (forvar532 + (1'h1)))
                    begin
                      reg533 = ((reg531 ?
                          $unsigned("8mtxVmit") : (|(reg529 ?
                              reg530 : reg502))) >> $signed(reg508[(3'h4):(2'h3)]));
                      reg534 <= (forvar500 >>> reg503);
                      reg535 = "CWp6POLh4O7mRP";
                      reg536 = $signed("");
                    end
                  reg537 = (^"J2pBSqX");
                  for (forvar538 = (1'h0); (forvar538 < (1'h0)); forvar538 = (forvar538 + (1'h1)))
                    begin
                      reg539 <= "2PayaFF8ZMenle";
                      reg540 = reg534[(1'h0):(1'h0)];
                      reg541 = {$unsigned($unsigned(reg508[(2'h2):(1'h1)]))};
                    end
                end
            end
        end
      reg542 = ($signed(reg529) ?
          $unsigned(forvar504[(3'h6):(3'h6)]) : (^~"FbV58BM45pe1rG"));
    end
  assign wire543 = $signed(reg502);
  module544 #() modinst1135 (wire1134, clk, wire543, reg529, reg527, reg502);
  assign wire1136 = $signed(reg529);
  always
    @(posedge clk) begin
      for (forvar1137 = (1'h0); (forvar1137 < (2'h2)); forvar1137 = (forvar1137 + (1'h1)))
        begin
          reg1138 = $signed($unsigned((8'hb5)));
        end
      if ({(+"a")})
        begin
          if (((8'ha5) ?
              ((^((8'h9e) * wire359)) && $unsigned("")) : $signed("iub")))
            begin
              reg1139 = (((^~(!wire1134)) <<< ($signed(reg523) >> (reg520 && reg539))) ?
                  wire498 : reg534);
              for (forvar1140 = (1'h0); (forvar1140 < (2'h2)); forvar1140 = (forvar1140 + (1'h1)))
                begin
                  reg1141 = $unsigned((($signed(wire498) ?
                      $unsigned((8'ha2)) : (reg523 * reg503)) >> ((reg534 ?
                          reg503 : wire362) ?
                      $signed((8'ha1)) : (wire360 != reg503))));
                end
              if (((~&($unsigned(wire361) ?
                  $unsigned(wire363) : $signed(reg502))) || $signed(("6GG" != $unsigned(wire1136)))))
                begin
                  for (forvar1142 = (1'h0); (forvar1142 < (2'h3)); forvar1142 = (forvar1142 + (1'h1)))
                    begin
                      reg1143 <= $signed(forvar1140);
                      reg1144 = wire359;
                    end
                  reg1145 <= {(~(^$unsigned(reg520)))};
                end
              else
                begin
                  reg1142 <= (reg1145[(4'hf):(1'h0)] | $signed($unsigned((wire498 - reg502))));
                  if ($unsigned("rk"))
                    begin
                      reg1144 = $signed($unsigned({wire1134[(3'h5):(2'h2)]}));
                      reg1145 <= $signed($signed(($signed(wire1134) | reg1145)));
                      reg1146 = wire498[(4'h9):(1'h0)];
                    end
                  else
                    begin
                      reg1143 <= $signed((~^(wire364 ?
                          (wire361 ?
                              reg1141 : reg1143) : wire498[(2'h3):(2'h3)])));
                      reg1145 <= {(~$signed("4AhrlyhV"))};
                      reg1146 = (wire361 ^~ (reg1146[(4'ha):(3'h4)] <<< $unsigned(((8'hab) + reg1139))));
                    end
                end
            end
          else
            begin
              reg1140 <= "2bMqm4g3Qwo9cXB";
            end
        end
      else
        begin
          reg1140 <= $unsigned($unsigned(wire362[(2'h2):(1'h1)]));
          for (forvar1141 = (1'h0); (forvar1141 < (1'h0)); forvar1141 = (forvar1141 + (1'h1)))
            begin
              for (forvar1142 = (1'h0); (forvar1142 < (2'h3)); forvar1142 = (forvar1142 + (1'h1)))
                begin
                  reg1144 = (($signed($unsigned(wire1134)) >>> (-$unsigned(wire364))) ?
                      $signed("06fJ2cDs") : (((reg520 & (8'hab)) <<< $unsigned(reg1144)) ?
                          $signed($signed((8'hac))) : $unsigned($unsigned(reg1138))));
                end
              if (((((reg515 ? reg1141 : forvar1141) ?
                      (+reg529) : (wire364 < reg523)) ?
                  reg530 : reg525[(4'hc):(4'h8)]) & $signed($signed((~reg1142)))))
                begin
                  reg1146 = (~^(wire498 == ((^~(8'hb8)) ?
                      (wire360 - reg530) : (reg503 <<< forvar1141))));
                  for (forvar1147 = (1'h0); (forvar1147 < (1'h1)); forvar1147 = (forvar1147 + (1'h1)))
                    begin
                      reg1148 = reg1144[(1'h0):(1'h0)];
                      reg1149 <= ("KP7MVJwy" >= {((reg530 * reg502) ?
                              (|reg534) : $unsigned((8'hb2)))});
                      reg1150 = "oQHA";
                    end
                  if (({((wire361 ?
                          wire1136 : wire362) >>> (reg1145 ^ reg525))} >>> $signed($unsigned(reg526[(4'hb):(4'h9)]))))
                    begin
                      reg1151 = reg1140[(3'h4):(1'h1)];
                      reg1152 <= (-(~((reg529 ? reg539 : (8'haf)) | (reg1143 ?
                          reg1139 : (8'hba)))));
                      reg1153 = reg529;
                    end
                  else
                    begin
                      reg1151 = $signed({(reg529 ^~ $unsigned(reg1139))});
                      reg1153 = wire1134[(3'h5):(3'h5)];
                      reg1154 <= reg1140;
                    end
                  if ((~|"6QVolCL4bNrF"))
                    begin
                      reg1155 = ("dVtP6Fz85y" ?
                          ($signed($signed(wire361)) <<< (~(reg526 ?
                              reg530 : reg539))) : (reg1142[(3'h5):(3'h5)] ~^ "HyIc177oHfpQd0"));
                      reg1156 = (wire361 ?
                          (wire1134[(1'h1):(1'h1)] == (forvar1141[(4'h8):(3'h5)] ?
                              "RYDln5eXfnC3Is" : reg1148)) : ("Eu2SX2gi" ?
                              wire1134[(4'ha):(2'h2)] : (&(-reg1146))));
                    end
                  else
                    begin
                      reg1155 = reg1153;
                      reg1156 = $signed(((reg1152 << (reg1140 > (8'h9d))) ?
                          ((!wire360) ?
                              "DoYGIeDqqJvkeT" : ((8'ha2) ?
                                  reg525 : forvar1147)) : $signed($signed(reg526))));
                      reg1157 = $unsigned((^~reg1154[(3'h7):(3'h4)]));
                      reg1158 <= (-reg1155[(2'h3):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar1145 = (1'h0); (forvar1145 < (2'h3)); forvar1145 = (forvar1145 + (1'h1)))
                    begin
                      reg1146 = $signed($signed(((+reg525) < (reg503 - reg1150))));
                      reg1147 <= ($signed(((reg1149 ^~ wire361) ?
                              reg1139 : (~&wire362))) ?
                          ((8'hba) ?
                              reg1142[(3'h5):(2'h3)] : (forvar1141 ?
                                  "HIY" : $signed(reg1149))) : $unsigned(($signed(reg525) ?
                              (forvar1147 ?
                                  reg526 : (8'hb5)) : $unsigned(reg1156))));
                    end
                  for (forvar1148 = (1'h0); (forvar1148 < (2'h3)); forvar1148 = (forvar1148 + (1'h1)))
                    begin
                      reg1150 = "";
                      reg1152 <= ($unsigned(((^~reg528) * reg529)) ?
                          "CwXTONGa0D9" : (~|$unsigned("49FGmifBs")));
                    end
                  reg1153 = "TrRioI";
                end
              if ($signed(reg1148[(4'ha):(1'h1)]))
                begin
                  reg1159 <= (^~reg502[(3'h6):(1'h1)]);
                  reg1160 <= (~&($unsigned(reg1153) && (~&(wire363 != reg534))));
                  if (reg1145[(2'h3):(2'h3)])
                    begin
                      reg1161 <= $unsigned((|forvar1147[(2'h3):(1'h0)]));
                      reg1162 = ((|((reg1159 <= reg1156) && $signed(reg502))) ?
                          $signed((reg1159[(3'h5):(2'h2)] ?
                              $unsigned(reg526) : wire359)) : $unsigned((forvar1147 ?
                              reg523[(3'h4):(2'h3)] : ((8'hb7) ?
                                  reg523 : reg1155))));
                      reg1163 = {$signed((reg539[(4'h9):(3'h7)] >= reg523))};
                    end
                  else
                    begin
                      reg1161 <= (reg1146[(1'h0):(1'h0)] || ((wire498[(4'ha):(3'h5)] >>> {reg1160}) < $unsigned(((8'ha8) ?
                          wire361 : reg515))));
                      reg1162 = $signed(reg1139);
                    end
                  if ({$unsigned($unsigned(reg1149))})
                    begin
                      reg1164 = $unsigned({$signed(wire364)});
                      reg1165 = wire1134;
                      reg1166 = reg526;
                      reg1167 = {({forvar1140} ?
                              reg1162[(1'h0):(1'h0)] : $unsigned($signed(reg1142)))};
                    end
                  else
                    begin
                      reg1164 = reg1162[(2'h2):(1'h0)];
                      reg1165 = "a77";
                    end
                end
              else
                begin
                  for (forvar1159 = (1'h0); (forvar1159 < (1'h0)); forvar1159 = (forvar1159 + (1'h1)))
                    begin
                      reg1162 = ((($unsigned(reg1166) ?
                          $unsigned(reg1165) : (forvar1137 == forvar1140)) > $unsigned(((8'hb7) ?
                          wire359 : forvar1147))) < reg1151);
                      reg1168 <= $unsigned(("TCdxSCP1EMa" | wire1136));
                      reg1169 = reg534[(2'h3):(1'h1)];
                    end
                  for (forvar1170 = (1'h0); (forvar1170 < (2'h2)); forvar1170 = (forvar1170 + (1'h1)))
                    begin
                      reg1171 = (reg1139 && wire362[(3'h4):(1'h0)]);
                      reg1172 = reg520[(4'h8):(2'h2)];
                      reg1173 <= {reg1171[(3'h7):(2'h3)]};
                    end
                  reg1174 <= $unsigned(((!(forvar1147 ? wire543 : reg1147)) ?
                      $unsigned($signed((8'haa))) : $signed((^~forvar1145))));
                end
              if ($unsigned(({(^~reg1142)} ? (~|{reg1144}) : "V8yiguUceidC")))
                begin
                  for (forvar1175 = (1'h0); (forvar1175 < (2'h3)); forvar1175 = (forvar1175 + (1'h1)))
                    begin
                      reg1176 = (~(reg1140 ? (8'hb9) : reg529[(3'h5):(1'h0)]));
                      reg1177 = reg1160;
                      reg1178 = ((reg520 * $signed((reg528 ?
                              (8'ha3) : reg1139))) ?
                          (8'had) : $signed(((reg539 ? reg528 : reg1141) ?
                              "bd" : {wire498})));
                    end
                  for (forvar1179 = (1'h0); (forvar1179 < (2'h3)); forvar1179 = (forvar1179 + (1'h1)))
                    begin
                      reg1180 = (~^"ds4pwAFLin");
                    end
                end
              else
                begin
                  reg1175 <= $unsigned(reg1144[(3'h4):(3'h4)]);
                  reg1179 <= "t7C";
                  reg1180 = forvar1170[(3'h4):(3'h4)];
                  if ((reg1179 ?
                      (($signed(wire364) ? (reg503 ^ reg1180) : {reg1179}) ?
                          ($unsigned(reg1164) - $unsigned(wire498)) : $unsigned((reg523 ?
                              (8'ha4) : reg523))) : {({(8'hb0)} || reg502[(3'h7):(3'h4)])}))
                    begin
                      reg1181 <= reg525[(4'hd):(1'h0)];
                      reg1182 <= $unsigned($signed(((reg529 ?
                              forvar1147 : reg1139) ?
                          (forvar1148 ?
                              wire364 : wire359) : (reg1164 <<< forvar1142))));
                      reg1183 = $unsigned(reg1148[(3'h5):(3'h4)]);
                      reg1184 <= wire1136;
                    end
                  else
                    begin
                      reg1181 <= reg515;
                      reg1182 <= reg503;
                      reg1183 = (({$unsigned(wire1134)} ?
                          (^(-reg1142)) : reg1141[(3'h4):(1'h0)]) - $signed($unsigned({(8'ha6)})));
                      reg1184 <= reg1153[(2'h2):(1'h0)];
                    end
                end
            end
        end
      reg1185 = "gbMMKtJmOrL5T04";
      if ($unsigned(reg520))
        begin
          reg1186 <= ($unsigned("6aO") ~^ (~|(~reg1168[(3'h5):(1'h1)])));
          for (forvar1187 = (1'h0); (forvar1187 < (2'h3)); forvar1187 = (forvar1187 + (1'h1)))
            begin
              reg1188 = ($signed($unsigned(reg1167)) > $unsigned({$unsigned(reg1169)}));
              for (forvar1189 = (1'h0); (forvar1189 < (2'h2)); forvar1189 = (forvar1189 + (1'h1)))
                begin
                  if ("mLVl")
                    begin
                      reg1190 <= "gG2N7uTSY8te9K";
                      reg1191 = (^~reg529[(3'h7):(3'h6)]);
                      reg1192 = ($unsigned(((!reg1191) <= reg539[(1'h0):(1'h0)])) & (|((wire361 != (8'ha5)) ?
                          reg1175 : (forvar1140 >= reg527))));
                    end
                  else
                    begin
                      reg1191 = (("1g4xHBDJS" ?
                              ({(8'ha4)} ?
                                  $unsigned(reg1188) : reg1192) : (!reg1153[(4'ha):(1'h1)])) ?
                          (+$unsigned(reg1192[(1'h0):(1'h0)])) : (("8mI6N3Udy" * (^reg502)) - {reg1176}));
                      reg1192 = reg1164[(1'h1):(1'h0)];
                      reg1193 <= forvar1159[(2'h2):(2'h2)];
                      reg1194 <= "dUcxud4FnExpi1b";
                    end
                  for (forvar1195 = (1'h0); (forvar1195 < (1'h0)); forvar1195 = (forvar1195 + (1'h1)))
                    begin
                      reg1196 = reg1161[(2'h2):(2'h2)];
                      reg1197 = ({(!reg526[(1'h0):(1'h0)])} ?
                          (^~(8'h9e)) : (((+(8'hb2)) <= reg1185) || $signed($unsigned(reg1160))));
                      reg1198 = forvar1145[(3'h7):(3'h4)];
                    end
                  reg1199 <= reg1160;
                  reg1200 <= reg1149[(4'hf):(4'ha)];
                end
              for (forvar1201 = (1'h0); (forvar1201 < (2'h2)); forvar1201 = (forvar1201 + (1'h1)))
                begin
                  for (forvar1202 = (1'h0); (forvar1202 < (2'h2)); forvar1202 = (forvar1202 + (1'h1)))
                    begin
                      reg1203 <= (~|{$unsigned((^wire363))});
                      reg1204 = "lI";
                    end
                end
            end
          reg1205 = "ha";
        end
      else
        begin
          if ((^~$unsigned(wire362[(2'h2):(1'h1)])))
            begin
              reg1186 <= (&reg1203[(3'h5):(3'h5)]);
              for (forvar1187 = (1'h0); (forvar1187 < (2'h2)); forvar1187 = (forvar1187 + (1'h1)))
                begin
                  reg1188 = ((+((reg1179 ? reg1172 : wire363) ?
                      reg1177 : $unsigned(reg526))) && $unsigned("lffrSMIO"));
                  for (forvar1189 = (1'h0); (forvar1189 < (1'h0)); forvar1189 = (forvar1189 + (1'h1)))
                    begin
                      reg1190 <= ($signed((~^(~|reg1181))) ?
                          $signed($unsigned((&wire498))) : reg1138[(1'h0):(1'h0)]);
                      reg1191 = (((-reg1163[(1'h0):(1'h0)]) ?
                          {reg526[(3'h5):(1'h0)]} : reg1160) == ($unsigned("gb") | (~&(+wire362))));
                      reg1193 <= ($unsigned({(~(8'ha3))}) * {($unsigned(reg1167) != reg1162[(3'h4):(2'h3)])});
                      reg1195 = wire498[(2'h3):(2'h3)];
                    end
                end
              reg1199 <= reg1169[(3'h6):(3'h4)];
              for (forvar1200 = (1'h0); (forvar1200 < (2'h3)); forvar1200 = (forvar1200 + (1'h1)))
                begin
                  for (forvar1201 = (1'h0); (forvar1201 < (2'h3)); forvar1201 = (forvar1201 + (1'h1)))
                    begin
                      reg1202 <= ((forvar1148 & {{(8'ha0)}}) >>> $unsigned(($signed((8'hb3)) ~^ {reg502})));
                      reg1204 = forvar1179;
                      reg1205 = $unsigned(wire543[(2'h3):(1'h0)]);
                      reg1206 = reg1185[(4'h8):(2'h3)];
                    end
                  reg1207 <= (reg1158 ?
                      (~(!$signed((8'ha7)))) : (((reg1194 ?
                                  forvar1187 : wire359) ?
                              (~reg1145) : (reg1180 || (8'ha5))) ?
                          {reg1203} : $unsigned($unsigned(forvar1200))));
                  for (forvar1208 = (1'h0); (forvar1208 < (1'h1)); forvar1208 = (forvar1208 + (1'h1)))
                    begin
                      reg1209 <= $unsigned((({reg1177} ~^ $signed(wire361)) ?
                          (~$signed(reg526)) : wire359[(4'he):(2'h3)]));
                    end
                end
            end
          else
            begin
              reg1187 = (^~(($unsigned(forvar1201) - reg1148) ?
                  reg1180 : "Fa"));
              for (forvar1188 = (1'h0); (forvar1188 < (1'h0)); forvar1188 = (forvar1188 + (1'h1)))
                begin
                  for (forvar1189 = (1'h0); (forvar1189 < (1'h0)); forvar1189 = (forvar1189 + (1'h1)))
                    begin
                      reg1191 = (8'hb0);
                    end
                  reg1193 <= reg1203;
                  if (reg1155)
                    begin
                      reg1194 <= "QwiTYe40kAf";
                      reg1195 = reg1142;
                    end
                  else
                    begin
                      reg1195 = $signed(($unsigned("pN4UBGZt") >>> reg1138));
                    end
                  for (forvar1196 = (1'h0); (forvar1196 < (2'h2)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 = "RMF0ER3VeCLp";
                      reg1198 = reg1187[(3'h4):(1'h0)];
                    end
                end
              for (forvar1199 = (1'h0); (forvar1199 < (2'h3)); forvar1199 = (forvar1199 + (1'h1)))
                begin
                  if ({{(8'haa)}})
                    begin
                      reg1200 <= ((|$unsigned((|reg1140))) ?
                          reg1194[(3'h4):(2'h2)] : "2Ka2EOQzCp94f");
                      reg1201 = $signed(((reg1153[(3'h4):(1'h0)] * forvar1188) ?
                          ((forvar1196 ?
                              forvar1189 : reg1178) * wire1136[(1'h1):(1'h0)]) : $unsigned(((8'hb2) ?
                              (8'haf) : reg1151))));
                      reg1202 <= $signed((wire498 ?
                          "UHLvl5QfMhyX3" : ({(8'hb9)} <<< reg1167[(3'h6):(1'h0)])));
                      reg1204 = "X6IXVsLlzuwoXiD";
                    end
                  else
                    begin
                      reg1201 = $signed(reg1148[(4'h8):(2'h2)]);
                      reg1204 = $unsigned("hnv8Lr5Qfff");
                      reg1207 <= (((^~forvar1142) ?
                              (8'hba) : $unsigned((reg1190 >> (8'hb0)))) ?
                          forvar1140 : (-((~reg534) <= reg1138)));
                      reg1208 = (8'h9c);
                    end
                  reg1209 <= $unsigned(($signed($signed(reg1174)) <<< reg1169[(4'h9):(1'h1)]));
                  reg1210 <= {(~&"daiu8s")};
                  for (forvar1211 = (1'h0); (forvar1211 < (2'h3)); forvar1211 = (forvar1211 + (1'h1)))
                    begin
                      reg1212 <= (|reg1161[(1'h1):(1'h1)]);
                      reg1213 = forvar1147;
                    end
                end
              reg1214 = {(!$signed((forvar1195 ? reg1141 : wire362)))};
            end
          if ((^~{reg1214[(3'h5):(1'h1)]}))
            begin
              for (forvar1215 = (1'h0); (forvar1215 < (2'h2)); forvar1215 = (forvar1215 + (1'h1)))
                begin
                  for (forvar1216 = (1'h0); (forvar1216 < (1'h1)); forvar1216 = (forvar1216 + (1'h1)))
                    begin
                      reg1217 <= (reg1196 ?
                          reg1142 : (($signed(reg1199) ?
                                  (reg1162 == reg1184) : (~^reg1165)) ?
                              ((reg1140 ?
                                  reg1196 : reg1161) != {reg1203}) : ((~reg525) | reg1188[(2'h2):(2'h2)])));
                      reg1218 <= $unsigned(reg1213);
                      reg1219 = (^(^("B60ISfSKAU8MtAA" ?
                          $signed(reg1161) : (forvar1189 ?
                              reg526 : forvar1140))));
                    end
                end
              reg1220 <= ($unsigned((+(~|forvar1147))) ?
                  ($unsigned((-reg1157)) ?
                      reg1180[(3'h4):(2'h3)] : ("7Qg1KNns" >> ((8'ha9) ?
                          (8'ha3) : forvar1179))) : (!forvar1211));
              for (forvar1221 = (1'h0); (forvar1221 < (1'h1)); forvar1221 = (forvar1221 + (1'h1)))
                begin
                  for (forvar1222 = (1'h0); (forvar1222 < (1'h1)); forvar1222 = (forvar1222 + (1'h1)))
                    begin
                      reg1223 = ((((^reg1190) <<< (reg1154 ?
                              reg1193 : reg1153)) ?
                          {(forvar1216 ?
                                  (8'hb5) : forvar1141)} : ($signed(reg1141) ?
                              (reg1144 ?
                                  reg1155 : reg1187) : reg1220[(4'he):(4'h8)])) >> ((&$unsigned((8'ha0))) ?
                          $signed((^reg1154)) : $signed((+(8'h9c)))));
                    end
                  for (forvar1224 = (1'h0); (forvar1224 < (1'h1)); forvar1224 = (forvar1224 + (1'h1)))
                    begin
                      reg1225 = (reg1191[(2'h3):(2'h3)] ?
                          ($unsigned((reg1152 ? forvar1140 : reg1173)) ?
                              reg1147 : "GWAh4QL") : (^{"Ron"}));
                      reg1226 = ((forvar1189 ?
                          ($signed(reg1168) == $signed(reg503)) : $unsigned((reg1172 ?
                              reg1171 : reg1203))) <<< reg1178[(1'h0):(1'h0)]);
                    end
                  reg1227 <= reg1159;
                  reg1228 = $unsigned($signed($unsigned(reg1174)));
                end
              if (wire1136[(3'h4):(3'h4)])
                begin
                  reg1229 = {($unsigned((~|reg1218)) ?
                          forvar1201[(2'h2):(2'h2)] : reg1188)};
                end
              else
                begin
                  for (forvar1229 = (1'h0); (forvar1229 < (2'h2)); forvar1229 = (forvar1229 + (1'h1)))
                    begin
                      reg1230 = $signed({$signed($unsigned(forvar1188))});
                    end
                end
            end
          else
            begin
              reg1215 <= reg1228;
              reg1216 = $signed((forvar1159 ?
                  $unsigned((wire362 >= wire543)) : "rY"));
              for (forvar1217 = (1'h0); (forvar1217 < (1'h0)); forvar1217 = (forvar1217 + (1'h1)))
                begin
                  reg1218 <= reg1202;
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module544
#(parameter param1133 = (~&(((~&(8'hac)) ? (-(8'ha4)) : ((8'had) && (8'h9c))) ? {{(8'hba)}} : (8'hb2))))
(y, clk, wire548, wire547, wire546, wire545);
  output wire [(32'h97e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire548;
  input wire [(3'h5):(1'h0)] wire547;
  input wire signed [(3'h6):(1'h0)] wire546;
  input wire [(4'h8):(1'h0)] wire545;
  wire [(5'h10):(1'h0)] wire1132;
  wire [(4'he):(1'h0)] wire977;
  wire signed [(2'h2):(1'h0)] wire650;
  wire [(3'h7):(1'h0)] wire649;
  wire signed [(5'h10):(1'h0)] wire648;
  wire signed [(4'hf):(1'h0)] wire647;
  wire signed [(4'ha):(1'h0)] wire645;
  wire signed [(2'h3):(1'h0)] wire619;
  wire [(4'ha):(1'h0)] wire549;
  reg signed [(4'hf):(1'h0)] reg1121 = (1'h0);
  reg [(5'h10):(1'h0)] reg1109 = (1'h0);
  reg [(4'he):(1'h0)] reg1103 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1129 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1115 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1114 = (1'h0);
  reg [(4'h8):(1'h0)] reg1113 = (1'h0);
  reg [(3'h6):(1'h0)] reg1110 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1105 = (1'h0);
  reg [(4'hf):(1'h0)] reg1085 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1075 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1100 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1099 = (1'h0);
  reg [(3'h4):(1'h0)] reg1097 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1094 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1088 = (1'h0);
  reg [(4'ha):(1'h0)] reg1087 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1086 = (1'h0);
  reg [(2'h3):(1'h0)] reg1083 = (1'h0);
  reg [(2'h2):(1'h0)] reg1082 = (1'h0);
  reg [(2'h2):(1'h0)] reg1079 = (1'h0);
  reg [(4'h8):(1'h0)] reg1077 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1072 = (1'h0);
  reg [(4'hb):(1'h0)] reg1071 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1062 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1069 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1057 = (1'h0);
  reg [(3'h5):(1'h0)] reg1056 = (1'h0);
  reg [(4'he):(1'h0)] reg1053 = (1'h0);
  reg [(3'h5):(1'h0)] reg1052 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1047 = (1'h0);
  reg [(4'hf):(1'h0)] reg1041 = (1'h0);
  reg [(3'h6):(1'h0)] reg1040 = (1'h0);
  reg [(2'h3):(1'h0)] reg1035 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1034 = (1'h0);
  reg [(3'h4):(1'h0)] reg1028 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1027 = (1'h0);
  reg [(2'h2):(1'h0)] reg1025 = (1'h0);
  reg [(3'h5):(1'h0)] reg1024 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1022 = (1'h0);
  reg [(2'h2):(1'h0)] reg1015 = (1'h0);
  reg [(4'he):(1'h0)] reg1007 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1005 = (1'h0);
  reg [(2'h3):(1'h0)] reg1002 = (1'h0);
  reg [(2'h3):(1'h0)] reg1001 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg998 = (1'h0);
  reg [(3'h4):(1'h0)] reg997 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg992 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg987 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg984 = (1'h0);
  reg [(3'h5):(1'h0)] reg983 = (1'h0);
  reg [(3'h6):(1'h0)] reg981 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg550 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg551 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg553 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg558 = (1'h0);
  reg [(4'hf):(1'h0)] reg561 = (1'h0);
  reg [(4'h9):(1'h0)] reg563 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg571 = (1'h0);
  reg [(2'h3):(1'h0)] reg579 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg577 = (1'h0);
  reg [(2'h2):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg585 = (1'h0);
  reg [(4'hc):(1'h0)] reg586 = (1'h0);
  reg [(4'hb):(1'h0)] reg590 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg575 = (1'h0);
  reg signed [(4'he):(1'h0)] reg583 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg598 = (1'h0);
  reg [(3'h6):(1'h0)] reg600 = (1'h0);
  reg [(4'hc):(1'h0)] reg608 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg612 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg616 = (1'h0);
  reg [(2'h2):(1'h0)] reg618 = (1'h0);
  reg [(2'h2):(1'h0)] reg1131 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1118 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1100 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1130 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1128 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1127 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1126 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1125 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1124 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1123 = (1'h0);
  reg [(2'h3):(1'h0)] reg1122 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1121 = (1'h0);
  reg [(4'he):(1'h0)] reg1120 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1119 = (1'h0);
  reg [(4'hd):(1'h0)] reg1118 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1117 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1116 = (1'h0);
  reg [(5'h10):(1'h0)] reg1112 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1111 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1112 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1111 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1109 = (1'h0);
  reg [(3'h5):(1'h0)] reg1108 = (1'h0);
  reg [(4'hb):(1'h0)] reg1107 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1106 = (1'h0);
  reg [(3'h6):(1'h0)] reg1104 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1103 = (1'h0);
  reg [(4'hd):(1'h0)] reg1102 = (1'h0);
  reg [(2'h3):(1'h0)] reg1101 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1096 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1091 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1081 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1080 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1077 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1076 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1072 = (1'h0);
  reg [(4'hf):(1'h0)] reg1073 = (1'h0);
  reg [(4'hf):(1'h0)] reg1098 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1096 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1095 = (1'h0);
  reg [(3'h5):(1'h0)] reg1093 = (1'h0);
  reg [(2'h2):(1'h0)] reg1092 = (1'h0);
  reg [(4'hc):(1'h0)] reg1091 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1090 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1089 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1085 = (1'h0);
  reg [(4'he):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1081 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1080 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1078 = (1'h0);
  reg [(2'h3):(1'h0)] reg1076 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1075 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1074 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1073 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1066 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1063 = (1'h0);
  reg [(2'h2):(1'h0)] reg1061 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1059 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1058 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1070 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1068 = (1'h0);
  reg [(4'hf):(1'h0)] reg1067 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1066 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1065 = (1'h0);
  reg [(4'hd):(1'h0)] reg1064 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1063 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1062 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1061 = (1'h0);
  reg [(4'hc):(1'h0)] reg1060 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1059 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1058 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1055 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1054 = (1'h0);
  reg [(2'h3):(1'h0)] reg1051 = (1'h0);
  reg [(4'hc):(1'h0)] reg1050 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1049 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1048 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1046 = (1'h0);
  reg [(4'hd):(1'h0)] reg1045 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1044 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1043 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1042 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1039 = (1'h0);
  reg [(3'h4):(1'h0)] reg1038 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1037 = (1'h0);
  reg [(2'h3):(1'h0)] reg1036 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1033 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1032 = (1'h0);
  reg [(2'h3):(1'h0)] reg1031 = (1'h0);
  reg [(3'h7):(1'h0)] reg1030 = (1'h0);
  reg [(4'h9):(1'h0)] reg1029 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1026 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1018 = (1'h0);
  reg [(3'h7):(1'h0)] reg1023 = (1'h0);
  reg [(4'h8):(1'h0)] reg1021 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1020 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1019 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1018 = (1'h0);
  reg [(3'h4):(1'h0)] reg1017 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1016 = (1'h0);
  reg [(3'h6):(1'h0)] reg1014 = (1'h0);
  reg [(3'h5):(1'h0)] reg1013 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1012 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1011 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1010 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1009 = (1'h0);
  reg [(4'h9):(1'h0)] reg1008 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1006 = (1'h0);
  reg [(4'ha):(1'h0)] reg1003 = (1'h0);
  reg signed [(4'he):(1'h0)] reg999 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1004 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1003 = (1'h0);
  reg [(3'h7):(1'h0)] reg1000 = (1'h0);
  reg [(4'hf):(1'h0)] forvar999 = (1'h0);
  reg [(4'hf):(1'h0)] forvar996 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg995 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg994 = (1'h0);
  reg signed [(4'he):(1'h0)] reg993 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar991 = (1'h0);
  reg [(4'he):(1'h0)] forvar990 = (1'h0);
  reg [(4'he):(1'h0)] reg989 = (1'h0);
  reg [(4'hb):(1'h0)] forvar988 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar986 = (1'h0);
  reg [(2'h2):(1'h0)] reg985 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg982 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg980 = (1'h0);
  reg [(4'ha):(1'h0)] forvar979 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg623 = (1'h0);
  reg [(4'hc):(1'h0)] reg622 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg621 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg620 = (1'h0);
  reg [(5'h10):(1'h0)] reg569 = (1'h0);
  reg [(4'hd):(1'h0)] reg617 = (1'h0);
  reg [(4'hd):(1'h0)] reg615 = (1'h0);
  reg [(2'h2):(1'h0)] reg614 = (1'h0);
  reg [(3'h6):(1'h0)] reg613 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar611 = (1'h0);
  reg [(3'h7):(1'h0)] reg610 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar609 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg607 = (1'h0);
  reg [(4'hb):(1'h0)] reg606 = (1'h0);
  reg [(4'hd):(1'h0)] reg605 = (1'h0);
  reg [(4'hd):(1'h0)] reg604 = (1'h0);
  reg [(4'h9):(1'h0)] reg603 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar602 = (1'h0);
  reg [(4'ha):(1'h0)] reg601 = (1'h0);
  reg [(4'hd):(1'h0)] reg599 = (1'h0);
  reg [(4'h9):(1'h0)] reg597 = (1'h0);
  reg [(5'h10):(1'h0)] reg596 = (1'h0);
  reg [(5'h10):(1'h0)] forvar595 = (1'h0);
  reg [(4'h9):(1'h0)] reg594 = (1'h0);
  reg [(2'h2):(1'h0)] forvar593 = (1'h0);
  reg [(4'hb):(1'h0)] forvar592 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg591 = (1'h0);
  reg [(4'h8):(1'h0)] reg589 = (1'h0);
  reg [(4'h8):(1'h0)] forvar588 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg587 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg584 = (1'h0);
  reg [(4'he):(1'h0)] forvar583 = (1'h0);
  reg [(2'h2):(1'h0)] reg578 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg574 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg581 = (1'h0);
  reg [(4'hc):(1'h0)] reg580 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar578 = (1'h0);
  reg [(5'h10):(1'h0)] forvar577 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg576 = (1'h0);
  reg [(2'h3):(1'h0)] forvar575 = (1'h0);
  reg [(5'h10):(1'h0)] forvar574 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg573 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg572 = (1'h0);
  reg [(4'ha):(1'h0)] reg570 = (1'h0);
  reg [(4'h9):(1'h0)] forvar569 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar568 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg567 = (1'h0);
  reg [(3'h4):(1'h0)] reg566 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg565 = (1'h0);
  reg signed [(4'he):(1'h0)] reg564 = (1'h0);
  reg [(4'h8):(1'h0)] reg562 = (1'h0);
  reg [(4'hf):(1'h0)] reg554 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar551 = (1'h0);
  reg [(4'hc):(1'h0)] forvar550 = (1'h0);
  reg [(4'hf):(1'h0)] reg552 = (1'h0);
  reg [(4'ha):(1'h0)] reg560 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg559 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar558 = (1'h0);
  reg [(4'h9):(1'h0)] reg557 = (1'h0);
  reg [(3'h6):(1'h0)] reg556 = (1'h0);
  reg [(3'h6):(1'h0)] reg555 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar554 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar553 = (1'h0);
  reg [(4'hd):(1'h0)] forvar552 = (1'h0);
  assign y = {wire977,
                 wire650,
                 wire647,
                 wire549,
                 reg1121,
                 reg1109,
                 reg1085,
                 reg1100,
                 reg1087,
                 reg1083,
                 reg1062,
                 reg1047,
                 reg1035,
                 reg1034,
                 reg1028,
                 reg1027,
                 reg1024,
                 reg1002,
                 reg1001,
                 reg998,
                 reg997,
                 reg981,
                 reg550,
                 reg558,
                 reg563,
                 reg577,
                 reg586,
                 reg616,
                 reg618,
                 reg1131,
                 reg1130,
                 reg1120,
                 reg1119,
                 reg1118,
                 reg1116,
                 reg1107,
                 reg1104,
                 reg1102,
                 reg1096,
                 reg1080,
                 reg1098,
                 forvar1081,
                 forvar1063,
                 forvar1059,
                 reg1058,
                 reg1064,
                 forvar1062,
                 reg1055,
                 reg1051,
                 forvar1044,
                 reg1043,
                 reg1039,
                 forvar1033,
                 reg1031,
                 reg1023,
                 reg1021,
                 reg1017,
                 reg1013,
                 reg1012,
                 reg1010,
                 forvar1003,
                 forvar999,
                 forvar991,
                 forvar988,
                 forvar979,
                 reg622,
                 reg617,
                 reg614,
                 reg613,
                 forvar611,
                 forvar602,
                 reg601,
                 reg597,
                 reg594,
                 forvar593,
                 reg591,
                 reg589,
                 reg587,
                 reg578,
                 reg574,
                 reg580,
                 forvar575,
                 forvar574,
                 forvar569,
                 forvar568,
                 reg554,
                 reg557,
                 forvar554,
                 forvar553,
                 (1'h0)};
  assign wire549 = (^$signed($signed($unsigned(wire547))));
  always
    @(posedge clk) begin
      if ((^$unsigned((wire549 ? wire548 : $signed(wire545)))))
        begin
          reg550 <= $unsigned(((wire545 >>> (wire545 ?
              wire549 : wire546)) <<< (wire546 != "nfc")));
          reg551 <= $unsigned(((~wire548[(4'hd):(3'h6)]) ?
              (&$signed(wire549)) : "HmYoDKkTF5bgy0"));
          for (forvar552 = (1'h0); (forvar552 < (2'h2)); forvar552 = (forvar552 + (1'h1)))
            begin
              for (forvar553 = (1'h0); (forvar553 < (1'h1)); forvar553 = (forvar553 + (1'h1)))
                begin
                  for (forvar554 = (1'h0); (forvar554 < (2'h2)); forvar554 = (forvar554 + (1'h1)))
                    begin
                      reg555 = wire547[(3'h4):(2'h2)];
                      reg556 = $signed(reg555);
                    end
                  reg557 = forvar552[(3'h6):(2'h2)];
                  for (forvar558 = (1'h0); (forvar558 < (1'h1)); forvar558 = (forvar558 + (1'h1)))
                    begin
                      reg559 = {wire545[(1'h0):(1'h0)]};
                    end
                end
            end
          reg560 = $unsigned(((reg557 ?
                  $unsigned(wire545) : (wire548 - forvar552)) ?
              $signed((forvar558 <<< reg559)) : $signed($unsigned(reg555))));
        end
      else
        begin
          if (reg560)
            begin
              reg552 = wire548[(4'ha):(4'h8)];
            end
          else
            begin
              for (forvar550 = (1'h0); (forvar550 < (2'h3)); forvar550 = (forvar550 + (1'h1)))
                begin
                  for (forvar551 = (1'h0); (forvar551 < (2'h3)); forvar551 = (forvar551 + (1'h1)))
                    begin
                      reg553 <= "drsZltknxzshX";
                      reg554 = $signed({$unsigned($signed(forvar558))});
                      reg555 = "k";
                      reg558 <= $unsigned($unsigned($unsigned({forvar553})));
                    end
                  reg559 = ($unsigned({"1rntqoK4x5Be7"}) + wire548);
                  if ((~"Uc"))
                    begin
                      reg561 <= ($signed($signed(reg553[(4'hc):(4'hb)])) | "qMozTe");
                      reg562 = ((~^$unsigned($unsigned((8'h9d)))) ?
                          $signed((~^reg555)) : $unsigned($signed((forvar552 || reg561))));
                      reg563 <= $unsigned((&$signed($signed(forvar552))));
                      reg564 = {"LGLXYPunBRrecC"};
                    end
                  else
                    begin
                      reg561 <= (wire548 ?
                          $signed((&reg562[(4'h8):(2'h2)])) : (reg563[(2'h2):(1'h0)] >>> forvar551[(2'h3):(2'h3)]));
                    end
                end
              reg565 = reg563[(4'h8):(2'h3)];
            end
          reg566 = (&($unsigned((^wire547)) ?
              ("" ? $unsigned(forvar553) : forvar553[(1'h1):(1'h0)]) : reg557));
          reg567 = ($unsigned(($signed(wire545) ?
              $signed(wire548) : wire549)) & {"hpog2tLCH"});
        end
      if ($unsigned($unsigned((^~wire547))))
        begin
          for (forvar568 = (1'h0); (forvar568 < (2'h3)); forvar568 = (forvar568 + (1'h1)))
            begin
              for (forvar569 = (1'h0); (forvar569 < (2'h2)); forvar569 = (forvar569 + (1'h1)))
                begin
                  if (reg555)
                    begin
                      reg570 = (({$unsigned(reg566)} >> (8'ha8)) ?
                          {"W"} : $signed(forvar569));
                    end
                  else
                    begin
                      reg571 <= {$signed((reg567[(1'h1):(1'h1)] ?
                              $signed(reg565) : (reg559 ? wire547 : wire549)))};
                      reg572 = ((~&("EE5RS7s9yag4" <= $signed(reg552))) ?
                          reg566[(3'h4):(2'h2)] : forvar554[(3'h6):(3'h6)]);
                    end
                  reg573 = $signed(($signed($unsigned(reg552)) & reg559[(1'h0):(1'h0)]));
                end
            end
          if ($unsigned($unsigned({reg564[(4'ha):(1'h1)]})))
            begin
              for (forvar574 = (1'h0); (forvar574 < (2'h2)); forvar574 = (forvar574 + (1'h1)))
                begin
                  for (forvar575 = (1'h0); (forvar575 < (2'h3)); forvar575 = (forvar575 + (1'h1)))
                    begin
                      reg576 = "c9FFadhhsis";
                    end
                end
              for (forvar577 = (1'h0); (forvar577 < (2'h3)); forvar577 = (forvar577 + (1'h1)))
                begin
                  for (forvar578 = (1'h0); (forvar578 < (1'h0)); forvar578 = (forvar578 + (1'h1)))
                    begin
                      reg579 <= reg551[(2'h3):(1'h0)];
                      reg580 = (reg565[(3'h6):(1'h1)] ^~ "YtpON9gzUwk");
                    end
                end
              reg581 = {"xYWg8XvpEA"};
            end
          else
            begin
              if ($signed(reg552[(4'hb):(4'h8)]))
                begin
                  reg574 = (forvar558[(2'h3):(2'h3)] != (forvar578[(1'h0):(1'h0)] ?
                      ($unsigned(reg570) == reg563) : ("USHdH" ?
                          "gsqYx6m0Z2p7d" : (^~reg564))));
                  for (forvar575 = (1'h0); (forvar575 < (1'h0)); forvar575 = (forvar575 + (1'h1)))
                    begin
                      reg577 <= (-reg573[(4'hb):(2'h3)]);
                      reg578 = $unsigned(($unsigned((wire547 && (8'hb8))) ?
                          $unsigned((8'ha3)) : (^$signed((8'ha0)))));
                      reg580 = {$unsigned((8'hae))};
                      reg582 <= reg550[(3'h7):(1'h0)];
                    end
                  for (forvar583 = (1'h0); (forvar583 < (1'h1)); forvar583 = (forvar583 + (1'h1)))
                    begin
                      reg584 = ({$signed(forvar568)} ?
                          forvar553[(2'h2):(2'h2)] : reg553);
                      reg585 <= ((8'ha3) ?
                          "2kvRABL0H3Wt5d" : reg571[(3'h4):(2'h2)]);
                      reg586 <= (-{"ToQh87"});
                      reg587 = forvar577;
                    end
                  for (forvar588 = (1'h0); (forvar588 < (1'h0)); forvar588 = (forvar588 + (1'h1)))
                    begin
                      reg589 = (~|((reg552[(4'hd):(4'hc)] ?
                              $signed(reg577) : {forvar553}) ?
                          $unsigned(reg552[(2'h2):(1'h0)]) : ($unsigned(reg567) | reg551)));
                      reg590 <= $signed((!reg589[(3'h5):(2'h3)]));
                    end
                end
              else
                begin
                  for (forvar574 = (1'h0); (forvar574 < (1'h1)); forvar574 = (forvar574 + (1'h1)))
                    begin
                      reg575 <= "yztfmZi";
                      reg576 = ($unsigned(reg572) < (reg573 ?
                          (|$signed(reg564)) : $unsigned(reg585[(3'h4):(1'h0)])));
                    end
                  if (reg566)
                    begin
                      reg577 <= ($unsigned((^~{reg590})) ?
                          (^{"xDULSSlDQXoA"}) : (($unsigned(reg561) ^~ $unsigned((8'hb9))) >>> (^reg555)));
                      reg578 = $unsigned((8'hba));
                      reg580 = (~reg559[(2'h2):(1'h0)]);
                      reg582 <= $unsigned($unsigned({(reg582 ?
                              (8'ha4) : reg562)}));
                    end
                  else
                    begin
                      reg578 = reg553;
                      reg580 = (~(forvar553 ? reg555 : {(|forvar558)}));
                    end
                  if (reg553)
                    begin
                      reg583 <= wire549;
                    end
                  else
                    begin
                      reg584 = ($signed($signed({reg587})) >= {($signed((8'h9f)) ?
                              (reg577 ? reg562 : reg589) : (+(8'hb5)))});
                    end
                  reg587 = $signed(wire545[(3'h7):(3'h4)]);
                end
              reg591 = $unsigned((~^(|reg567[(4'hf):(4'he)])));
              for (forvar592 = (1'h0); (forvar592 < (1'h0)); forvar592 = (forvar592 + (1'h1)))
                begin
                  for (forvar593 = (1'h0); (forvar593 < (2'h3)); forvar593 = (forvar593 + (1'h1)))
                    begin
                      reg594 = ({$signed((~|reg558))} >= (&($signed((8'hab)) ^ (reg555 >>> reg577))));
                    end
                end
              for (forvar595 = (1'h0); (forvar595 < (2'h2)); forvar595 = (forvar595 + (1'h1)))
                begin
                  reg596 = (!reg582[(2'h2):(1'h0)]);
                  if ("Tx0rN7cw9yzap")
                    begin
                      reg597 = (forvar588[(2'h3):(1'h1)] ?
                          $signed(($unsigned(reg577) ~^ "zIYo1Mgk903xbR")) : (-(~^reg584[(2'h2):(1'h1)])));
                      reg598 <= reg579[(2'h3):(1'h1)];
                      reg599 = reg560[(3'h6):(2'h2)];
                      reg600 <= reg577;
                    end
                  else
                    begin
                      reg597 = (((8'hb9) ? {(~|reg566)} : reg598) ?
                          $unsigned($signed((reg561 ?
                              (8'ha8) : (8'hab)))) : {reg577[(4'hb):(4'h9)]});
                      reg599 = $signed(reg554[(2'h3):(1'h0)]);
                      reg600 <= (wire545 ?
                          forvar577 : {$signed($unsigned(forvar551))});
                      reg601 = (+("IfDc9" ?
                          $unsigned($signed(forvar583)) : "b3K7"));
                    end
                  for (forvar602 = (1'h0); (forvar602 < (1'h0)); forvar602 = (forvar602 + (1'h1)))
                    begin
                      reg603 = $unsigned(reg582);
                      reg604 = ("pSDMTr" && $signed((reg579 <<< "yDhi2Mh")));
                      reg605 = {$unsigned(reg558)};
                    end
                  if ((~^reg575))
                    begin
                      reg606 = ($signed($unsigned((reg585 ?
                          forvar593 : reg563))) != $signed((-(reg586 ?
                          reg586 : (8'ha8)))));
                    end
                  else
                    begin
                      reg606 = {$unsigned(reg583)};
                      reg607 = (~&$unsigned(forvar553[(1'h1):(1'h0)]));
                      reg608 <= forvar568;
                    end
                end
            end
          for (forvar609 = (1'h0); (forvar609 < (2'h3)); forvar609 = (forvar609 + (1'h1)))
            begin
              reg610 = "CJWIDvnb7nk8";
              if ($signed((^~(reg606 * forvar578[(2'h3):(2'h3)]))))
                begin
                  for (forvar611 = (1'h0); (forvar611 < (1'h1)); forvar611 = (forvar611 + (1'h1)))
                    begin
                      reg612 <= (reg590[(2'h2):(2'h2)] ? reg583 : wire545);
                      reg613 = $unsigned(reg604);
                      reg614 = $signed($signed(reg596[(1'h0):(1'h0)]));
                    end
                  if ((^(8'hb7)))
                    begin
                      reg615 = ((~&(8'haf)) ?
                          (($unsigned(forvar550) >> (forvar602 ?
                                  (8'ha6) : reg584)) ?
                              (!(reg581 | reg605)) : reg590) : reg579);
                      reg616 <= {"lsxyNu"};
                      reg617 = $signed(("b" > reg558));
                    end
                  else
                    begin
                      reg615 = $unsigned(forvar609[(4'he):(4'hc)]);
                      reg617 = $unsigned(reg575);
                      reg618 <= $unsigned($unsigned(("Fl9Qzbf0OBE" ?
                          forvar611 : $signed(reg561))));
                    end
                end
              else
                begin
                  for (forvar611 = (1'h0); (forvar611 < (1'h0)); forvar611 = (forvar611 + (1'h1)))
                    begin
                      reg613 = ($unsigned("9XqJqz") - reg558[(3'h4):(2'h3)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar568 = (1'h0); (forvar568 < (1'h0)); forvar568 = (forvar568 + (1'h1)))
            begin
              reg569 = ($signed($unsigned((reg580 ? reg590 : reg596))) ?
                  reg599[(1'h1):(1'h0)] : reg582);
            end
        end
    end
  assign wire619 = wire546[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg620 = (!"bRRn7N1qrGkG");
      reg621 = reg612[(2'h2):(1'h1)];
      reg622 = reg620[(1'h1):(1'h1)];
      reg623 = (reg571 ?
          ({(!reg586)} ?
              {reg575[(4'hb):(4'hb)]} : reg579) : ((reg608 < (&reg551)) ?
              {((8'ha2) == reg571)} : ((reg585 ? reg585 : reg586) ?
                  "uX" : $signed(reg553))));
    end
  module624 #() modinst646 (.wire626(reg583), .wire628(wire549), .clk(clk), .wire625(reg590), .y(wire645), .wire627(wire548), .wire629(reg550));
  assign wire647 = ((+("d" <<< reg579)) - $unsigned(((reg590 ?
                       (8'hb8) : reg550) >= reg583)));
  assign wire648 = ((~|(~^((8'ha2) ? reg558 : reg571))) >= $unsigned(((8'ha1) ?
                       $unsigned(reg608) : (wire546 << (8'ha7)))));
  assign wire649 = reg612[(3'h4):(1'h0)];
  assign wire650 = wire547[(3'h5):(3'h5)];
  module651 #() modinst978 (.clk(clk), .wire653(wire545), .wire652(reg612), .wire654(wire648), .y(wire977), .wire655(reg585));
  always
    @(posedge clk) begin
      for (forvar979 = (1'h0); (forvar979 < (2'h2)); forvar979 = (forvar979 + (1'h1)))
        begin
          if ($signed(wire546[(1'h0):(1'h0)]))
            begin
              if (($signed((wire649[(2'h2):(1'h1)] ?
                      (reg585 ? wire645 : reg618) : wire647)) ?
                  "Xk5" : $signed(((reg551 ?
                      forvar979 : wire546) << {reg598}))))
                begin
                  if ((reg550 ?
                      (((8'hab) ?
                          wire546[(3'h4):(2'h3)] : (wire549 & wire648)) ^ wire650[(1'h0):(1'h0)]) : {reg577}))
                    begin
                      reg980 = ($unsigned({{wire645}}) >> reg551);
                      reg981 <= $signed({(~^reg600[(1'h1):(1'h1)])});
                    end
                  else
                    begin
                      reg980 = $unsigned($unsigned($unsigned($unsigned((8'hae)))));
                      reg982 = reg583[(3'h7):(1'h1)];
                      reg983 <= $unsigned($unsigned($signed((!reg598))));
                    end
                end
              else
                begin
                  if (wire649)
                    begin
                      reg981 <= reg583[(4'h8):(2'h3)];
                      reg983 <= $signed((reg582[(1'h0):(1'h0)] * reg579));
                      reg984 <= ({{wire619}} ?
                          (8'hb3) : (wire547[(2'h2):(1'h0)] >= ((reg571 <<< reg590) * (8'hb4))));
                    end
                  else
                    begin
                      reg981 <= wire546;
                      reg982 = {(({(8'ha2)} ?
                              "PCQd" : (8'h9d)) <= (~^(~wire545)))};
                      reg985 = reg984;
                    end
                  for (forvar986 = (1'h0); (forvar986 < (2'h2)); forvar986 = (forvar986 + (1'h1)))
                    begin
                      reg987 <= (^~$unsigned(((reg579 ? reg985 : reg985) ?
                          $signed(reg612) : (reg612 ? (8'hab) : (8'ha3)))));
                    end
                  for (forvar988 = (1'h0); (forvar988 < (1'h0)); forvar988 = (forvar988 + (1'h1)))
                    begin
                      reg989 = reg590;
                    end
                end
              for (forvar990 = (1'h0); (forvar990 < (2'h2)); forvar990 = (forvar990 + (1'h1)))
                begin
                  for (forvar991 = (1'h0); (forvar991 < (2'h3)); forvar991 = (forvar991 + (1'h1)))
                    begin
                      reg992 <= {"7vqB0XxK8pEygCf"};
                      reg993 = reg571[(2'h2):(1'h1)];
                      reg994 = reg987[(3'h4):(1'h0)];
                    end
                  reg995 = (^~reg612[(3'h6):(3'h5)]);
                  for (forvar996 = (1'h0); (forvar996 < (2'h2)); forvar996 = (forvar996 + (1'h1)))
                    begin
                      reg997 <= $signed((~&{reg993[(3'h6):(1'h0)]}));
                    end
                end
              if (($unsigned(($unsigned(reg585) ^ (reg987 >> reg982))) & $signed(($signed(reg598) ?
                  (reg551 <<< reg583) : $unsigned(wire649)))))
                begin
                  reg998 <= reg575;
                  for (forvar999 = (1'h0); (forvar999 < (2'h2)); forvar999 = (forvar999 + (1'h1)))
                    begin
                      reg1000 = ($unsigned(reg995) - $signed("iUv"));
                      reg1001 <= ($signed(wire647) != reg618[(1'h0):(1'h0)]);
                      reg1002 <= ($unsigned($unsigned(wire650)) > ($signed((reg608 >>> reg997)) == (&$signed(reg598))));
                    end
                  for (forvar1003 = (1'h0); (forvar1003 < (1'h1)); forvar1003 = (forvar1003 + (1'h1)))
                    begin
                      reg1004 = $signed(((+$signed(reg582)) ?
                          ((reg980 ?
                              reg571 : wire645) ~^ (reg994 ~^ wire546)) : $signed(wire977)));
                    end
                end
              else
                begin
                  if ("oPx2")
                    begin
                      reg999 = {($unsigned(((8'hb1) > reg997)) <<< ((reg983 ?
                                  reg980 : (8'hb8)) ?
                              $unsigned(wire648) : (wire619 | reg1000)))};
                      reg1000 = (~wire545);
                      reg1003 = reg579;
                      reg1004 = $unsigned(($unsigned($signed(wire977)) ?
                          ("5VqdERlG2UCdfw" ?
                              reg561[(4'ha):(1'h0)] : ((8'ha3) ?
                                  reg997 : (8'ha5))) : (8'haf)));
                    end
                  else
                    begin
                      reg999 = "4ChPqFTmid";
                      reg1001 <= (~^$signed($signed((~&forvar991))));
                      reg1002 <= forvar990;
                      reg1005 <= $unsigned(reg583[(4'hd):(4'hd)]);
                    end
                  for (forvar1006 = (1'h0); (forvar1006 < (2'h2)); forvar1006 = (forvar1006 + (1'h1)))
                    begin
                      reg1007 <= {({{forvar991}} > ((reg993 + wire649) >>> $signed(reg981)))};
                      reg1008 = (8'ha5);
                    end
                  for (forvar1009 = (1'h0); (forvar1009 < (1'h0)); forvar1009 = (forvar1009 + (1'h1)))
                    begin
                      reg1010 = (reg563 || {(forvar986 ?
                              $unsigned(reg1004) : reg987[(3'h6):(3'h4)])});
                    end
                  for (forvar1011 = (1'h0); (forvar1011 < (1'h0)); forvar1011 = (forvar1011 + (1'h1)))
                    begin
                      reg1012 = $signed(($signed("Km2") ?
                          $signed((+(8'had))) : reg550));
                      reg1013 = ((($unsigned((8'h9d)) ?
                          $signed(forvar996) : $signed((8'had))) >>> ($unsigned(reg989) ?
                          (&reg998) : (~|reg1008))) >>> (^(^$unsigned(forvar996))));
                      reg1014 = ({{(reg550 - reg980)}} ?
                          $unsigned(({wire650} + $signed(reg1000))) : reg998[(1'h0):(1'h0)]);
                      reg1015 <= (~&$unsigned(({wire549} ? reg1007 : reg586)));
                    end
                end
            end
          else
            begin
              reg981 <= forvar979;
            end
          for (forvar1016 = (1'h0); (forvar1016 < (2'h2)); forvar1016 = (forvar1016 + (1'h1)))
            begin
              reg1017 = $signed((~&$signed((+reg582))));
              if (((wire546[(1'h0):(1'h0)] ?
                  reg550[(4'ha):(4'h8)] : {$signed(reg577)}) != (8'had)))
                begin
                  for (forvar1018 = (1'h0); (forvar1018 < (1'h1)); forvar1018 = (forvar1018 + (1'h1)))
                    begin
                      reg1019 = reg558[(3'h4):(3'h4)];
                      reg1020 = ((-wire547) && (~(~|(reg583 || reg1008))));
                    end
                  if (($signed(reg1020[(3'h4):(1'h0)]) ?
                      $signed(((reg586 ?
                          reg984 : reg1001) >>> $signed(forvar991))) : $unsigned((8'ha6))))
                    begin
                      reg1021 = $signed({{reg1001}});
                    end
                  else
                    begin
                      reg1021 = ($signed($signed((reg616 ?
                          forvar1011 : reg585))) && $signed(forvar979[(4'h8):(1'h0)]));
                      reg1022 <= {"U0uSVtXLCR"};
                    end
                  reg1023 = ($unsigned(((reg1013 ? forvar996 : reg561) ?
                      {reg992} : $signed((8'ha1)))) <<< wire650[(1'h0):(1'h0)]);
                end
              else
                begin
                  if (reg1004[(4'h8):(2'h2)])
                    begin
                      reg1018 = ($unsigned($signed((reg1013 << reg1007))) + (!(~reg553)));
                      reg1019 = (reg1007[(3'h6):(3'h6)] << reg608);
                      reg1020 = (^($signed(((8'h9f) > wire645)) << ((reg994 >> (8'hac)) || forvar986)));
                    end
                  else
                    begin
                      reg1022 <= $signed((((wire548 ? reg984 : reg980) ?
                              (forvar986 > reg582) : "DBo") ?
                          forvar986[(4'hb):(3'h7)] : wire545[(3'h6):(3'h4)]));
                      reg1024 <= "J5hxo6XhkGr0kAD";
                      reg1025 <= (reg987[(3'h6):(1'h0)] ?
                          reg1005[(3'h7):(2'h2)] : "QcKtn8u");
                    end
                  for (forvar1026 = (1'h0); (forvar1026 < (2'h3)); forvar1026 = (forvar1026 + (1'h1)))
                    begin
                      reg1027 <= (~|"MYPNDP");
                      reg1028 <= ({$unsigned($signed(reg1022))} ~^ reg1024);
                    end
                  reg1029 = reg1007[(4'ha):(1'h0)];
                  if (reg982[(3'h4):(2'h2)])
                    begin
                      reg1030 = forvar986[(3'h5):(1'h1)];
                      reg1031 = $signed(($signed($unsigned(reg995)) ?
                          ((8'hb1) ^~ (forvar1003 ?
                              reg983 : forvar999)) : (reg583 + (~(8'hb6)))));
                      reg1032 = forvar979[(3'h6):(3'h4)];
                    end
                  else
                    begin
                      reg1030 = (|forvar979);
                      reg1031 = ({reg551} ?
                          $unsigned({$unsigned((8'hb7))}) : $unsigned($signed($unsigned((8'hb4)))));
                      reg1032 = "M";
                    end
                end
              for (forvar1033 = (1'h0); (forvar1033 < (1'h1)); forvar1033 = (forvar1033 + (1'h1)))
                begin
                  if ($signed($signed("w0FBL0gR")))
                    begin
                      reg1034 <= ({wire648[(1'h0):(1'h0)]} * $unsigned(reg1015));
                      reg1035 <= $unsigned(forvar1026);
                      reg1036 = reg583[(4'he):(3'h5)];
                    end
                  else
                    begin
                      reg1034 <= (8'ha0);
                    end
                  for (forvar1037 = (1'h0); (forvar1037 < (2'h2)); forvar1037 = (forvar1037 + (1'h1)))
                    begin
                      reg1038 = {$signed(reg1032[(2'h2):(1'h0)])};
                      reg1039 = ((-(~^(&reg992))) ?
                          "2oLx" : (~^$unsigned(reg981[(3'h4):(1'h1)])));
                      reg1040 <= (wire977 > {$unsigned({reg1007})});
                    end
                  reg1041 <= "Guz3kdinSVH8";
                end
            end
          for (forvar1042 = (1'h0); (forvar1042 < (1'h0)); forvar1042 = (forvar1042 + (1'h1)))
            begin
              reg1043 = (forvar990 ?
                  $signed($signed((forvar979 ? (8'hb5) : wire645))) : reg586);
              for (forvar1044 = (1'h0); (forvar1044 < (2'h3)); forvar1044 = (forvar1044 + (1'h1)))
                begin
                  reg1045 = reg1018[(1'h0):(1'h0)];
                  if (("iAPyBgYzzF" << forvar1042[(1'h0):(1'h0)]))
                    begin
                      reg1046 = (8'h9f);
                      reg1047 <= "Kk";
                      reg1048 = reg1018[(4'h9):(1'h0)];
                    end
                  else
                    begin
                      reg1046 = ((|(((8'hba) ~^ (8'ha3)) ?
                          {forvar1009} : {reg1032})) > $signed(reg1001));
                    end
                  if ($signed("bWYMXbl"))
                    begin
                      reg1049 = (($unsigned((^reg981)) >> "6KTZ5vn") ?
                          reg1017[(1'h0):(1'h0)] : (wire647 ?
                              $signed(reg997) : ({forvar1009} ?
                                  (^reg558) : wire546[(2'h3):(2'h2)])));
                      reg1050 = (~$signed($signed($signed(reg577))));
                      reg1051 = "sRnT2Nbc8";
                      reg1052 <= reg1035[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg1049 = (~&($signed({reg1018}) ?
                          "A" : (+reg987[(3'h5):(3'h4)])));
                      reg1050 = {$unsigned($signed(reg600[(2'h2):(1'h0)]))};
                      reg1052 <= $unsigned((^(~&$unsigned((8'h9e)))));
                    end
                end
              reg1053 <= reg1008;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1054 = (1'h0); (forvar1054 < (1'h0)); forvar1054 = (forvar1054 + (1'h1)))
        begin
          reg1055 = {reg575};
          reg1056 <= $signed(reg558);
        end
      reg1057 <= reg1002[(1'h0):(1'h0)];
      if ($unsigned({$signed((-reg981))}))
        begin
          if ("pJGtsL")
            begin
              for (forvar1058 = (1'h0); (forvar1058 < (2'h2)); forvar1058 = (forvar1058 + (1'h1)))
                begin
                  reg1059 = reg997[(3'h4):(2'h2)];
                end
              reg1060 = (reg582 <<< "udeQduYc");
              for (forvar1061 = (1'h0); (forvar1061 < (1'h1)); forvar1061 = (forvar1061 + (1'h1)))
                begin
                  for (forvar1062 = (1'h0); (forvar1062 < (1'h1)); forvar1062 = (forvar1062 + (1'h1)))
                    begin
                      reg1063 = reg1024[(1'h0):(1'h0)];
                      reg1064 = {(((reg612 ? reg998 : wire648) ?
                                  ((8'hae) >= reg1035) : wire547[(1'h0):(1'h0)]) ?
                              (reg575[(1'h1):(1'h1)] ?
                                  (reg608 ?
                                      forvar1058 : reg1005) : reg608[(4'h9):(1'h0)]) : ($unsigned(reg981) ?
                                  (reg598 ?
                                      wire548 : reg984) : (reg1028 || reg577)))};
                      reg1065 = ((reg582[(1'h0):(1'h0)] ?
                              $unsigned("4") : ({wire549} && "uVck")) ?
                          forvar1062 : reg551[(1'h1):(1'h0)]);
                    end
                  for (forvar1066 = (1'h0); (forvar1066 < (1'h0)); forvar1066 = (forvar1066 + (1'h1)))
                    begin
                      reg1067 = ($signed(reg983) ?
                          $signed(reg1015) : (~|{"dHkFxhaHD"}));
                      reg1068 = ("JURPwYDdc2SCT" ~^ $unsigned($unsigned(wire649)));
                      reg1069 <= ((wire648[(4'h8):(1'h0)] ?
                              ($signed((8'hb7)) + (^reg558)) : (^reg1001[(1'h0):(1'h0)])) ?
                          $unsigned((8'ha4)) : reg1040[(1'h1):(1'h1)]);
                    end
                  reg1070 = reg997;
                end
            end
          else
            begin
              if (({reg553[(2'h2):(1'h1)]} > ((|$unsigned(forvar1061)) != ($signed(reg577) <<< (~^reg1002)))))
                begin
                  reg1058 = (reg608[(2'h2):(1'h0)] ^ (^~$unsigned(((8'had) ?
                      (8'ha3) : forvar1058))));
                  for (forvar1059 = (1'h0); (forvar1059 < (2'h3)); forvar1059 = (forvar1059 + (1'h1)))
                    begin
                      reg1060 = $signed(wire549[(3'h6):(1'h0)]);
                      reg1061 = reg1068[(3'h6):(3'h4)];
                      reg1062 <= $signed((((+reg553) <<< ((8'ha2) < reg616)) ?
                          wire547 : (!$unsigned((8'hb8)))));
                    end
                end
              else
                begin
                  for (forvar1058 = (1'h0); (forvar1058 < (2'h3)); forvar1058 = (forvar1058 + (1'h1)))
                    begin
                      reg1059 = reg590;
                      reg1062 <= $unsigned((~^"NysR"));
                    end
                end
              for (forvar1063 = (1'h0); (forvar1063 < (1'h0)); forvar1063 = (forvar1063 + (1'h1)))
                begin
                  if ((~&((^~{forvar1059}) ^ "E9Ke")))
                    begin
                      reg1064 = ($unsigned((!(reg1063 >>> reg1060))) - $signed($signed(reg586)));
                      reg1065 = (~|"MoKrex5hIAuqR0");
                      reg1066 = $unsigned((wire549 < wire547));
                    end
                  else
                    begin
                      reg1064 = wire649;
                      reg1065 = $signed(($signed($unsigned((8'h9f))) ?
                          (reg1053 - wire649[(3'h7):(3'h7)]) : reg1007[(4'h8):(1'h0)]));
                      reg1066 = {$signed("Uz3oRGWNTu")};
                    end
                  reg1069 <= "0KJ9fDJftgEiB2Y";
                  if (($unsigned(reg1057) << $signed(($signed(reg1056) * reg1068[(1'h1):(1'h1)]))))
                    begin
                      reg1071 <= $signed((~&"IDzTNXHUm4qJ0yI"));
                      reg1072 <= reg553[(4'h8):(1'h1)];
                    end
                  else
                    begin
                      reg1070 = {$signed((reg1067[(4'h8):(3'h7)] ?
                              $unsigned(reg1069) : {reg1052}))};
                    end
                  for (forvar1073 = (1'h0); (forvar1073 < (2'h2)); forvar1073 = (forvar1073 + (1'h1)))
                    begin
                      reg1074 = "4ED";
                    end
                end
            end
          for (forvar1075 = (1'h0); (forvar1075 < (1'h0)); forvar1075 = (forvar1075 + (1'h1)))
            begin
              if ((&reg561))
                begin
                  reg1076 = (((&(reg1067 ?
                          reg983 : reg1041)) <= ((reg558 >> reg575) & $signed((8'ha1)))) ?
                      reg992 : (reg1056 >>> reg1069));
                end
              else
                begin
                  reg1076 = reg583;
                end
            end
          reg1077 <= reg1027;
          for (forvar1078 = (1'h0); (forvar1078 < (1'h1)); forvar1078 = (forvar1078 + (1'h1)))
            begin
              reg1079 <= {wire548};
              for (forvar1080 = (1'h0); (forvar1080 < (2'h3)); forvar1080 = (forvar1080 + (1'h1)))
                begin
                  for (forvar1081 = (1'h0); (forvar1081 < (1'h1)); forvar1081 = (forvar1081 + (1'h1)))
                    begin
                      reg1082 <= "wLcGASaurwcX";
                      reg1083 <= ((8'hba) ? reg575 : wire549[(4'h8):(3'h4)]);
                      reg1084 = (((-reg1015) ?
                          $unsigned("C88q") : reg1041[(4'hf):(4'hc)]) <= $signed({reg1079}));
                    end
                  for (forvar1085 = (1'h0); (forvar1085 < (1'h1)); forvar1085 = (forvar1085 + (1'h1)))
                    begin
                      reg1086 <= "853MfJ9Q";
                      reg1087 <= (wire649[(2'h2):(1'h1)] != (reg600 && $signed(reg1002[(1'h0):(1'h0)])));
                      reg1088 <= (($signed((wire548 <= wire549)) ?
                              "Blz" : ((8'hac) ? reg1053 : $signed(reg1015))) ?
                          $signed(reg577[(4'ha):(3'h6)]) : reg1059[(3'h5):(3'h5)]);
                      reg1089 = "uv";
                    end
                  if ((wire545 >>> "q"))
                    begin
                      reg1090 = reg1005;
                      reg1091 = $unsigned($signed("pd64qZEq"));
                      reg1092 = (reg1089 + "25o851ZQP");
                      reg1093 = ($unsigned((~forvar1063[(4'h8):(4'h8)])) - (-wire650));
                    end
                  else
                    begin
                      reg1090 = wire977[(3'h4):(3'h4)];
                      reg1094 <= reg1066[(1'h1):(1'h0)];
                    end
                end
              for (forvar1095 = (1'h0); (forvar1095 < (2'h2)); forvar1095 = (forvar1095 + (1'h1)))
                begin
                  for (forvar1096 = (1'h0); (forvar1096 < (1'h1)); forvar1096 = (forvar1096 + (1'h1)))
                    begin
                      reg1097 <= reg1092;
                      reg1098 = {($unsigned("wOx7bBp7") << $unsigned((8'ha6)))};
                      reg1099 <= $unsigned((reg550 << reg1061));
                      reg1100 <= reg983[(3'h5):(3'h5)];
                    end
                end
            end
        end
      else
        begin
          reg1058 = (|({reg1077} ~^ (+$signed(wire619))));
          for (forvar1059 = (1'h0); (forvar1059 < (1'h0)); forvar1059 = (forvar1059 + (1'h1)))
            begin
              reg1060 = (~(|$signed(reg571)));
              for (forvar1061 = (1'h0); (forvar1061 < (2'h3)); forvar1061 = (forvar1061 + (1'h1)))
                begin
                  if ($signed($unsigned("1h")))
                    begin
                      reg1063 = (~&reg1060[(4'h9):(3'h4)]);
                    end
                  else
                    begin
                      reg1062 <= $signed($unsigned({{reg1090}}));
                      reg1069 <= "";
                    end
                end
              if ($unsigned(reg984[(3'h5):(2'h3)]))
                begin
                  reg1070 = (+(~{reg616[(2'h2):(2'h2)]}));
                  reg1073 = (8'hb3);
                end
              else
                begin
                  reg1071 <= reg558;
                  for (forvar1072 = (1'h0); (forvar1072 < (2'h3)); forvar1072 = (forvar1072 + (1'h1)))
                    begin
                      reg1073 = reg1083[(1'h1):(1'h0)];
                      reg1074 = ({$unsigned("OvMh")} ?
                          ($signed((wire977 ? (8'hb8) : reg1074)) ?
                              $unsigned(reg1053) : "LN") : (-({forvar1095} >>> ((8'haf) ^~ forvar1073))));
                      reg1075 <= $signed((~(reg1067 ?
                          (^reg550) : $unsigned(reg586))));
                    end
                end
            end
          for (forvar1076 = (1'h0); (forvar1076 < (2'h2)); forvar1076 = (forvar1076 + (1'h1)))
            begin
              for (forvar1077 = (1'h0); (forvar1077 < (2'h2)); forvar1077 = (forvar1077 + (1'h1)))
                begin
                  for (forvar1078 = (1'h0); (forvar1078 < (1'h1)); forvar1078 = (forvar1078 + (1'h1)))
                    begin
                      reg1080 = reg1056[(3'h4):(2'h3)];
                      reg1081 = wire547;
                      reg1084 = ({(~&$unsigned(wire549))} ?
                          reg571[(2'h2):(1'h0)] : ($signed($unsigned(forvar1081)) <<< (+(forvar1075 ^ reg1035))));
                      reg1085 <= reg1005[(4'h8):(4'h8)];
                    end
                  reg1086 <= (~|forvar1085);
                  reg1089 = $signed(((|$signed(forvar1059)) * forvar1077));
                  reg1090 = forvar1081[(4'h9):(3'h7)];
                end
              for (forvar1091 = (1'h0); (forvar1091 < (1'h1)); forvar1091 = (forvar1091 + (1'h1)))
                begin
                  reg1094 <= wire648[(4'hc):(4'hb)];
                end
            end
          if ($unsigned(reg1075))
            begin
              for (forvar1095 = (1'h0); (forvar1095 < (1'h1)); forvar1095 = (forvar1095 + (1'h1)))
                begin
                  if (reg1022)
                    begin
                      reg1096 = $signed({reg1002});
                      reg1097 <= $unsigned((reg551[(2'h3):(1'h0)] ?
                          (~|((8'hb1) || reg551)) : $signed($signed((8'ha7)))));
                    end
                  else
                    begin
                      reg1097 <= reg1073;
                      reg1099 <= {forvar1063[(4'hd):(4'ha)]};
                      reg1101 = reg1047[(2'h3):(2'h2)];
                    end
                  reg1102 = (reg585[(4'ha):(4'h8)] ?
                      forvar1095[(2'h3):(2'h3)] : ({reg1034[(3'h6):(3'h4)]} ?
                          reg612 : $unsigned($unsigned(reg1100))));
                end
              for (forvar1103 = (1'h0); (forvar1103 < (2'h2)); forvar1103 = (forvar1103 + (1'h1)))
                begin
                  if ({(^{reg1088})})
                    begin
                      reg1104 = "UNfmKRO66dxnv";
                    end
                  else
                    begin
                      reg1105 <= (8'ha3);
                    end
                  for (forvar1106 = (1'h0); (forvar1106 < (2'h3)); forvar1106 = (forvar1106 + (1'h1)))
                    begin
                      reg1107 = {(~((!reg1063) ?
                              reg1077[(3'h6):(3'h5)] : (~&reg1015)))};
                      reg1108 = (+"oieDNeuJmyW");
                    end
                  for (forvar1109 = (1'h0); (forvar1109 < (2'h3)); forvar1109 = (forvar1109 + (1'h1)))
                    begin
                      reg1110 <= "fpqRfrD";
                    end
                end
              if (reg583[(4'hd):(4'h8)])
                begin
                  reg1111 = wire546;
                  for (forvar1112 = (1'h0); (forvar1112 < (1'h1)); forvar1112 = (forvar1112 + (1'h1)))
                    begin
                      reg1113 <= "dUA8xElmDI";
                      reg1114 <= $signed((wire649 ?
                          (~(8'h9f)) : "iZuB7VwJ5hk"));
                    end
                  reg1115 <= wire548[(4'hb):(1'h1)];
                end
              else
                begin
                  for (forvar1111 = (1'h0); (forvar1111 < (2'h2)); forvar1111 = (forvar1111 + (1'h1)))
                    begin
                      reg1112 = (~$unsigned(reg1007[(4'ha):(3'h6)]));
                    end
                  reg1116 = (~^reg984[(1'h1):(1'h1)]);
                  for (forvar1117 = (1'h0); (forvar1117 < (2'h2)); forvar1117 = (forvar1117 + (1'h1)))
                    begin
                      reg1118 = (wire647[(1'h1):(1'h1)] <= (("39T1RUkAs" ?
                              reg1065[(2'h3):(1'h1)] : (&reg582)) ?
                          reg1052 : (8'hb3)));
                      reg1119 = $unsigned($signed((+{forvar1081})));
                      reg1120 = reg1104;
                    end
                  for (forvar1121 = (1'h0); (forvar1121 < (2'h3)); forvar1121 = (forvar1121 + (1'h1)))
                    begin
                      reg1122 = $signed(reg1091[(3'h5):(2'h2)]);
                      reg1123 = (|"cw4JsC6Yg");
                      reg1124 = (8'hb0);
                      reg1125 = (~wire549);
                    end
                end
              for (forvar1126 = (1'h0); (forvar1126 < (2'h3)); forvar1126 = (forvar1126 + (1'h1)))
                begin
                  for (forvar1127 = (1'h0); (forvar1127 < (2'h3)); forvar1127 = (forvar1127 + (1'h1)))
                    begin
                      reg1128 = $signed($signed($unsigned(reg1027)));
                      reg1129 <= (((~^((8'h9e) || forvar1091)) || reg1113[(3'h4):(1'h0)]) ?
                          forvar1081[(2'h3):(2'h2)] : "AvrtWPZeBbgR");
                      reg1130 = wire547;
                    end
                end
            end
          else
            begin
              for (forvar1095 = (1'h0); (forvar1095 < (2'h3)); forvar1095 = (forvar1095 + (1'h1)))
                begin
                  reg1097 <= ((reg1102 ?
                      ((reg987 ?
                          forvar1126 : reg1114) << reg571[(3'h6):(3'h4)]) : forvar1066) ^ "DDtfStD7WfH");
                  reg1099 <= (reg575[(4'h8):(4'h8)] && (((8'haf) * reg1064[(1'h0):(1'h0)]) ?
                      ((reg1081 ^~ forvar1076) == $signed(reg1001)) : $unsigned((wire650 ?
                          wire548 : reg1080))));
                  for (forvar1100 = (1'h0); (forvar1100 < (1'h1)); forvar1100 = (forvar1100 + (1'h1)))
                    begin
                      reg1103 <= $unsigned((((reg1116 ?
                          reg1125 : reg1087) + reg612[(2'h2):(1'h0)]) * ($signed(reg1102) * {wire547})));
                      reg1105 <= reg1087[(1'h0):(1'h0)];
                    end
                  for (forvar1106 = (1'h0); (forvar1106 < (2'h3)); forvar1106 = (forvar1106 + (1'h1)))
                    begin
                      reg1109 <= reg585[(3'h5):(1'h0)];
                      reg1111 = (8'hae);
                      reg1112 = "";
                      reg1113 <= ((reg579[(2'h2):(1'h0)] > (~(reg550 ?
                          reg992 : (8'h9d)))) ~^ $unsigned(("7VX2b" ?
                          (reg1097 - reg1076) : (reg1073 ~^ reg1077))));
                    end
                end
              reg1116 = reg550;
              for (forvar1117 = (1'h0); (forvar1117 < (2'h3)); forvar1117 = (forvar1117 + (1'h1)))
                begin
                  for (forvar1118 = (1'h0); (forvar1118 < (2'h3)); forvar1118 = (forvar1118 + (1'h1)))
                    begin
                      reg1121 <= ("FlIXkl4" ? (~reg616) : $signed(reg1099));
                    end
                end
            end
        end
      reg1131 = {$signed(reg1098)};
    end
  assign wire1132 = (!($signed((reg586 <<< reg583)) ^~ (~^"XbGP6Slp0GW")));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module365
#(parameter param497 = ({(8'ha6)} ? (&(((8'hb4) >>> (8'hae)) || {(8'hae)})) : {(((8'ha8) ? (8'ha8) : (8'hab)) ? {(8'hb5)} : (~&(8'hb1)))}))
(y, clk, wire369, wire368, wire367, wire366);
  output wire [(32'h5a6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire369;
  input wire signed [(4'he):(1'h0)] wire368;
  input wire [(4'hf):(1'h0)] wire367;
  input wire signed [(3'h4):(1'h0)] wire366;
  wire signed [(4'h8):(1'h0)] wire496;
  wire signed [(3'h7):(1'h0)] wire370;
  reg signed [(5'h10):(1'h0)] reg495 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg446 = (1'h0);
  reg [(3'h4):(1'h0)] reg437 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg436 = (1'h0);
  reg [(4'hd):(1'h0)] reg427 = (1'h0);
  reg [(4'hc):(1'h0)] reg490 = (1'h0);
  reg [(4'hf):(1'h0)] reg487 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg486 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg485 = (1'h0);
  reg [(2'h2):(1'h0)] reg483 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg479 = (1'h0);
  reg [(4'h8):(1'h0)] reg466 = (1'h0);
  reg signed [(4'he):(1'h0)] reg472 = (1'h0);
  reg [(3'h4):(1'h0)] reg470 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg469 = (1'h0);
  reg [(4'he):(1'h0)] reg465 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg464 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg462 = (1'h0);
  reg [(3'h6):(1'h0)] reg459 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg453 = (1'h0);
  reg signed [(4'he):(1'h0)] reg451 = (1'h0);
  reg signed [(4'he):(1'h0)] reg450 = (1'h0);
  reg [(5'h10):(1'h0)] reg449 = (1'h0);
  reg [(5'h10):(1'h0)] reg443 = (1'h0);
  reg [(4'h9):(1'h0)] reg442 = (1'h0);
  reg [(4'hb):(1'h0)] reg440 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg439 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg434 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg429 = (1'h0);
  reg [(2'h3):(1'h0)] reg424 = (1'h0);
  reg [(4'he):(1'h0)] reg423 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg421 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg420 = (1'h0);
  reg [(3'h5):(1'h0)] reg418 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg417 = (1'h0);
  reg [(3'h6):(1'h0)] reg411 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg406 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg403 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg398 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg395 = (1'h0);
  reg [(3'h6):(1'h0)] reg388 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg386 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg383 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg381 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg380 = (1'h0);
  reg [(3'h4):(1'h0)] reg377 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg376 = (1'h0);
  reg [(4'hc):(1'h0)] reg494 = (1'h0);
  reg [(4'hc):(1'h0)] forvar493 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg492 = (1'h0);
  reg [(3'h6):(1'h0)] reg457 = (1'h0);
  reg [(3'h4):(1'h0)] reg455 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar453 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg452 = (1'h0);
  reg signed [(4'he):(1'h0)] reg448 = (1'h0);
  reg [(4'he):(1'h0)] forvar447 = (1'h0);
  reg [(4'hf):(1'h0)] forvar443 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg441 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar438 = (1'h0);
  reg [(4'h8):(1'h0)] reg431 = (1'h0);
  reg [(4'hf):(1'h0)] reg426 = (1'h0);
  reg signed [(4'he):(1'h0)] reg491 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg489 = (1'h0);
  reg [(4'ha):(1'h0)] reg488 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg484 = (1'h0);
  reg [(4'hf):(1'h0)] reg482 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg481 = (1'h0);
  reg [(3'h6):(1'h0)] reg480 = (1'h0);
  reg [(2'h3):(1'h0)] reg478 = (1'h0);
  reg [(4'h9):(1'h0)] forvar477 = (1'h0);
  reg [(4'h8):(1'h0)] reg476 = (1'h0);
  reg [(4'h9):(1'h0)] reg475 = (1'h0);
  reg [(4'hc):(1'h0)] forvar474 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg471 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar462 = (1'h0);
  reg [(4'hb):(1'h0)] reg474 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg473 = (1'h0);
  reg [(3'h6):(1'h0)] forvar471 = (1'h0);
  reg [(4'hc):(1'h0)] reg468 = (1'h0);
  reg [(4'hc):(1'h0)] reg467 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar466 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg463 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg461 = (1'h0);
  reg [(4'hb):(1'h0)] reg460 = (1'h0);
  reg [(3'h4):(1'h0)] reg458 = (1'h0);
  reg [(3'h6):(1'h0)] forvar457 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg456 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar455 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg454 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar452 = (1'h0);
  reg [(4'he):(1'h0)] forvar448 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg447 = (1'h0);
  reg [(3'h6):(1'h0)] forvar446 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar445 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg445 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg444 = (1'h0);
  reg [(3'h6):(1'h0)] forvar441 = (1'h0);
  reg [(2'h2):(1'h0)] reg438 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar437 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar436 = (1'h0);
  reg [(3'h5):(1'h0)] reg435 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg433 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar431 = (1'h0);
  reg [(3'h7):(1'h0)] reg430 = (1'h0);
  reg [(5'h10):(1'h0)] reg428 = (1'h0);
  reg [(4'ha):(1'h0)] forvar427 = (1'h0);
  reg [(2'h2):(1'h0)] forvar426 = (1'h0);
  reg [(4'he):(1'h0)] forvar425 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar413 = (1'h0);
  reg [(4'hf):(1'h0)] reg422 = (1'h0);
  reg [(4'hb):(1'h0)] forvar419 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar416 = (1'h0);
  reg [(4'hc):(1'h0)] reg415 = (1'h0);
  reg [(4'hb):(1'h0)] reg410 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar408 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar405 = (1'h0);
  reg [(4'h9):(1'h0)] reg414 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg413 = (1'h0);
  reg [(4'h8):(1'h0)] reg412 = (1'h0);
  reg [(3'h5):(1'h0)] forvar410 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg409 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg408 = (1'h0);
  reg [(4'hf):(1'h0)] reg407 = (1'h0);
  reg [(3'h4):(1'h0)] reg404 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg402 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg401 = (1'h0);
  reg [(4'he):(1'h0)] reg400 = (1'h0);
  reg [(5'h10):(1'h0)] reg399 = (1'h0);
  reg signed [(4'he):(1'h0)] reg397 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar396 = (1'h0);
  reg [(3'h4):(1'h0)] reg391 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg396 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar395 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg394 = (1'h0);
  reg [(3'h5):(1'h0)] reg393 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg392 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar391 = (1'h0);
  reg [(4'hc):(1'h0)] reg390 = (1'h0);
  reg [(2'h3):(1'h0)] forvar389 = (1'h0);
  reg [(4'he):(1'h0)] forvar387 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg375 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg385 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg384 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg382 = (1'h0);
  reg [(4'he):(1'h0)] reg379 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg378 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar375 = (1'h0);
  reg [(3'h5):(1'h0)] reg374 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar373 = (1'h0);
  reg [(4'hb):(1'h0)] forvar372 = (1'h0);
  reg [(4'h8):(1'h0)] reg371 = (1'h0);
  assign y = {wire496,
                 reg495,
                 reg446,
                 reg437,
                 reg436,
                 reg490,
                 reg483,
                 reg453,
                 reg443,
                 reg440,
                 reg439,
                 reg434,
                 reg421,
                 reg403,
                 reg380,
                 reg377,
                 reg494,
                 reg492,
                 reg455,
                 forvar453,
                 reg448,
                 forvar443,
                 reg491,
                 reg489,
                 reg482,
                 reg481,
                 reg480,
                 reg478,
                 reg475,
                 reg471,
                 forvar462,
                 forvar471,
                 reg461,
                 forvar452,
                 forvar448,
                 forvar441,
                 forvar437,
                 forvar436,
                 reg430,
                 forvar405,
                 reg412,
                 forvar410,
                 reg397,
                 forvar396,
                 forvar395,
                 forvar389,
                 reg385,
                 reg384,
                 reg382,
                 reg378,
                 reg374,
                 forvar372,
                 (1'h0)};
  assign wire370 = {wire368};
  always
    @(posedge clk) begin
      reg371 = "R8dwcAHzY2czR";
      if (reg371[(1'h0):(1'h0)])
        begin
          for (forvar372 = (1'h0); (forvar372 < (2'h3)); forvar372 = (forvar372 + (1'h1)))
            begin
              for (forvar373 = (1'h0); (forvar373 < (2'h3)); forvar373 = (forvar373 + (1'h1)))
                begin
                  reg374 = (&((^~wire368[(4'h9):(1'h1)]) >>> "G4x"));
                  for (forvar375 = (1'h0); (forvar375 < (2'h2)); forvar375 = (forvar375 + (1'h1)))
                    begin
                      reg376 <= wire368[(3'h7):(3'h4)];
                      reg377 <= "8";
                      reg378 = forvar372;
                      reg379 = ({((~&wire370) << forvar375[(2'h3):(2'h2)])} ?
                          $unsigned((!"GTp9MgIdX")) : $signed("p"));
                    end
                  reg380 <= $unsigned("Ydvv");
                  if (((($signed(reg379) ?
                          (&reg377) : (reg376 ? (8'hb9) : wire366)) ?
                      reg371 : $signed("K7HceCRJ4JzD3")) != $unsigned(((wire366 && wire370) ?
                      {reg379} : $signed(reg379)))))
                    begin
                      reg381 <= reg371;
                      reg382 = (^reg381);
                    end
                  else
                    begin
                      reg382 = wire367[(4'he):(4'ha)];
                    end
                end
              reg383 <= ("VYtkz" && "YY");
              reg384 = (($unsigned((+reg378)) ?
                  wire370[(1'h0):(1'h0)] : reg374[(1'h0):(1'h0)]) != (^~$unsigned((wire370 << (8'ha1)))));
            end
          reg385 = forvar375;
        end
      else
        begin
          for (forvar372 = (1'h0); (forvar372 < (1'h0)); forvar372 = (forvar372 + (1'h1)))
            begin
              for (forvar373 = (1'h0); (forvar373 < (1'h0)); forvar373 = (forvar373 + (1'h1)))
                begin
                  if ({$unsigned(forvar375)})
                    begin
                      reg374 = $unsigned(({((8'hb1) >= reg382)} == reg377));
                      reg375 = ($unsigned(($signed(reg383) ?
                              $signed(reg371) : (~^wire368))) ?
                          {(^(reg380 ?
                                  reg379 : reg383))} : (wire370[(1'h0):(1'h0)] ?
                              wire370[(1'h0):(1'h0)] : $unsigned($signed((8'hb2)))));
                    end
                  else
                    begin
                      reg374 = $unsigned($unsigned(""));
                      reg375 = $signed((reg384 * (reg380 ~^ (+reg375))));
                      reg376 <= "SBZ";
                      reg378 = "K";
                    end
                  if (forvar372)
                    begin
                      reg379 = $unsigned((!wire367));
                      reg380 <= $unsigned((8'ha3));
                      reg381 <= (!"NB");
                      reg382 = $unsigned((-((~|forvar373) ?
                          reg371[(4'h8):(1'h0)] : $signed(wire369))));
                    end
                  else
                    begin
                      reg380 <= ($signed({$unsigned(reg376)}) ?
                          $unsigned($unsigned(wire369)) : ($unsigned((8'hb4)) ?
                              ($signed(wire367) ?
                                  $unsigned(reg381) : reg380[(2'h2):(2'h2)]) : (reg377 ^ (reg377 & reg385))));
                      reg381 <= $unsigned($signed(wire367[(4'he):(4'hd)]));
                      reg382 = reg374;
                      reg384 = (|"1apaqgCmRlFZBX");
                    end
                  reg385 = reg375;
                  reg386 <= "Sb";
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar387 = (1'h0); (forvar387 < (2'h3)); forvar387 = (forvar387 + (1'h1)))
        begin
          reg388 <= (reg381 ? "IXGK7fl" : {reg386[(1'h0):(1'h0)]});
          for (forvar389 = (1'h0); (forvar389 < (2'h3)); forvar389 = (forvar389 + (1'h1)))
            begin
              reg390 = $unsigned($signed($unsigned(reg376[(4'hd):(4'hd)])));
              if (((|(^(forvar389 + forvar389))) ?
                  (~|$unsigned(wire366[(1'h0):(1'h0)])) : "f"))
                begin
                  for (forvar391 = (1'h0); (forvar391 < (2'h2)); forvar391 = (forvar391 + (1'h1)))
                    begin
                      reg392 = $unsigned($signed($signed(reg377)));
                      reg393 = ($signed((8'hb9)) <<< (~|(^~(8'hb0))));
                    end
                  reg394 = $signed((+reg388));
                  for (forvar395 = (1'h0); (forvar395 < (1'h1)); forvar395 = (forvar395 + (1'h1)))
                    begin
                      reg396 = ($unsigned(((forvar391 ?
                              reg388 : forvar387) & (8'hab))) ?
                          $unsigned($signed(reg386)) : (8'hb6));
                    end
                end
              else
                begin
                  reg391 = reg388[(1'h1):(1'h0)];
                  reg395 <= $unsigned(((8'hb7) > (|((8'ha0) ?
                      reg383 : forvar391))));
                  for (forvar396 = (1'h0); (forvar396 < (2'h3)); forvar396 = (forvar396 + (1'h1)))
                    begin
                      reg397 = "C83xZkSqeRVlCI";
                      reg398 <= {(+$signed(((8'hb0) ^ reg383)))};
                    end
                  if ("DL08691")
                    begin
                      reg399 = reg392[(1'h0):(1'h0)];
                      reg400 = {({(^(8'hb1))} ?
                              $unsigned($signed(reg399)) : reg394)};
                      reg401 = forvar387;
                      reg402 = wire367;
                    end
                  else
                    begin
                      reg399 = $unsigned(reg397);
                    end
                end
              reg403 <= (~&(~$unsigned(reg396[(1'h1):(1'h0)])));
              reg404 = $unsigned((~^reg402));
            end
          if ("RgTwYk")
            begin
              if (($signed(reg395) ?
                  {$unsigned(wire368)} : ($unsigned("VMp2Je") ?
                      $unsigned("FgPRIJ") : $signed($signed(forvar389)))))
                begin
                  if (($signed((8'hb8)) ?
                      $signed({"QL"}) : (({wire369} ? (!(8'hb3)) : (^~reg391)) ?
                          ($unsigned(reg395) ?
                              (~&reg397) : (wire367 ?
                                  (8'ha1) : wire370)) : {$signed((8'hb6))})))
                    begin
                      reg405 <= reg377[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg405 <= $unsigned("nuoXn5tUxp");
                    end
                  if (reg391[(2'h3):(2'h3)])
                    begin
                      reg406 <= ($unsigned({(wire369 ?
                              wire368 : reg392)}) >= reg398);
                      reg407 = forvar396[(2'h2):(2'h2)];
                      reg408 = $signed("fboF1gJOB");
                      reg409 = reg395[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg407 = ("MnfmbRAukGHXd2z" ?
                          reg388 : (reg391[(1'h0):(1'h0)] ?
                              (reg395[(3'h5):(2'h2)] ?
                                  reg401 : ((8'hb1) ?
                                      forvar389 : reg376)) : (forvar387[(4'he):(4'hb)] ?
                                  $unsigned(reg405) : (~^wire369))));
                      reg408 = reg403;
                      reg409 = (((reg403[(4'hd):(2'h2)] ?
                              (8'hb7) : (reg388 << reg408)) ?
                          (((8'ha4) * (8'ha4)) ?
                              (reg390 ~^ reg377) : $unsigned(reg396)) : (|$unsigned(reg396))) * reg394);
                    end
                  for (forvar410 = (1'h0); (forvar410 < (2'h2)); forvar410 = (forvar410 + (1'h1)))
                    begin
                      reg411 <= {("8w3X" || (~(|reg399)))};
                      reg412 = {($unsigned("r6rRJq") ~^ $signed({(8'hb0)}))};
                      reg413 = reg399;
                    end
                  if ((~|$unsigned({(-forvar389)})))
                    begin
                      reg414 = reg397;
                    end
                  else
                    begin
                      reg414 = $unsigned(($unsigned((reg407 ?
                              reg401 : reg383)) ?
                          (^{(8'ha5)}) : reg390));
                    end
                end
              else
                begin
                  for (forvar405 = (1'h0); (forvar405 < (1'h0)); forvar405 = (forvar405 + (1'h1)))
                    begin
                      reg406 <= $signed({$signed("xXYA4KX")});
                      reg407 = reg396;
                    end
                  for (forvar408 = (1'h0); (forvar408 < (2'h2)); forvar408 = (forvar408 + (1'h1)))
                    begin
                      reg409 = {{((reg413 ?
                                  (8'h9c) : (8'ha1)) << $signed(forvar408))}};
                      reg410 = ((forvar410 ?
                          reg388 : {$unsigned((8'ha1))}) == reg398[(2'h2):(1'h0)]);
                    end
                  reg412 = (8'ha0);
                end
              reg415 = ({reg405} ?
                  (^~(~^reg411[(1'h0):(1'h0)])) : $signed($unsigned(wire366[(1'h0):(1'h0)])));
              for (forvar416 = (1'h0); (forvar416 < (1'h0)); forvar416 = (forvar416 + (1'h1)))
                begin
                  reg417 <= reg414[(4'h8):(4'h8)];
                  reg418 <= (&(($unsigned((8'ha8)) < {reg397}) + (&"Butqu4tAMkLAp")));
                  for (forvar419 = (1'h0); (forvar419 < (1'h1)); forvar419 = (forvar419 + (1'h1)))
                    begin
                      reg420 <= $signed($signed(reg404[(2'h2):(2'h2)]));
                      reg421 <= $signed($unsigned(reg380[(1'h1):(1'h0)]));
                      reg422 = $signed(("CKuV" ?
                          reg420 : ({reg398} ?
                              reg417[(3'h5):(3'h5)] : reg380[(1'h0):(1'h0)])));
                      reg423 <= (+{$signed($signed(forvar391))});
                    end
                end
            end
          else
            begin
              for (forvar405 = (1'h0); (forvar405 < (1'h0)); forvar405 = (forvar405 + (1'h1)))
                begin
                  reg407 = ($unsigned({$unsigned(reg398)}) << reg402);
                  if ($unsigned(((~(reg395 + (8'ha8))) <<< (forvar405[(4'h9):(3'h5)] - (forvar391 - wire369)))))
                    begin
                      reg408 = (&(((reg417 ?
                              forvar396 : (8'hb8)) <<< (~|reg386)) ?
                          $signed($signed(forvar416)) : ((~|(8'ha7)) ?
                              (reg390 == reg402) : (forvar395 ?
                                  (8'hb1) : reg376))));
                    end
                  else
                    begin
                      reg408 = reg393[(3'h5):(2'h2)];
                      reg411 <= reg403[(3'h6):(2'h2)];
                      reg412 = reg421[(2'h3):(2'h3)];
                    end
                end
              for (forvar413 = (1'h0); (forvar413 < (2'h3)); forvar413 = (forvar413 + (1'h1)))
                begin
                  reg414 = reg413[(2'h3):(1'h0)];
                end
              reg415 = $unsigned(reg408[(2'h3):(2'h2)]);
            end
          reg424 <= (reg403[(4'h8):(3'h7)] ?
              reg377 : (reg391[(2'h2):(1'h0)] ?
                  ((reg401 * (8'ha4)) - $unsigned((8'haa))) : forvar389[(2'h3):(1'h1)]));
        end
      if ((8'ha3))
        begin
          for (forvar425 = (1'h0); (forvar425 < (1'h0)); forvar425 = (forvar425 + (1'h1)))
            begin
              for (forvar426 = (1'h0); (forvar426 < (2'h2)); forvar426 = (forvar426 + (1'h1)))
                begin
                  for (forvar427 = (1'h0); (forvar427 < (2'h3)); forvar427 = (forvar427 + (1'h1)))
                    begin
                      reg428 = {$signed($unsigned(reg413[(1'h0):(1'h0)]))};
                      reg429 <= {reg403[(1'h0):(1'h0)]};
                      reg430 = ((!forvar410[(2'h2):(1'h1)]) >= $signed($unsigned(reg412)));
                    end
                  for (forvar431 = (1'h0); (forvar431 < (2'h2)); forvar431 = (forvar431 + (1'h1)))
                    begin
                      reg432 = (8'hb6);
                      reg433 = ((reg407[(3'h5):(3'h4)] > (-$unsigned(reg430))) ?
                          ($signed({reg383}) + (reg410[(4'h9):(3'h6)] + $signed(reg409))) : reg391);
                      reg434 <= $signed("2v4YO19xguzVg");
                      reg435 = forvar419;
                    end
                end
              for (forvar436 = (1'h0); (forvar436 < (2'h3)); forvar436 = (forvar436 + (1'h1)))
                begin
                  for (forvar437 = (1'h0); (forvar437 < (2'h3)); forvar437 = (forvar437 + (1'h1)))
                    begin
                      reg438 = (reg420 && (&reg423));
                      reg439 <= "a";
                      reg440 <= reg380;
                    end
                  for (forvar441 = (1'h0); (forvar441 < (1'h0)); forvar441 = (forvar441 + (1'h1)))
                    begin
                      reg442 <= "9M";
                    end
                  reg443 <= (8'ha2);
                end
            end
          reg444 = "Ag";
          if ({(^~("fngqUZ5H" << (~&reg405)))})
            begin
              reg445 = (forvar413 ? (|reg417[(3'h7):(3'h7)]) : {reg411});
            end
          else
            begin
              for (forvar445 = (1'h0); (forvar445 < (2'h3)); forvar445 = (forvar445 + (1'h1)))
                begin
                  for (forvar446 = (1'h0); (forvar446 < (1'h0)); forvar446 = (forvar446 + (1'h1)))
                    begin
                      reg447 = (reg413 >>> (~|$signed($unsigned(reg414))));
                    end
                  for (forvar448 = (1'h0); (forvar448 < (2'h2)); forvar448 = (forvar448 + (1'h1)))
                    begin
                      reg449 <= {{($unsigned((8'hb0)) <<< (~forvar431))}};
                      reg450 <= ({reg432[(1'h0):(1'h0)]} >= {$unsigned(((8'ha1) + reg381))});
                      reg451 <= (~^(+(8'hb6)));
                    end
                  for (forvar452 = (1'h0); (forvar452 < (1'h0)); forvar452 = (forvar452 + (1'h1)))
                    begin
                      reg453 <= (reg432 ?
                          {reg383} : {(forvar410 | (~&reg421))});
                      reg454 = ($unsigned("htHFI4") ?
                          $signed(reg447[(2'h2):(1'h0)]) : reg443[(4'hd):(4'h9)]);
                    end
                end
              for (forvar455 = (1'h0); (forvar455 < (1'h1)); forvar455 = (forvar455 + (1'h1)))
                begin
                  reg456 = ("zTxLmIa" == (reg445 ?
                      ($unsigned(forvar437) ?
                          {reg392} : $unsigned((8'h9c))) : "stHqN5tV2"));
                  for (forvar457 = (1'h0); (forvar457 < (1'h0)); forvar457 = (forvar457 + (1'h1)))
                    begin
                      reg458 = (reg404[(1'h1):(1'h1)] ?
                          (|((^~reg435) & $signed(reg429))) : $unsigned(reg412[(1'h0):(1'h0)]));
                      reg459 <= reg414;
                      reg460 = reg408;
                      reg461 = $signed(reg438);
                    end
                end
              if (forvar441)
                begin
                  if (("El1P" ?
                      forvar391[(3'h4):(1'h1)] : reg377[(2'h2):(1'h0)]))
                    begin
                      reg462 <= {$signed("")};
                      reg463 = $unsigned({reg440});
                      reg464 <= $signed((-$unsigned("954m")));
                      reg465 <= (((-"rSgiIXS") ?
                          (((8'ha5) >>> reg459) >= ((8'hb2) ?
                              forvar416 : wire367)) : reg429) <= ($signed(reg410[(4'hb):(1'h0)]) ?
                          "HnxO5IzOeVIm0gn" : (~reg388)));
                    end
                  else
                    begin
                      reg462 <= $unsigned(forvar436);
                    end
                  for (forvar466 = (1'h0); (forvar466 < (2'h3)); forvar466 = (forvar466 + (1'h1)))
                    begin
                      reg467 = (~|($unsigned((8'ha3)) >> {$signed(forvar441)}));
                      reg468 = reg444[(4'h9):(2'h2)];
                      reg469 <= (~($unsigned(forvar446[(2'h3):(1'h0)]) ?
                          (reg451 ~^ reg386[(3'h4):(3'h4)]) : (reg383 > ((8'hb4) ?
                              (8'had) : forvar408))));
                    end
                  reg470 <= $signed((($unsigned(reg412) + (forvar391 ?
                      reg462 : reg442)) >> ((reg468 ?
                      (8'ha4) : reg434) < forvar452[(1'h1):(1'h0)])));
                  for (forvar471 = (1'h0); (forvar471 < (1'h0)); forvar471 = (forvar471 + (1'h1)))
                    begin
                      reg472 <= "";
                      reg473 = (("3JptszPaQa5Wa" > $signed((forvar410 ?
                              reg442 : reg467))) ?
                          (8'h9c) : $signed({{(8'ha8)}}));
                      reg474 = reg434[(2'h2):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar462 = (1'h0); (forvar462 < (1'h0)); forvar462 = (forvar462 + (1'h1)))
                    begin
                      reg464 <= {$signed(forvar466[(1'h1):(1'h1)])};
                      reg465 <= $signed((~&{{forvar445}}));
                    end
                  if ((!reg454[(5'h10):(3'h5)]))
                    begin
                      reg466 <= (reg434 <<< ((-"sBXk4VwBLClhFpC") > forvar408));
                      reg469 <= ($unsigned(($unsigned(reg465) ?
                              (+forvar441) : (|reg449))) ?
                          (reg463 ^~ reg402) : (~|((8'ha6) ?
                              (reg409 ?
                                  forvar436 : forvar457) : reg376[(3'h7):(1'h0)])));
                      reg471 = {reg472[(1'h0):(1'h0)]};
                      reg473 = reg381[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg467 = forvar419[(2'h2):(1'h0)];
                      reg468 = (((8'ha8) ?
                              $signed($unsigned(forvar419)) : (+$signed((8'h9c)))) ?
                          reg376 : $unsigned(((reg459 << reg466) * (8'h9c))));
                    end
                  for (forvar474 = (1'h0); (forvar474 < (2'h2)); forvar474 = (forvar474 + (1'h1)))
                    begin
                      reg475 = $signed((~forvar431[(4'hd):(4'hb)]));
                      reg476 = (^$unsigned(((^~(8'ha6)) ?
                          reg392 : reg394[(4'h9):(4'h8)])));
                    end
                  for (forvar477 = (1'h0); (forvar477 < (1'h1)); forvar477 = (forvar477 + (1'h1)))
                    begin
                      reg478 = "z0q297vMF";
                      reg479 <= ($signed(($unsigned(reg430) + (reg451 != reg470))) ?
                          $unsigned($unsigned($unsigned(reg458))) : $unsigned($signed({forvar445})));
                      reg480 = $unsigned((!{{(8'haa)}}));
                    end
                end
              if ($signed($signed(((forvar455 << reg418) ?
                  (&forvar396) : forvar446[(1'h0):(1'h0)]))))
                begin
                  reg481 = $unsigned(((|(forvar389 ~^ (8'ha6))) & $unsigned({wire370})));
                  reg482 = ($signed("uotuBWoouB1W") ?
                      forvar445[(3'h5):(2'h2)] : ($signed(((8'hac) ?
                          reg428 : reg453)) >= "rub3sTZDQwgeEp"));
                end
              else
                begin
                  if ((~^($signed(((8'hab) == reg475)) & $signed((reg391 ?
                      reg433 : reg481)))))
                    begin
                      reg483 <= $unsigned({(forvar455[(3'h7):(3'h5)] ?
                              (^~(8'h9f)) : (^~reg411))});
                      reg484 = {((reg458 <<< (~|reg377)) * ((reg376 ?
                              forvar391 : reg402) || (reg445 ?
                              forvar471 : forvar455)))};
                    end
                  else
                    begin
                      reg483 <= reg481;
                      reg485 <= "ny";
                    end
                  if (((+reg429[(3'h5):(3'h4)]) + $unsigned("g")))
                    begin
                      reg486 <= ($signed(reg410[(4'hb):(3'h4)]) ?
                          reg458[(3'h4):(2'h3)] : $signed(((forvar391 ^ forvar446) & $signed(forvar466))));
                      reg487 <= ($signed(($unsigned(reg393) >> (-reg399))) ?
                          ($unsigned(forvar431) <= {(reg391 ?
                                  (8'hb8) : (8'hac))}) : $unsigned($unsigned({reg381})));
                      reg488 = reg450;
                      reg489 = "";
                    end
                  else
                    begin
                      reg488 = $signed({$unsigned((&reg478))});
                      reg490 <= reg443;
                      reg491 = forvar437[(2'h3):(2'h3)];
                    end
                end
            end
        end
      else
        begin
          for (forvar425 = (1'h0); (forvar425 < (1'h0)); forvar425 = (forvar425 + (1'h1)))
            begin
              if ({"3lnwYTmkGa4"})
                begin
                  reg426 = $signed(reg435[(1'h1):(1'h1)]);
                end
              else
                begin
                  reg427 <= $unsigned($unsigned({$signed(reg439)}));
                  if ((((8'h9d) ?
                          ($signed(reg430) ?
                              $signed(reg484) : $signed(reg403)) : wire367) ?
                      (forvar413 ?
                          ((forvar477 ?
                              (8'hb1) : reg426) ^ reg406) : reg408) : $unsigned((|(reg490 >> (8'hb1))))))
                    begin
                      reg428 = $unsigned($signed(reg426[(1'h0):(1'h0)]));
                      reg429 <= $unsigned($unsigned({{forvar436}}));
                      reg430 = $unsigned($unsigned((forvar437[(1'h0):(1'h0)] ^~ reg463)));
                      reg431 = reg398;
                    end
                  else
                    begin
                      reg429 <= (($unsigned((8'ha9)) ?
                          forvar466[(1'h0):(1'h0)] : forvar413) >> ((^~forvar387) ?
                          (+forvar425[(1'h1):(1'h1)]) : ($signed(reg381) << ((8'had) ?
                              (8'had) : reg415))));
                      reg430 = reg399[(4'hb):(4'ha)];
                      reg434 <= {(~&(~|((8'hb4) & reg397)))};
                      reg436 <= (8'ha7);
                    end
                end
              reg437 <= (reg485 >>> reg485);
              if (reg478)
                begin
                  for (forvar438 = (1'h0); (forvar438 < (1'h0)); forvar438 = (forvar438 + (1'h1)))
                    begin
                      reg441 = $signed((($signed(forvar395) || reg413[(1'h0):(1'h0)]) ?
                          reg476[(4'h8):(3'h5)] : "P5GxpNbWt"));
                    end
                end
              else
                begin
                  for (forvar438 = (1'h0); (forvar438 < (1'h0)); forvar438 = (forvar438 + (1'h1)))
                    begin
                      reg441 = reg480;
                    end
                  reg442 <= ($unsigned(((reg451 ?
                          reg462 : reg443) | {reg439})) ?
                      $unsigned(((forvar455 - forvar445) ?
                          reg410[(3'h4):(2'h2)] : (wire367 + reg376))) : (|$unsigned({reg460})));
                end
              if (((~^((-forvar452) < $unsigned((8'had)))) > reg417))
                begin
                  for (forvar443 = (1'h0); (forvar443 < (2'h3)); forvar443 = (forvar443 + (1'h1)))
                    begin
                      reg444 = reg377;
                      reg445 = {reg430[(3'h6):(3'h5)]};
                    end
                  reg446 <= "wS";
                end
              else
                begin
                  reg444 = ((reg438 && (-reg454[(4'hf):(4'hf)])) ?
                      reg461 : (^reg478[(2'h3):(1'h0)]));
                  reg446 <= forvar446;
                  for (forvar447 = (1'h0); (forvar447 < (2'h2)); forvar447 = (forvar447 + (1'h1)))
                    begin
                      reg448 = {(^reg437)};
                      reg452 = reg399;
                    end
                  for (forvar453 = (1'h0); (forvar453 < (2'h3)); forvar453 = (forvar453 + (1'h1)))
                    begin
                      reg454 = $signed($unsigned($signed((~|forvar408))));
                      reg455 = "JWbwEQ";
                      reg456 = (8'ha0);
                    end
                end
            end
          reg457 = (|$signed($unsigned((~^reg386))));
        end
      reg492 = $unsigned(($unsigned("") - (-(reg458 ? (8'haa) : reg394))));
    end
  always
    @(posedge clk) begin
      for (forvar493 = (1'h0); (forvar493 < (2'h2)); forvar493 = (forvar493 + (1'h1)))
        begin
          reg494 = {reg437};
          reg495 <= (|(&$signed((reg388 ? reg464 : reg395))));
        end
    end
  assign wire496 = (~&$signed((reg424 ?
                       $signed((8'hb9)) : reg490[(1'h1):(1'h0)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module651
#(parameter param976 = ((!(~|((8'ha5) & (8'hb4)))) ? ((|((8'ha7) ? (8'h9d) : (8'hb4))) ? {{(8'h9f)}} : (((8'hb4) ? (8'ha0) : (8'hb9)) ? (!(8'h9d)) : (&(8'hb2)))) : ((^~{(8'h9c)}) > ({(8'hb1)} * ((8'hb1) ? (8'haf) : (8'hac))))))
(y, clk, wire655, wire654, wire653, wire652);
  output wire [(32'hd4d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire655;
  input wire [(4'h8):(1'h0)] wire654;
  input wire signed [(4'h8):(1'h0)] wire653;
  input wire [(4'h9):(1'h0)] wire652;
  wire signed [(4'h8):(1'h0)] wire737;
  wire signed [(3'h5):(1'h0)] wire656;
  reg [(4'h9):(1'h0)] reg971 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg968 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg966 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg961 = (1'h0);
  reg [(3'h4):(1'h0)] reg957 = (1'h0);
  reg [(3'h7):(1'h0)] reg958 = (1'h0);
  reg [(5'h10):(1'h0)] reg951 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg947 = (1'h0);
  reg [(3'h5):(1'h0)] reg945 = (1'h0);
  reg [(4'ha):(1'h0)] reg943 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg942 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg937 = (1'h0);
  reg [(4'h8):(1'h0)] reg934 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg933 = (1'h0);
  reg [(4'h9):(1'h0)] reg932 = (1'h0);
  reg [(4'hd):(1'h0)] reg929 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg924 = (1'h0);
  reg [(3'h4):(1'h0)] reg913 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg923 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg921 = (1'h0);
  reg [(4'hc):(1'h0)] reg915 = (1'h0);
  reg [(4'hf):(1'h0)] reg914 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg907 = (1'h0);
  reg [(3'h4):(1'h0)] reg895 = (1'h0);
  reg [(4'hb):(1'h0)] reg902 = (1'h0);
  reg [(3'h4):(1'h0)] reg898 = (1'h0);
  reg [(4'ha):(1'h0)] reg892 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg890 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg882 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg888 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg884 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg883 = (1'h0);
  reg [(5'h10):(1'h0)] reg879 = (1'h0);
  reg [(4'hf):(1'h0)] reg877 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg876 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg875 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg873 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg871 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg867 = (1'h0);
  reg [(4'he):(1'h0)] reg865 = (1'h0);
  reg [(4'hd):(1'h0)] reg864 = (1'h0);
  reg [(4'h8):(1'h0)] reg863 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg859 = (1'h0);
  reg [(4'ha):(1'h0)] reg858 = (1'h0);
  reg [(4'hf):(1'h0)] reg845 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg842 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg811 = (1'h0);
  reg [(2'h3):(1'h0)] reg813 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg855 = (1'h0);
  reg [(3'h7):(1'h0)] reg854 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg851 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg850 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg847 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg839 = (1'h0);
  reg [(3'h5):(1'h0)] reg836 = (1'h0);
  reg [(2'h2):(1'h0)] reg835 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg830 = (1'h0);
  reg signed [(4'he):(1'h0)] reg825 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg823 = (1'h0);
  reg [(2'h2):(1'h0)] reg821 = (1'h0);
  reg [(3'h5):(1'h0)] reg820 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg818 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg814 = (1'h0);
  reg [(3'h4):(1'h0)] reg809 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg808 = (1'h0);
  reg [(3'h5):(1'h0)] reg804 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg794 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg793 = (1'h0);
  reg [(4'he):(1'h0)] reg792 = (1'h0);
  reg [(4'hd):(1'h0)] reg786 = (1'h0);
  reg [(3'h4):(1'h0)] reg784 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg781 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg775 = (1'h0);
  reg [(4'ha):(1'h0)] reg773 = (1'h0);
  reg [(4'he):(1'h0)] reg758 = (1'h0);
  reg [(3'h4):(1'h0)] reg757 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg755 = (1'h0);
  reg [(4'h9):(1'h0)] reg754 = (1'h0);
  reg [(3'h4):(1'h0)] reg752 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg750 = (1'h0);
  reg [(4'h8):(1'h0)] reg747 = (1'h0);
  reg [(5'h10):(1'h0)] reg746 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg744 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg740 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg736 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg733 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg732 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg729 = (1'h0);
  reg [(5'h10):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg722 = (1'h0);
  reg [(2'h3):(1'h0)] reg721 = (1'h0);
  reg [(4'h9):(1'h0)] reg718 = (1'h0);
  reg [(4'hc):(1'h0)] reg711 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg709 = (1'h0);
  reg [(3'h7):(1'h0)] reg708 = (1'h0);
  reg [(5'h10):(1'h0)] reg706 = (1'h0);
  reg [(4'h8):(1'h0)] reg704 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg701 = (1'h0);
  reg [(3'h4):(1'h0)] reg699 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg696 = (1'h0);
  reg [(3'h6):(1'h0)] reg686 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg685 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg694 = (1'h0);
  reg [(4'h8):(1'h0)] reg691 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg689 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg684 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg683 = (1'h0);
  reg [(3'h4):(1'h0)] reg681 = (1'h0);
  reg [(3'h7):(1'h0)] reg667 = (1'h0);
  reg [(4'hd):(1'h0)] reg662 = (1'h0);
  reg signed [(4'he):(1'h0)] reg658 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg678 = (1'h0);
  reg [(3'h5):(1'h0)] reg677 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg673 = (1'h0);
  reg [(4'hc):(1'h0)] reg669 = (1'h0);
  reg [(3'h6):(1'h0)] reg668 = (1'h0);
  reg [(3'h6):(1'h0)] reg665 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg664 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg661 = (1'h0);
  reg [(3'h7):(1'h0)] reg975 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg974 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg973 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar972 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar970 = (1'h0);
  reg [(4'hb):(1'h0)] reg969 = (1'h0);
  reg [(5'h10):(1'h0)] reg967 = (1'h0);
  reg [(4'hc):(1'h0)] reg965 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg964 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar963 = (1'h0);
  reg [(4'hb):(1'h0)] reg962 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg960 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg959 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar957 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg956 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg955 = (1'h0);
  reg [(4'hb):(1'h0)] reg954 = (1'h0);
  reg [(4'h9):(1'h0)] reg953 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg952 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg950 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg949 = (1'h0);
  reg [(3'h6):(1'h0)] reg948 = (1'h0);
  reg [(4'hb):(1'h0)] reg935 = (1'h0);
  reg [(3'h7):(1'h0)] forvar933 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg941 = (1'h0);
  reg [(4'h9):(1'h0)] reg946 = (1'h0);
  reg [(4'he):(1'h0)] reg944 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar941 = (1'h0);
  reg signed [(4'he):(1'h0)] reg940 = (1'h0);
  reg [(2'h3):(1'h0)] reg939 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg938 = (1'h0);
  reg [(3'h5):(1'h0)] reg936 = (1'h0);
  reg [(4'hb):(1'h0)] forvar935 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg931 = (1'h0);
  reg [(4'hc):(1'h0)] forvar930 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg928 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg927 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar926 = (1'h0);
  reg [(4'he):(1'h0)] forvar925 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg916 = (1'h0);
  reg [(4'hf):(1'h0)] reg922 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg920 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg919 = (1'h0);
  reg [(2'h3):(1'h0)] reg918 = (1'h0);
  reg [(4'he):(1'h0)] reg917 = (1'h0);
  reg [(4'ha):(1'h0)] forvar916 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar913 = (1'h0);
  reg [(4'ha):(1'h0)] reg912 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg911 = (1'h0);
  reg [(4'hb):(1'h0)] reg910 = (1'h0);
  reg [(4'hf):(1'h0)] forvar909 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar908 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg906 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg905 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg904 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar903 = (1'h0);
  reg [(3'h4):(1'h0)] reg901 = (1'h0);
  reg [(2'h2):(1'h0)] forvar900 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg899 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg897 = (1'h0);
  reg [(4'hc):(1'h0)] reg896 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar895 = (1'h0);
  reg [(4'hb):(1'h0)] reg894 = (1'h0);
  reg [(3'h4):(1'h0)] reg893 = (1'h0);
  reg [(4'he):(1'h0)] forvar891 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg885 = (1'h0);
  reg [(4'hd):(1'h0)] forvar876 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg891 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar890 = (1'h0);
  reg [(3'h7):(1'h0)] reg889 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg887 = (1'h0);
  reg [(5'h10):(1'h0)] forvar886 = (1'h0);
  reg [(5'h10):(1'h0)] forvar885 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar882 = (1'h0);
  reg [(3'h6):(1'h0)] reg881 = (1'h0);
  reg [(4'h8):(1'h0)] reg880 = (1'h0);
  reg [(4'ha):(1'h0)] reg878 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg872 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg874 = (1'h0);
  reg [(4'h9):(1'h0)] forvar872 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg870 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg869 = (1'h0);
  reg [(4'h9):(1'h0)] reg868 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg866 = (1'h0);
  reg [(4'hd):(1'h0)] reg862 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg861 = (1'h0);
  reg [(4'h9):(1'h0)] forvar860 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg857 = (1'h0);
  reg [(4'hc):(1'h0)] reg856 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar853 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar851 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar841 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar835 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar825 = (1'h0);
  reg signed [(4'he):(1'h0)] reg824 = (1'h0);
  reg [(2'h3):(1'h0)] forvar815 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg853 = (1'h0);
  reg [(4'hf):(1'h0)] reg852 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg849 = (1'h0);
  reg [(4'ha):(1'h0)] reg848 = (1'h0);
  reg [(3'h5):(1'h0)] reg846 = (1'h0);
  reg [(4'hd):(1'h0)] forvar845 = (1'h0);
  reg [(4'he):(1'h0)] reg844 = (1'h0);
  reg [(3'h5):(1'h0)] reg843 = (1'h0);
  reg [(4'h8):(1'h0)] forvar842 = (1'h0);
  reg [(3'h6):(1'h0)] reg837 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg833 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg841 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg840 = (1'h0);
  reg [(4'hd):(1'h0)] reg838 = (1'h0);
  reg [(4'ha):(1'h0)] forvar837 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg834 = (1'h0);
  reg [(3'h6):(1'h0)] forvar833 = (1'h0);
  reg [(3'h7):(1'h0)] reg819 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg832 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg831 = (1'h0);
  reg [(3'h4):(1'h0)] reg829 = (1'h0);
  reg [(4'hd):(1'h0)] reg828 = (1'h0);
  reg [(5'h10):(1'h0)] reg827 = (1'h0);
  reg [(5'h10):(1'h0)] reg826 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar824 = (1'h0);
  reg [(4'ha):(1'h0)] reg822 = (1'h0);
  reg [(4'hd):(1'h0)] forvar819 = (1'h0);
  reg [(3'h4):(1'h0)] reg817 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg816 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg815 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar813 = (1'h0);
  reg [(4'hb):(1'h0)] reg812 = (1'h0);
  reg [(4'he):(1'h0)] forvar811 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar810 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg807 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg806 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar805 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg803 = (1'h0);
  reg [(4'hc):(1'h0)] forvar802 = (1'h0);
  reg [(4'hc):(1'h0)] reg801 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar800 = (1'h0);
  reg [(4'hc):(1'h0)] forvar799 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg798 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg797 = (1'h0);
  reg [(4'hd):(1'h0)] reg796 = (1'h0);
  reg [(3'h6):(1'h0)] forvar795 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar791 = (1'h0);
  reg [(4'h9):(1'h0)] reg790 = (1'h0);
  reg [(3'h5):(1'h0)] reg789 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg788 = (1'h0);
  reg [(2'h2):(1'h0)] reg787 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar785 = (1'h0);
  reg [(3'h4):(1'h0)] forvar783 = (1'h0);
  reg [(3'h4):(1'h0)] reg782 = (1'h0);
  reg [(3'h7):(1'h0)] forvar780 = (1'h0);
  reg [(2'h2):(1'h0)] reg779 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar778 = (1'h0);
  reg [(3'h6):(1'h0)] reg777 = (1'h0);
  reg signed [(4'he):(1'h0)] reg776 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg774 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg772 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg771 = (1'h0);
  reg [(4'hd):(1'h0)] reg770 = (1'h0);
  reg [(4'hc):(1'h0)] reg769 = (1'h0);
  reg [(4'hc):(1'h0)] reg768 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar767 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar766 = (1'h0);
  reg signed [(4'he):(1'h0)] reg761 = (1'h0);
  reg [(4'he):(1'h0)] forvar760 = (1'h0);
  reg [(3'h7):(1'h0)] forvar743 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar742 = (1'h0);
  reg [(4'hc):(1'h0)] reg765 = (1'h0);
  reg [(2'h2):(1'h0)] reg764 = (1'h0);
  reg [(4'hb):(1'h0)] reg763 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg762 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar761 = (1'h0);
  reg [(2'h3):(1'h0)] reg760 = (1'h0);
  reg [(3'h7):(1'h0)] reg759 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar755 = (1'h0);
  reg [(3'h5):(1'h0)] forvar753 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg756 = (1'h0);
  reg [(4'hc):(1'h0)] reg753 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg751 = (1'h0);
  reg [(4'hb):(1'h0)] reg749 = (1'h0);
  reg [(4'hd):(1'h0)] forvar748 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg745 = (1'h0);
  reg [(3'h7):(1'h0)] reg743 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg742 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg741 = (1'h0);
  reg [(4'h9):(1'h0)] forvar739 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar738 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg714 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg705 = (1'h0);
  reg [(3'h7):(1'h0)] forvar699 = (1'h0);
  reg [(3'h6):(1'h0)] forvar698 = (1'h0);
  reg [(5'h10):(1'h0)] forvar696 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg735 = (1'h0);
  reg [(4'hb):(1'h0)] reg734 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar731 = (1'h0);
  reg [(5'h10):(1'h0)] forvar730 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg728 = (1'h0);
  reg [(3'h6):(1'h0)] reg727 = (1'h0);
  reg [(3'h6):(1'h0)] forvar726 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar725 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar723 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar720 = (1'h0);
  reg [(3'h7):(1'h0)] forvar719 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg717 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar716 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg715 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar714 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg713 = (1'h0);
  reg [(4'h9):(1'h0)] reg712 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg710 = (1'h0);
  reg [(3'h7):(1'h0)] reg707 = (1'h0);
  reg [(3'h7):(1'h0)] forvar705 = (1'h0);
  reg [(2'h2):(1'h0)] reg703 = (1'h0);
  reg [(4'hd):(1'h0)] reg702 = (1'h0);
  reg [(5'h10):(1'h0)] reg700 = (1'h0);
  reg [(4'he):(1'h0)] forvar697 = (1'h0);
  reg [(4'he):(1'h0)] forvar700 = (1'h0);
  reg [(3'h4):(1'h0)] reg698 = (1'h0);
  reg [(3'h5):(1'h0)] reg697 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg695 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg693 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar692 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg690 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg688 = (1'h0);
  reg [(2'h3):(1'h0)] reg687 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar686 = (1'h0);
  reg [(4'ha):(1'h0)] forvar685 = (1'h0);
  reg [(4'ha):(1'h0)] reg682 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar665 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar664 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg657 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar668 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg663 = (1'h0);
  reg [(4'h9):(1'h0)] forvar661 = (1'h0);
  reg [(4'h8):(1'h0)] reg680 = (1'h0);
  reg [(3'h4):(1'h0)] reg679 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar671 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg676 = (1'h0);
  reg [(4'hd):(1'h0)] reg675 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg674 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg672 = (1'h0);
  reg [(4'he):(1'h0)] reg671 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg670 = (1'h0);
  reg [(4'hc):(1'h0)] forvar667 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg666 = (1'h0);
  reg [(2'h3):(1'h0)] forvar663 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar662 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg660 = (1'h0);
  reg [(3'h5):(1'h0)] reg659 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar658 = (1'h0);
  reg [(5'h10):(1'h0)] forvar657 = (1'h0);
  assign y = {wire656,
                 reg968,
                 reg951,
                 reg945,
                 reg943,
                 reg934,
                 reg933,
                 reg923,
                 reg921,
                 reg907,
                 reg895,
                 reg898,
                 reg888,
                 reg877,
                 reg876,
                 reg867,
                 reg863,
                 reg858,
                 reg845,
                 reg813,
                 reg847,
                 reg835,
                 reg809,
                 reg808,
                 reg804,
                 reg792,
                 reg786,
                 reg773,
                 reg758,
                 reg754,
                 reg746,
                 reg733,
                 reg732,
                 reg729,
                 reg721,
                 reg711,
                 reg709,
                 reg701,
                 reg699,
                 reg696,
                 reg685,
                 reg689,
                 reg677,
                 reg668,
                 reg665,
                 forvar970,
                 reg962,
                 reg960,
                 reg959,
                 reg950,
                 reg940,
                 reg938,
                 forvar930,
                 reg928,
                 forvar925,
                 reg920,
                 reg918,
                 forvar913,
                 reg910,
                 forvar909,
                 reg905,
                 reg901,
                 reg899,
                 reg896,
                 reg894,
                 reg885,
                 forvar876,
                 reg891,
                 forvar890,
                 reg887,
                 reg881,
                 reg872,
                 reg874,
                 reg869,
                 forvar851,
                 forvar835,
                 reg853,
                 forvar845,
                 reg841,
                 reg827,
                 reg826,
                 forvar819,
                 reg816,
                 reg812,
                 forvar811,
                 forvar810,
                 reg806,
                 reg803,
                 reg801,
                 forvar799,
                 forvar795,
                 reg788,
                 reg787,
                 reg779,
                 reg777,
                 reg776,
                 reg771,
                 reg768,
                 forvar766,
                 forvar760,
                 forvar743,
                 forvar742,
                 reg765,
                 reg762,
                 forvar761,
                 reg760,
                 reg749,
                 reg742,
                 forvar739,
                 reg735,
                 reg727,
                 forvar726,
                 forvar725,
                 forvar720,
                 reg717,
                 forvar714,
                 reg712,
                 reg707,
                 forvar705,
                 forvar697,
                 forvar700,
                 reg698,
                 reg695,
                 forvar692,
                 reg687,
                 forvar686,
                 forvar665,
                 reg657,
                 reg680,
                 reg672,
                 reg660,
                 reg659,
                 (1'h0)};
  assign wire656 = $unsigned(wire654);
  always
    @(posedge clk) begin
      if ((&$unsigned(wire653[(3'h5):(2'h2)])))
        begin
          for (forvar657 = (1'h0); (forvar657 < (1'h1)); forvar657 = (forvar657 + (1'h1)))
            begin
              for (forvar658 = (1'h0); (forvar658 < (1'h0)); forvar658 = (forvar658 + (1'h1)))
                begin
                  if (forvar658)
                    begin
                      reg659 = {((8'hb3) <= wire656[(2'h3):(1'h0)])};
                      reg660 = ($unsigned(($signed(wire654) < $unsigned(forvar658))) ?
                          (|$unsigned(wire654[(1'h1):(1'h0)])) : ({$unsigned(wire653)} ?
                              (^~(-wire656)) : ({wire655} ?
                                  $unsigned(forvar658) : wire654)));
                      reg661 <= (-reg659[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg659 = $unsigned(reg661);
                    end
                end
            end
          for (forvar662 = (1'h0); (forvar662 < (1'h0)); forvar662 = (forvar662 + (1'h1)))
            begin
              for (forvar663 = (1'h0); (forvar663 < (1'h1)); forvar663 = (forvar663 + (1'h1)))
                begin
                  if ("wszn")
                    begin
                      reg664 <= {((+(~|forvar657)) | {wire654})};
                    end
                  else
                    begin
                      reg664 <= $signed(forvar658);
                    end
                end
              reg665 <= wire654;
              if (wire656[(2'h3):(1'h1)])
                begin
                  reg666 = wire653;
                  for (forvar667 = (1'h0); (forvar667 < (1'h0)); forvar667 = (forvar667 + (1'h1)))
                    begin
                      reg668 <= wire654;
                      reg669 <= $unsigned("");
                      reg670 = (8'ha9);
                      reg671 = reg668;
                    end
                  reg672 = ((^("Gbh8ydfx" < forvar663)) ?
                      wire656 : $signed("Uddr"));
                  if (($signed(forvar663) <<< (~{(!wire654)})))
                    begin
                      reg673 <= reg659[(1'h1):(1'h1)];
                      reg674 = ((wire653[(1'h1):(1'h0)] ?
                              (wire656 << (wire654 ?
                                  wire654 : reg673)) : forvar658[(2'h2):(1'h1)]) ?
                          reg664 : (~reg660));
                    end
                  else
                    begin
                      reg674 = reg668[(3'h4):(1'h0)];
                      reg675 = "xSeZ";
                      reg676 = (reg668[(2'h2):(2'h2)] ?
                          reg672 : $unsigned({forvar667}));
                      reg677 <= ({(-(reg664 >= reg660))} ?
                          (!((~reg671) ?
                              (reg672 ?
                                  forvar663 : (8'h9d)) : $unsigned(reg675))) : {$unsigned($signed(forvar663))});
                    end
                end
              else
                begin
                  reg666 = {reg668};
                  for (forvar667 = (1'h0); (forvar667 < (2'h3)); forvar667 = (forvar667 + (1'h1)))
                    begin
                      reg670 = (!$signed(((^(8'hae)) ?
                          {wire654} : (&forvar667))));
                    end
                  for (forvar671 = (1'h0); (forvar671 < (1'h1)); forvar671 = (forvar671 + (1'h1)))
                    begin
                      reg673 <= $unsigned((-((reg665 << (8'h9e)) ~^ reg666)));
                    end
                end
              reg678 <= $signed($signed($signed({reg676})));
            end
          reg679 = "";
          reg680 = (-($signed({reg668}) >>> "bmZnIYgx"));
        end
      else
        begin
          if (($signed(reg676[(2'h2):(1'h0)]) | ($signed(reg674[(2'h2):(1'h0)]) || reg674[(1'h1):(1'h0)])))
            begin
              if (forvar662)
                begin
                  for (forvar657 = (1'h0); (forvar657 < (2'h3)); forvar657 = (forvar657 + (1'h1)))
                    begin
                      reg658 <= (!$signed($unsigned((-forvar667))));
                      reg659 = (!{$signed({reg679})});
                    end
                  reg660 = wire655;
                  for (forvar661 = (1'h0); (forvar661 < (1'h1)); forvar661 = (forvar661 + (1'h1)))
                    begin
                      reg662 <= (&(reg659[(2'h2):(1'h0)] <<< (reg680 & "Ml")));
                      reg663 = $unsigned($signed(reg665));
                      reg666 = $unsigned(reg669);
                    end
                  reg667 <= {$signed(("VL" <<< (^reg677)))};
                end
              else
                begin
                  for (forvar657 = (1'h0); (forvar657 < (2'h2)); forvar657 = (forvar657 + (1'h1)))
                    begin
                      reg659 = {(^reg663)};
                      reg660 = "Q7ZEqVV";
                    end
                end
              if ("NoTAmLIcu0U")
                begin
                  reg670 = "srED";
                  if ("2zFuemT8o2AnZ")
                    begin
                      reg671 = reg677[(3'h4):(1'h1)];
                      reg673 <= $signed($signed(reg678[(2'h2):(2'h2)]));
                      reg677 <= $signed($unsigned((&(~reg669))));
                      reg679 = ($unsigned(reg677[(1'h0):(1'h0)]) ?
                          "TYeo9g5eL" : (+reg658));
                    end
                  else
                    begin
                      reg671 = reg661[(1'h0):(1'h0)];
                      reg672 = (|reg661[(3'h5):(1'h0)]);
                      reg674 = $unsigned($unsigned(((~^wire655) ?
                          $unsigned(reg670) : $unsigned(reg672))));
                      reg677 <= ((($signed(reg676) & $signed(reg674)) > wire653[(1'h1):(1'h0)]) ^~ $signed((8'h9d)));
                    end
                end
              else
                begin
                  for (forvar668 = (1'h0); (forvar668 < (1'h1)); forvar668 = (forvar668 + (1'h1)))
                    begin
                      reg670 = forvar661[(1'h0):(1'h0)];
                    end
                  for (forvar671 = (1'h0); (forvar671 < (1'h0)); forvar671 = (forvar671 + (1'h1)))
                    begin
                      reg673 <= "4l";
                      reg674 = ((reg665[(3'h4):(3'h4)] | (8'ha9)) * $unsigned(((reg673 ?
                          (8'hb7) : (8'hb9)) & $unsigned(forvar667))));
                      reg677 <= (~($unsigned((reg670 ?
                          wire652 : (8'h9c))) && (reg670[(2'h3):(1'h0)] ?
                          wire656 : (-reg671))));
                      reg679 = $unsigned((((reg677 == reg662) ?
                              {(8'ha2)} : {(8'ha8)}) ?
                          reg670 : $signed($unsigned(reg673))));
                    end
                end
            end
          else
            begin
              if (($unsigned((-(&wire652))) ^~ {$unsigned((forvar667 - reg671))}))
                begin
                  for (forvar657 = (1'h0); (forvar657 < (1'h1)); forvar657 = (forvar657 + (1'h1)))
                    begin
                      reg659 = (({(|reg662)} ?
                              ((|forvar668) ?
                                  reg669[(1'h1):(1'h1)] : $unsigned((8'ha4))) : $unsigned({wire655})) ?
                          (("w41xm7J55Ouxl" | wire656[(2'h3):(2'h3)]) != (&$unsigned(forvar657))) : $unsigned((^~$signed((8'hb6)))));
                      reg661 <= $signed($unsigned(reg672[(2'h2):(2'h2)]));
                    end
                end
              else
                begin
                  reg657 = ("wNLpVCbhQQDkL" >= (~|reg667[(1'h1):(1'h1)]));
                  reg659 = $signed((-{$signed(reg677)}));
                end
              reg663 = $signed(reg666);
              for (forvar664 = (1'h0); (forvar664 < (2'h3)); forvar664 = (forvar664 + (1'h1)))
                begin
                  for (forvar665 = (1'h0); (forvar665 < (1'h0)); forvar665 = (forvar665 + (1'h1)))
                    begin
                      reg666 = (+(+reg664));
                      reg670 = ($unsigned(reg680) ^ reg659);
                      reg671 = forvar668;
                    end
                  if (reg679[(1'h1):(1'h1)])
                    begin
                      reg672 = ("v5QHK57t2c" + ("rVDxWTge5FRo" && (~^"Uti9ihqCzkNrym")));
                      reg673 <= ((+reg661[(3'h6):(2'h2)]) ?
                          $signed(($unsigned(reg674) ?
                              reg665[(1'h1):(1'h1)] : (forvar661 ?
                                  (8'ha4) : reg660))) : $signed($signed("HyEmUheWt")));
                      reg674 = wire654[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg672 = $unsigned("31QC8x");
                      reg674 = (reg669 ?
                          wire654[(3'h4):(3'h4)] : ((reg660 ^ reg675) ?
                              ((~reg666) ?
                                  $unsigned(reg679) : $signed(reg668)) : forvar668));
                      reg675 = ({(reg658[(3'h5):(1'h0)] >> reg662[(4'hd):(4'hc)])} <<< ($unsigned({forvar668}) >> ({(8'h9d)} ?
                          forvar668 : (forvar661 ? (8'ha7) : wire652))));
                    end
                  if ($unsigned(wire655[(4'h8):(3'h7)]))
                    begin
                      reg676 = ("lmzSu" == ($signed($signed(forvar671)) << ((forvar664 ?
                          reg672 : reg658) ~^ (reg669 | reg667))));
                      reg677 <= $signed($signed(reg673[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg676 = $signed(((((8'hb9) & (8'ha2)) ?
                          (~|wire655) : reg665) & (^~{reg672})));
                      reg677 <= $unsigned((((forvar661 ?
                              reg673 : reg670) >= $unsigned(reg673)) ?
                          $unsigned(reg664) : (^~forvar668[(1'h0):(1'h0)])));
                      reg679 = "mTxJVLkCyu";
                    end
                  if ("")
                    begin
                      reg680 = reg671[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg680 = ($signed($signed($unsigned(reg663))) || (8'h9d));
                      reg681 <= "toKPYTZcCQh73O9";
                      reg682 = ({$signed({reg665})} & wire652);
                      reg683 <= ("ewQdEb" ?
                          (reg663 <= $signed(wire652)) : {({reg665} ?
                                  (forvar657 * reg671) : {forvar662})});
                    end
                end
              reg684 <= $unsigned(reg671);
            end
          if ($signed($unsigned((~&$unsigned((8'ha3))))))
            begin
              for (forvar685 = (1'h0); (forvar685 < (1'h1)); forvar685 = (forvar685 + (1'h1)))
                begin
                  for (forvar686 = (1'h0); (forvar686 < (2'h2)); forvar686 = (forvar686 + (1'h1)))
                    begin
                      reg687 = $unsigned((($unsigned(reg667) >= ((8'ha7) ?
                              forvar658 : reg660)) ?
                          (((8'ha9) <<< forvar668) ~^ (!wire656)) : {(reg658 ?
                                  reg678 : reg677)}));
                      reg688 = reg676[(2'h3):(1'h1)];
                      reg689 <= "V0pynf7AOYED9V";
                    end
                  reg690 = $signed(reg687[(2'h3):(1'h1)]);
                  reg691 <= $unsigned($unsigned((reg657[(2'h2):(1'h1)] >>> $signed(forvar664))));
                  for (forvar692 = (1'h0); (forvar692 < (2'h2)); forvar692 = (forvar692 + (1'h1)))
                    begin
                      reg693 = (($signed((forvar685 ? reg667 : wire656)) ?
                          reg659[(1'h1):(1'h1)] : {(forvar657 ?
                                  reg689 : reg672)}) * $unsigned(wire655[(3'h4):(2'h2)]));
                      reg694 <= $signed((8'hb8));
                    end
                end
              reg695 = forvar662;
            end
          else
            begin
              if ("U9TJVkhOu")
                begin
                  reg685 <= $unsigned("DY");
                  reg686 <= {{reg694}};
                end
              else
                begin
                  reg687 = (wire652 ? reg689 : "VmBpV");
                end
            end
        end
      if ($unsigned($unsigned($signed((reg676 ? reg671 : reg679)))))
        begin
          if (((~|$unsigned(((8'ha2) ? reg684 : reg680))) ?
              reg669[(4'ha):(4'ha)] : wire653))
            begin
              reg696 <= reg671;
              if ($unsigned((^$signed((~&reg666)))))
                begin
                  if ($unsigned(reg672))
                    begin
                      reg697 = (reg669 ?
                          forvar685[(1'h1):(1'h0)] : (($unsigned(reg691) ?
                                  forvar685[(1'h0):(1'h0)] : {reg668}) ?
                              (&(^~reg690)) : {""}));
                      reg698 = (~&($signed($unsigned(forvar663)) ?
                          reg659 : (-forvar671[(1'h1):(1'h1)])));
                      reg699 <= $signed((-reg660[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg697 = reg680[(2'h3):(2'h3)];
                      reg699 <= ($unsigned((&$unsigned(reg677))) <= {(!reg657[(1'h0):(1'h0)])});
                    end
                  for (forvar700 = (1'h0); (forvar700 < (1'h1)); forvar700 = (forvar700 + (1'h1)))
                    begin
                      reg701 <= "KDO";
                    end
                end
              else
                begin
                  for (forvar697 = (1'h0); (forvar697 < (1'h0)); forvar697 = (forvar697 + (1'h1)))
                    begin
                      reg698 = $unsigned("y");
                    end
                  if (forvar661)
                    begin
                      reg699 <= $unsigned("SINS4oJaPF0");
                    end
                  else
                    begin
                      reg700 = {(wire653[(1'h1):(1'h0)] * forvar667)};
                      reg702 = reg688;
                      reg703 = $unsigned(($signed((|reg691)) ^~ "cS234r"));
                      reg704 <= (~&(reg677 ?
                          reg657 : $unsigned((reg662 <= reg687))));
                    end
                  for (forvar705 = (1'h0); (forvar705 < (2'h2)); forvar705 = (forvar705 + (1'h1)))
                    begin
                      reg706 <= "";
                      reg707 = {$signed((&wire652[(1'h1):(1'h0)]))};
                      reg708 <= ((&reg684[(1'h0):(1'h0)]) ?
                          (forvar661 ?
                              {(forvar692 <= reg681)} : ((reg674 * reg663) && (wire655 ?
                                  reg681 : forvar663))) : reg696[(3'h4):(2'h3)]);
                    end
                  if ((forvar667[(2'h3):(1'h1)] && (^~$unsigned("sFf7CTibB"))))
                    begin
                      reg709 <= forvar658[(1'h0):(1'h0)];
                      reg710 = (8'hb7);
                      reg711 <= "yzYCCkbwb";
                      reg712 = ($unsigned(reg689) ?
                          (|(reg696[(1'h0):(1'h0)] || (reg660 ?
                              reg703 : (8'hb1)))) : (|(((8'h9d) ?
                              reg665 : forvar657) > (reg683 | reg699))));
                    end
                  else
                    begin
                      reg709 <= (forvar705[(3'h6):(1'h1)] == (~($unsigned(forvar686) ^ forvar705)));
                    end
                end
              reg713 = "";
              for (forvar714 = (1'h0); (forvar714 < (1'h1)); forvar714 = (forvar714 + (1'h1)))
                begin
                  reg715 = (((reg708[(3'h6):(1'h1)] ?
                          reg676[(1'h1):(1'h1)] : reg672) ?
                      ({reg676} + (!reg704)) : reg695[(4'hf):(4'h9)]) <<< $signed($unsigned($signed((8'hab)))));
                  for (forvar716 = (1'h0); (forvar716 < (1'h1)); forvar716 = (forvar716 + (1'h1)))
                    begin
                      reg717 = reg694[(1'h0):(1'h0)];
                    end
                  reg718 <= $signed((~|reg660[(3'h5):(3'h5)]));
                end
            end
          else
            begin
              reg696 <= "r";
              reg697 = reg712[(4'h9):(1'h0)];
            end
          for (forvar719 = (1'h0); (forvar719 < (1'h0)); forvar719 = (forvar719 + (1'h1)))
            begin
              for (forvar720 = (1'h0); (forvar720 < (1'h0)); forvar720 = (forvar720 + (1'h1)))
                begin
                  reg721 <= {{reg715}};
                  reg722 <= $unsigned($signed(($signed(reg658) ?
                      reg658 : forvar720[(2'h2):(2'h2)])));
                  for (forvar723 = (1'h0); (forvar723 < (2'h3)); forvar723 = (forvar723 + (1'h1)))
                    begin
                      reg724 <= $signed(($signed((forvar658 == reg691)) ?
                          (~^$signed((8'haa))) : $signed(forvar658[(2'h3):(1'h1)])));
                    end
                end
              for (forvar725 = (1'h0); (forvar725 < (1'h0)); forvar725 = (forvar725 + (1'h1)))
                begin
                  for (forvar726 = (1'h0); (forvar726 < (1'h0)); forvar726 = (forvar726 + (1'h1)))
                    begin
                      reg727 = "AkS891";
                      reg728 = reg701;
                      reg729 <= $unsigned(("HaqQ" ?
                          $signed($signed(reg724)) : $unsigned({reg680})));
                    end
                end
              for (forvar730 = (1'h0); (forvar730 < (1'h0)); forvar730 = (forvar730 + (1'h1)))
                begin
                  for (forvar731 = (1'h0); (forvar731 < (1'h1)); forvar731 = (forvar731 + (1'h1)))
                    begin
                      reg732 <= forvar730;
                      reg733 <= (~&(!((8'hb3) <<< {forvar685})));
                      reg734 = ((reg709 ?
                          (~^(reg680 - reg718)) : (|$unsigned(reg673))) == $signed(forvar705));
                    end
                  reg735 = forvar697;
                end
            end
        end
      else
        begin
          for (forvar696 = (1'h0); (forvar696 < (1'h1)); forvar696 = (forvar696 + (1'h1)))
            begin
              reg697 = "4GQ";
            end
          for (forvar698 = (1'h0); (forvar698 < (2'h2)); forvar698 = (forvar698 + (1'h1)))
            begin
              for (forvar699 = (1'h0); (forvar699 < (1'h0)); forvar699 = (forvar699 + (1'h1)))
                begin
                  for (forvar700 = (1'h0); (forvar700 < (1'h1)); forvar700 = (forvar700 + (1'h1)))
                    begin
                      reg702 = (reg735 ?
                          $signed(((forvar730 + reg672) ?
                              $signed(wire652) : (-forvar731))) : (($unsigned(reg659) ?
                                  (&reg734) : ((8'hb4) ? forvar698 : (8'hb5))) ?
                              ($signed(reg657) != (reg679 < reg668)) : (8'h9e)));
                    end
                end
              if (forvar730[(4'ha):(3'h6)])
                begin
                  if (reg733[(2'h3):(1'h0)])
                    begin
                      reg704 <= (($unsigned({forvar698}) ?
                          $unsigned(reg704) : ((^~(8'hb9)) >>> forvar725)) - (reg733[(2'h3):(1'h0)] > $signed(reg694)));
                      reg705 = ((forvar723 ^~ $signed(reg699)) && forvar697);
                    end
                  else
                    begin
                      reg703 = (reg694 ?
                          $unsigned("wqMJV952N") : (^($unsigned(reg696) ?
                              (forvar671 >= reg696) : (~wire655))));
                      reg705 = reg676[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  if (({($signed(reg717) - $unsigned(reg735))} ?
                      reg734[(4'h9):(4'h9)] : $unsigned((~^$signed(reg668)))))
                    begin
                      reg703 = "BiUk";
                      reg704 <= (8'hb8);
                      reg705 = reg699;
                    end
                  else
                    begin
                      reg704 <= ($signed(reg732) ?
                          "aluFRCOgXnH" : ($signed($unsigned(reg722)) ?
                              reg672[(3'h4):(3'h4)] : (reg687 ^~ (^~reg669))));
                      reg705 = (8'hab);
                      reg707 = {(~^(+$unsigned(reg664)))};
                      reg710 = $unsigned(((forvar685[(3'h7):(1'h1)] ?
                          (~(8'hb2)) : wire652) * reg713[(4'h8):(2'h3)]));
                    end
                  reg712 = ("nYTveAh15i" ?
                      ("yo7eB" ?
                          ($signed(reg705) * reg682[(4'ha):(3'h6)]) : $signed($unsigned(forvar698))) : (($signed(reg715) - $unsigned(forvar705)) != "bF2wNVWFeeVtH"));
                  reg713 = $signed(reg667[(3'h6):(1'h1)]);
                end
            end
          reg714 = ($signed($signed(((8'hba) ?
              reg670 : (8'hb2)))) || reg690[(2'h3):(2'h2)]);
        end
      reg736 <= reg662;
    end
  assign wire737 = $signed({$signed({reg667})});
  always
    @(posedge clk) begin
      for (forvar738 = (1'h0); (forvar738 < (2'h2)); forvar738 = (forvar738 + (1'h1)))
        begin
          for (forvar739 = (1'h0); (forvar739 < (2'h3)); forvar739 = (forvar739 + (1'h1)))
            begin
              reg740 <= (~^("FK8RxX5y8NaLTmW" << wire655[(3'h6):(1'h0)]));
            end
          reg741 = $signed({({reg677} && (~|forvar738))});
        end
      if (((8'hae) >>> {((+forvar738) ?
              reg722[(4'ha):(4'h9)] : $unsigned(reg733))}))
        begin
          reg742 = reg701;
        end
      else
        begin
          if ({(8'hb8)})
            begin
              if ($signed(((reg667 > (^reg665)) ?
                  (8'h9d) : (~|(reg661 ? reg704 : (8'ha1))))))
                begin
                  if (reg733[(1'h0):(1'h0)])
                    begin
                      reg742 = $signed($unsigned((^~(reg668 ?
                          reg691 : wire737))));
                      reg743 = {(~&$unsigned(reg683))};
                      reg744 <= $signed((reg669 ~^ reg696[(2'h3):(2'h2)]));
                      reg745 = reg678;
                    end
                  else
                    begin
                      reg744 <= $unsigned($signed(reg699));
                      reg745 = (reg741 ?
                          $signed((reg709[(4'h9):(1'h1)] - ((8'hb2) == wire737))) : reg677);
                      reg746 <= ({$unsigned((~reg667))} ^~ ({(~|reg681)} ?
                          wire653 : {"eak9F2b0ztc4"}));
                      reg747 <= (^~(&{(reg732 < (8'hb4))}));
                    end
                  for (forvar748 = (1'h0); (forvar748 < (1'h0)); forvar748 = (forvar748 + (1'h1)))
                    begin
                      reg749 = $unsigned(reg681);
                      reg750 <= $unsigned(reg706);
                      reg751 = {reg665[(1'h0):(1'h0)]};
                      reg752 <= (|(|(|(reg750 < reg667))));
                    end
                end
              else
                begin
                  reg742 = (reg750 ? "J" : "ZAT5pYpSuDx");
                end
              if (((($unsigned((8'ha0)) ?
                  (~^reg709) : (^~(8'h9f))) <<< "dQGXNYMTI") & reg721))
                begin
                  if ("9pOYFow9axvW")
                    begin
                      reg753 = reg711[(4'hb):(4'h9)];
                      reg754 <= {reg701[(3'h4):(2'h3)]};
                      reg755 <= $signed(reg753);
                    end
                  else
                    begin
                      reg754 <= ((($unsigned(reg684) | reg662) ?
                              (~&(reg699 ?
                                  reg751 : (8'hb6))) : $unsigned((&reg704))) ?
                          $unsigned((~{reg669})) : ({"6cxrnadCpcW"} ?
                              ((wire655 == reg684) ?
                                  (8'hb0) : reg733) : ((8'h9d) ?
                                  "q5hx5Y4KvEFlWT3" : reg684[(1'h1):(1'h0)])));
                      reg755 <= $unsigned((($signed(reg742) ^ reg724) ?
                          $unsigned((reg745 ?
                              (8'h9f) : reg709)) : $unsigned((reg678 ?
                              reg683 : reg681))));
                      reg756 = reg685[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar753 = (1'h0); (forvar753 < (2'h2)); forvar753 = (forvar753 + (1'h1)))
                    begin
                      reg754 <= (reg753[(2'h2):(1'h1)] ? "ILFgZdLKt" : "BU2WT");
                    end
                  for (forvar755 = (1'h0); (forvar755 < (1'h1)); forvar755 = (forvar755 + (1'h1)))
                    begin
                      reg757 <= {wire737};
                      reg758 <= {"XcfZBFBD8E74"};
                      reg759 = ("bYgBxuRyTy9" && reg701);
                      reg760 = (~$signed(((reg709 ? reg753 : reg744) ?
                          (forvar755 || reg744) : (reg684 >= reg759))));
                    end
                  for (forvar761 = (1'h0); (forvar761 < (2'h3)); forvar761 = (forvar761 + (1'h1)))
                    begin
                      reg762 = $unsigned(($unsigned((reg699 << reg741)) <= reg704[(1'h1):(1'h0)]));
                      reg763 = $signed(($unsigned(reg744) ^ $unsigned((reg699 << reg709))));
                      reg764 = ((-(&(reg755 ? reg665 : reg743))) ?
                          (reg691[(3'h5):(3'h4)] <<< (^~{reg756})) : ({(^~wire655)} * $unsigned({(8'hb2)})));
                    end
                end
              reg765 = {"h1HipYAkNB2vO"};
            end
          else
            begin
              for (forvar742 = (1'h0); (forvar742 < (1'h0)); forvar742 = (forvar742 + (1'h1)))
                begin
                  for (forvar743 = (1'h0); (forvar743 < (2'h3)); forvar743 = (forvar743 + (1'h1)))
                    begin
                      reg744 <= (reg684 ?
                          (-(~&(reg686 >> reg677))) : ($unsigned($unsigned((8'ha1))) ?
                              (8'hb6) : (~^{reg673})));
                      reg745 = (wire653[(2'h3):(2'h2)] ?
                          "uEtuI" : reg665[(1'h0):(1'h0)]);
                      reg746 <= $unsigned($unsigned(forvar742));
                      reg747 <= ("SGZp3izk2v94R" ?
                          ($unsigned($signed(reg752)) ?
                              reg729 : "ixBHJ") : reg677);
                    end
                  for (forvar748 = (1'h0); (forvar748 < (2'h3)); forvar748 = (forvar748 + (1'h1)))
                    begin
                      reg749 = ((((reg724 ? forvar755 : reg686) ?
                                  (reg677 + reg736) : $signed(reg757)) ?
                              $signed(forvar748[(4'ha):(3'h5)]) : forvar742) ?
                          reg686 : reg736[(3'h6):(3'h4)]);
                      reg750 <= reg757[(1'h0):(1'h0)];
                      reg751 = $unsigned((8'h9c));
                      reg752 <= "2kwVbUMAtLxx";
                    end
                  for (forvar753 = (1'h0); (forvar753 < (1'h0)); forvar753 = (forvar753 + (1'h1)))
                    begin
                      reg754 <= {reg746[(2'h2):(1'h1)]};
                      reg756 = (((&(~^reg677)) ?
                              reg751 : reg736[(2'h3):(1'h0)]) ?
                          reg704 : ((+(~&reg760)) && "QZqXuZf7"));
                      reg757 <= (reg678[(2'h3):(1'h0)] ?
                          (("rYVl7HUxrIbLH4" ?
                              (reg729 ~^ wire654) : (reg689 ?
                                  reg683 : reg745)) | ($signed(reg747) ^ reg729)) : reg678);
                      reg759 = reg764[(1'h0):(1'h0)];
                    end
                  for (forvar760 = (1'h0); (forvar760 < (1'h0)); forvar760 = (forvar760 + (1'h1)))
                    begin
                      reg761 = ((reg681[(2'h3):(2'h3)] ?
                              reg740 : "y07pAALkA8") ?
                          "ZT3OxJLGqRT" : "Q0c9o");
                      reg762 = $signed($unsigned(((reg747 & forvar738) << $signed(reg744))));
                      reg763 = $signed((|(^{wire655})));
                    end
                end
            end
          for (forvar766 = (1'h0); (forvar766 < (1'h0)); forvar766 = (forvar766 + (1'h1)))
            begin
              for (forvar767 = (1'h0); (forvar767 < (1'h0)); forvar767 = (forvar767 + (1'h1)))
                begin
                  reg768 = $signed((!((reg758 ? forvar753 : reg685) ?
                      reg762 : reg744)));
                  if ($unsigned(wire655))
                    begin
                      reg769 = $signed(reg699);
                      reg770 = ({$unsigned((8'hb0))} & wire656[(1'h1):(1'h1)]);
                      reg771 = "MfO9VtbHUOBm";
                      reg772 = ((^~((reg721 ? reg743 : reg759) ?
                              reg706 : $signed(reg685))) ?
                          $unsigned(((8'hba) ?
                              wire656 : $unsigned(reg724))) : reg762);
                    end
                  else
                    begin
                      reg769 = reg729[(2'h2):(1'h1)];
                      reg773 <= reg681[(1'h0):(1'h0)];
                      reg774 = $signed({$unsigned((~reg741))});
                      reg775 <= (~|(&{((8'ha3) - reg662)}));
                    end
                end
              reg776 = forvar766;
            end
          reg777 = reg756;
        end
      for (forvar778 = (1'h0); (forvar778 < (2'h3)); forvar778 = (forvar778 + (1'h1)))
        begin
          reg779 = (&reg709[(4'hd):(3'h6)]);
          for (forvar780 = (1'h0); (forvar780 < (1'h1)); forvar780 = (forvar780 + (1'h1)))
            begin
              reg781 <= ("m" ?
                  "dz5U816u" : ($unsigned(((8'hb5) ? (8'had) : reg722)) ?
                      "QxZg" : $signed($signed((8'had)))));
              reg782 = reg706;
            end
          for (forvar783 = (1'h0); (forvar783 < (2'h2)); forvar783 = (forvar783 + (1'h1)))
            begin
              reg784 <= reg763[(3'h4):(2'h2)];
              for (forvar785 = (1'h0); (forvar785 < (1'h1)); forvar785 = (forvar785 + (1'h1)))
                begin
                  reg786 <= (reg743[(3'h5):(2'h2)] >>> reg772);
                  if ((reg752 ?
                      ($unsigned(reg701[(3'h4):(1'h0)]) ?
                          (reg765[(2'h2):(1'h1)] ?
                              "OsWRxqyxskhcuiL" : reg758) : (~(wire737 >>> (8'ha9)))) : ({reg777} ?
                          reg681 : $unsigned("nak"))))
                    begin
                      reg787 = (&(({reg764} ?
                          {reg668} : forvar743) == wire655[(3'h5):(3'h5)]));
                    end
                  else
                    begin
                      reg787 = $signed((&$signed($unsigned((8'h9e)))));
                      reg788 = $unsigned((reg732 != $unsigned((reg706 ?
                          wire654 : (8'hba)))));
                      reg789 = $unsigned(reg721[(1'h1):(1'h1)]);
                    end
                  reg790 = ($unsigned($unsigned("MkDGvlK5En")) ^~ "Iw1DXNIUxaZkSI2");
                  for (forvar791 = (1'h0); (forvar791 < (1'h1)); forvar791 = (forvar791 + (1'h1)))
                    begin
                      reg792 <= reg762;
                      reg793 <= "30l";
                      reg794 <= (!$signed($signed($unsigned((8'hb6)))));
                    end
                end
              for (forvar795 = (1'h0); (forvar795 < (1'h0)); forvar795 = (forvar795 + (1'h1)))
                begin
                  reg796 = forvar783[(1'h1):(1'h1)];
                  reg797 = reg774[(1'h1):(1'h0)];
                end
              reg798 = (~&(reg668 ?
                  ((reg701 + reg661) ?
                      ((8'hb0) + reg746) : (reg793 < (8'hb6))) : ($unsigned(reg668) ?
                      forvar753 : $signed(reg662))));
            end
          for (forvar799 = (1'h0); (forvar799 < (1'h1)); forvar799 = (forvar799 + (1'h1)))
            begin
              for (forvar800 = (1'h0); (forvar800 < (2'h3)); forvar800 = (forvar800 + (1'h1)))
                begin
                  reg801 = "gyeW";
                  for (forvar802 = (1'h0); (forvar802 < (2'h2)); forvar802 = (forvar802 + (1'h1)))
                    begin
                      reg803 = reg736[(1'h1):(1'h0)];
                    end
                  reg804 <= ((((reg718 ? reg770 : reg793) ?
                              {reg751} : $unsigned(reg752)) ?
                          wire656[(3'h5):(1'h0)] : {reg684}) ?
                      (~&(^~((8'hb0) >= reg749))) : ((|"IDoA") ^~ ""));
                  for (forvar805 = (1'h0); (forvar805 < (2'h2)); forvar805 = (forvar805 + (1'h1)))
                    begin
                      reg806 = ($unsigned((+reg788[(2'h2):(1'h0)])) < $signed($unsigned($unsigned(reg775))));
                      reg807 = ("5g2" ?
                          $signed(($unsigned(reg733) ?
                              reg701 : reg685[(4'hb):(4'h8)])) : reg661[(1'h0):(1'h0)]);
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      reg808 <= reg689;
    end
  always
    @(posedge clk) begin
      reg809 <= $unsigned(reg699[(3'h4):(3'h4)]);
      if (reg683)
        begin
          for (forvar810 = (1'h0); (forvar810 < (1'h1)); forvar810 = (forvar810 + (1'h1)))
            begin
              for (forvar811 = (1'h0); (forvar811 < (1'h0)); forvar811 = (forvar811 + (1'h1)))
                begin
                  reg812 = {reg755};
                  for (forvar813 = (1'h0); (forvar813 < (2'h3)); forvar813 = (forvar813 + (1'h1)))
                    begin
                      reg814 <= ("PWrNW2f5wqstsOo" ?
                          ($unsigned((!reg808)) ?
                              ({reg793} ?
                                  (reg664 ?
                                      reg711 : reg740) : (~&wire654)) : $unsigned($signed(reg699))) : "mwQUO");
                      reg815 = reg750[(3'h4):(2'h2)];
                    end
                  reg816 = $unsigned(($unsigned(reg792[(4'hb):(4'h9)]) || ((reg681 == reg701) ?
                      (reg746 - (8'hab)) : $signed(wire737))));
                  reg817 = (($signed(reg721) ?
                      $signed((reg678 ?
                          reg781 : reg665)) : ((&reg794) & reg699[(3'h4):(1'h0)])) >= reg665);
                end
              if ($unsigned($unsigned(reg784[(3'h4):(3'h4)])))
                begin
                  reg818 <= reg794;
                  for (forvar819 = (1'h0); (forvar819 < (2'h2)); forvar819 = (forvar819 + (1'h1)))
                    begin
                      reg820 <= ({$signed(wire655[(4'h9):(1'h1)])} ?
                          ($unsigned((forvar819 * reg683)) ?
                              ($signed(reg686) ?
                                  wire653 : (-reg662)) : $unsigned((reg815 ?
                                  reg683 : reg658))) : reg746[(2'h2):(1'h0)]);
                      reg821 <= wire737[(1'h0):(1'h0)];
                      reg822 = (reg758[(2'h3):(2'h3)] ?
                          reg681[(3'h4):(2'h3)] : (^~(reg689 ?
                              ((8'hba) ?
                                  reg758 : (8'hab)) : $signed((8'ha6)))));
                      reg823 <= (^reg677);
                    end
                  for (forvar824 = (1'h0); (forvar824 < (2'h2)); forvar824 = (forvar824 + (1'h1)))
                    begin
                      reg825 <= (({reg681} ?
                          $signed($unsigned(reg733)) : (~(~wire655))) >>> ((forvar811 >>> reg665[(2'h3):(2'h2)]) ?
                          reg665 : {(reg750 >= reg804)}));
                      reg826 = ((reg718[(1'h1):(1'h0)] * reg706[(4'he):(2'h3)]) ?
                          wire652[(2'h3):(2'h3)] : ($signed($unsigned(reg732)) ?
                              $unsigned(((8'had) ?
                                  reg754 : forvar819)) : (+(reg758 ?
                                  reg711 : reg821))));
                      reg827 = $signed((!reg699[(2'h3):(2'h3)]));
                    end
                  if (forvar819[(3'h6):(3'h5)])
                    begin
                      reg828 = ((&reg817[(3'h4):(1'h1)]) ^~ $unsigned({$signed(reg752)}));
                      reg829 = ((({reg822} <<< (-(8'hb3))) ?
                          ((^~reg664) | reg746[(3'h4):(1'h1)]) : reg808) & ("EJNF1o" ^~ forvar811));
                    end
                  else
                    begin
                      reg828 = reg827;
                      reg830 <= $signed((8'ha3));
                      reg831 = $unsigned($signed((&$unsigned((8'had)))));
                      reg832 = {$unsigned((~{reg804}))};
                    end
                end
              else
                begin
                  reg819 = ({$unsigned((+wire655))} * reg694);
                end
              if ((&(&reg752)))
                begin
                  for (forvar833 = (1'h0); (forvar833 < (2'h3)); forvar833 = (forvar833 + (1'h1)))
                    begin
                      reg834 = "pVdRp8kK3no9Tq";
                      reg835 <= $signed($unsigned((^~(reg808 ?
                          (8'hb1) : reg815))));
                      reg836 <= reg677[(1'h1):(1'h1)];
                    end
                  for (forvar837 = (1'h0); (forvar837 < (2'h2)); forvar837 = (forvar837 + (1'h1)))
                    begin
                      reg838 = {(8'h9d)};
                      reg839 <= (reg722 ^~ ((|reg822[(1'h1):(1'h0)]) <= ((~&(8'ha5)) < $unsigned((8'ha3)))));
                      reg840 = ((8'hb0) < (~$unsigned($unsigned(reg736))));
                      reg841 = "wWBiCtEmku";
                    end
                end
              else
                begin
                  if (reg662[(4'h8):(1'h1)])
                    begin
                      reg833 = {({reg838} & {$signed(wire654)})};
                      reg834 = reg694;
                      reg835 <= reg708[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg835 <= $unsigned($signed(reg830[(2'h3):(2'h3)]));
                      reg837 = $signed(reg699[(2'h2):(1'h0)]);
                      reg838 = reg804;
                    end
                  reg840 = {$unsigned(reg718[(3'h6):(3'h4)])};
                end
              for (forvar842 = (1'h0); (forvar842 < (1'h1)); forvar842 = (forvar842 + (1'h1)))
                begin
                  reg843 = (~(8'ha7));
                  reg844 = (forvar810 ?
                      $unsigned("L6hTW53l") : (-((^~reg733) - reg747[(3'h4):(3'h4)])));
                  for (forvar845 = (1'h0); (forvar845 < (2'h3)); forvar845 = (forvar845 + (1'h1)))
                    begin
                      reg846 = reg754[(3'h7):(1'h0)];
                      reg847 <= (-reg752);
                      reg848 = ((8'hac) ?
                          (~&((^reg804) ?
                              "g9WLwq0htQrwB1" : ((8'ha2) <<< reg819))) : (reg818[(4'h8):(1'h0)] ^~ (8'ha8)));
                      reg849 = reg833;
                    end
                  if (reg696[(2'h3):(1'h0)])
                    begin
                      reg850 <= (^(reg706 ^~ $unsigned((reg846 ~^ reg830))));
                      reg851 <= $unsigned((reg699[(3'h4):(3'h4)] ?
                          (~^reg815) : {(~&reg792)}));
                      reg852 = $signed($signed((forvar811[(4'h9):(2'h2)] ?
                          forvar824[(2'h2):(1'h0)] : reg826)));
                      reg853 = (!{{"XBRs7y2QSwL"}});
                    end
                  else
                    begin
                      reg852 = {reg755[(3'h7):(2'h2)]};
                      reg853 = (((~&reg831) == $unsigned((reg775 ^ (8'ha2)))) != {($unsigned(reg848) ?
                              $unsigned(wire653) : reg696[(3'h6):(2'h2)])});
                    end
                end
            end
          reg854 <= ({(!reg849[(3'h6):(3'h5)])} >> $unsigned($signed($signed(reg683))));
          reg855 <= ((!($unsigned(reg668) <= reg804)) ?
              ($signed((reg754 ^~ reg669)) ?
                  "dgbeJHJ" : "2v2iPzwEkQuw3Xh") : $unsigned((forvar833[(3'h5):(3'h5)] || reg828)));
        end
      else
        begin
          for (forvar810 = (1'h0); (forvar810 < (1'h1)); forvar810 = (forvar810 + (1'h1)))
            begin
              if (("aXebl" ? reg822[(4'ha):(1'h0)] : (~reg754)))
                begin
                  for (forvar811 = (1'h0); (forvar811 < (2'h2)); forvar811 = (forvar811 + (1'h1)))
                    begin
                      reg813 <= $unsigned($unsigned(($unsigned(reg729) << $signed(forvar813))));
                      reg814 <= forvar813[(1'h1):(1'h1)];
                    end
                  for (forvar815 = (1'h0); (forvar815 < (2'h3)); forvar815 = (forvar815 + (1'h1)))
                    begin
                      reg816 = $unsigned(forvar813);
                      reg817 = {reg662};
                      reg819 = (~reg847[(5'h10):(4'ha)]);
                    end
                  reg822 = forvar819[(4'h8):(2'h3)];
                  reg824 = ((($signed(reg754) >> ((8'hb9) ?
                              forvar815 : wire737)) ?
                          $signed(reg699[(2'h3):(2'h2)]) : $signed($signed(reg750))) ?
                      $unsigned(reg732) : {reg661[(3'h5):(2'h2)]});
                end
              else
                begin
                  reg811 <= (($unsigned($unsigned(reg736)) >= "4vQJYyl") >>> ({$signed(reg701)} ?
                      $unsigned((reg824 != (8'hac))) : reg855[(2'h2):(1'h1)]));
                end
              for (forvar825 = (1'h0); (forvar825 < (2'h2)); forvar825 = (forvar825 + (1'h1)))
                begin
                  if ($signed({$unsigned((wire655 * reg744))}))
                    begin
                      reg826 = "dcIhF";
                      reg830 <= {reg667[(1'h1):(1'h1)]};
                      reg831 = ((reg678[(1'h1):(1'h1)] >= ($unsigned(reg828) > $unsigned(reg855))) ?
                          $unsigned($signed($unsigned(reg729))) : "Jg1iZu5cQp09");
                    end
                  else
                    begin
                      reg830 <= (8'hb1);
                      reg831 = (&reg837);
                      reg832 = (^~(reg825[(3'h4):(1'h0)] ?
                          $signed((reg685 ?
                              reg758 : reg706)) : wire655[(4'hd):(3'h6)]));
                      reg833 = (8'ha1);
                    end
                  reg834 = {$signed(wire653)};
                  for (forvar835 = (1'h0); (forvar835 < (1'h1)); forvar835 = (forvar835 + (1'h1)))
                    begin
                      reg837 = $unsigned((((forvar845 ? (8'hb5) : reg811) ?
                              ((8'ha9) >> reg829) : reg841[(4'hb):(4'h8)]) ?
                          (^~$signed((8'ha4))) : (~&(~^(8'hba)))));
                      reg838 = reg729;
                    end
                  reg840 = $unsigned((+reg831));
                end
            end
          for (forvar841 = (1'h0); (forvar841 < (2'h2)); forvar841 = (forvar841 + (1'h1)))
            begin
              if ("4yWRXsdiuoXE")
                begin
                  if ({$unsigned($unsigned((reg850 >> reg664)))})
                    begin
                      reg842 <= $signed(reg828);
                      reg843 = reg786;
                      reg844 = reg721;
                      reg845 <= $signed($unsigned(reg773));
                    end
                  else
                    begin
                      reg842 <= "snp2Iuh4EbeWU";
                      reg845 <= reg740;
                    end
                  reg846 = $signed(forvar813);
                end
              else
                begin
                  for (forvar842 = (1'h0); (forvar842 < (2'h3)); forvar842 = (forvar842 + (1'h1)))
                    begin
                      reg843 = reg721[(2'h3):(1'h0)];
                      reg845 <= reg658;
                      reg847 <= reg757;
                      reg848 = wire652[(1'h1):(1'h0)];
                    end
                end
              reg850 <= (8'hb8);
              for (forvar851 = (1'h0); (forvar851 < (2'h2)); forvar851 = (forvar851 + (1'h1)))
                begin
                  reg852 = $unsigned($signed(((8'ha4) == forvar845)));
                end
              for (forvar853 = (1'h0); (forvar853 < (2'h2)); forvar853 = (forvar853 + (1'h1)))
                begin
                  if ({$unsigned(($unsigned(reg833) ^~ $signed(forvar853)))})
                    begin
                      reg856 = $signed("Vs91736XtLq");
                      reg857 = reg834[(3'h7):(3'h6)];
                      reg858 <= reg696;
                    end
                  else
                    begin
                      reg856 = (forvar842 ?
                          reg752[(2'h2):(2'h2)] : (forvar842 > ({wire656} ?
                              {reg829} : {reg708})));
                      reg857 = $signed($unsigned((reg732[(1'h1):(1'h0)] ?
                          (reg829 ? reg815 : reg843) : $signed(reg746))));
                    end
                  reg859 <= $signed($signed(reg833[(4'hb):(2'h3)]));
                  for (forvar860 = (1'h0); (forvar860 < (1'h0)); forvar860 = (forvar860 + (1'h1)))
                    begin
                      reg861 = wire652[(2'h2):(2'h2)];
                      reg862 = reg711[(1'h0):(1'h0)];
                      reg863 <= $unsigned({(reg662 - reg827)});
                      reg864 <= ($unsigned(reg850[(1'h1):(1'h0)]) + $unsigned(($unsigned(reg752) ?
                          reg732 : $signed(reg683))));
                    end
                  if (((~$unsigned(((8'hb5) ?
                      reg658 : (8'ha0)))) ^~ reg747[(2'h3):(1'h0)]))
                    begin
                      reg865 <= reg662;
                      reg866 = $unsigned($unsigned(((&reg814) & reg669[(2'h2):(2'h2)])));
                      reg867 <= {$unsigned(($unsigned(reg811) < {(8'hb4)}))};
                    end
                  else
                    begin
                      reg866 = {$signed((reg836 ?
                              reg862[(3'h5):(2'h2)] : $signed(reg834)))};
                    end
                end
            end
          if ({$signed(reg694)})
            begin
              if ((8'hb1))
                begin
                  reg868 = reg793[(2'h2):(2'h2)];
                  if ($unsigned($unsigned(reg857)))
                    begin
                      reg869 = (~|forvar845[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg869 = $unsigned(forvar825);
                      reg870 = (($signed({reg827}) <<< "DDiKvsd92a0E7m") ?
                          (~($signed(reg691) ?
                              reg858[(2'h2):(2'h2)] : (8'had))) : $unsigned(reg664[(2'h2):(2'h2)]));
                      reg871 <= (!$unsigned({reg662[(2'h2):(2'h2)]}));
                    end
                  for (forvar872 = (1'h0); (forvar872 < (1'h1)); forvar872 = (forvar872 + (1'h1)))
                    begin
                      reg873 <= $unsigned((forvar833 & $signed((!forvar837))));
                      reg874 = {$signed("GmFmzueUyEOm")};
                      reg875 <= ($unsigned((&$unsigned(forvar860))) ?
                          reg861 : "MUb8HC");
                      reg876 <= reg868[(4'h8):(3'h5)];
                    end
                  reg877 <= $signed((reg793 >>> reg876[(3'h7):(2'h2)]));
                end
              else
                begin
                  if ($unsigned(reg733[(2'h3):(2'h3)]))
                    begin
                      reg871 <= (reg844[(4'hb):(3'h6)] ?
                          $signed($signed((reg842 ^ reg792))) : $signed((8'ha7)));
                      reg872 = reg775[(4'ha):(1'h0)];
                      reg874 = {$unsigned((-(reg875 > reg866)))};
                    end
                  else
                    begin
                      reg868 = (((-(^~reg658)) ?
                              (-forvar842[(3'h7):(2'h3)]) : {(reg856 ?
                                      forvar811 : reg832)}) ?
                          (8'ha2) : (^~("R5l1Vy" ?
                              (+forvar833) : $signed(reg792))));
                      reg869 = $unsigned(wire653);
                      reg871 <= (^(({reg775} ?
                          {reg775} : "QpP5Ov5QZNMa") & $unsigned((reg835 < reg721))));
                      reg872 = reg733[(2'h2):(2'h2)];
                    end
                  if ((8'hb1))
                    begin
                      reg875 <= $unsigned(reg775[(3'h6):(3'h5)]);
                      reg878 = ((&reg808) ?
                          reg818[(1'h1):(1'h1)] : reg685[(2'h3):(1'h1)]);
                      reg879 <= {reg851[(3'h7):(3'h4)]};
                    end
                  else
                    begin
                      reg878 = ((($signed(forvar845) && $unsigned(reg843)) >= (^~{reg724})) ?
                          {$unsigned((reg732 + forvar837))} : ($signed($signed(reg839)) || $signed((-reg669))));
                      reg879 <= reg875;
                      reg880 = {reg677};
                      reg881 = $unsigned($unsigned($signed({reg872})));
                    end
                end
              for (forvar882 = (1'h0); (forvar882 < (1'h0)); forvar882 = (forvar882 + (1'h1)))
                begin
                  reg883 <= $unsigned("D4BXzOdfXgA");
                  reg884 <= $unsigned(($signed((~&reg871)) > {(reg853 ^~ reg881)}));
                end
              for (forvar885 = (1'h0); (forvar885 < (2'h3)); forvar885 = (forvar885 + (1'h1)))
                begin
                  for (forvar886 = (1'h0); (forvar886 < (1'h1)); forvar886 = (forvar886 + (1'h1)))
                    begin
                      reg887 = (reg732[(1'h1):(1'h1)] * (-(+$signed(reg784))));
                      reg888 <= (^{$signed({reg662})});
                    end
                  reg889 = $unsigned(($signed($unsigned(reg662)) ?
                      reg845 : ((reg871 + reg701) * forvar845)));
                  for (forvar890 = (1'h0); (forvar890 < (2'h3)); forvar890 = (forvar890 + (1'h1)))
                    begin
                      reg891 = $signed("RRieLVx4");
                    end
                end
            end
          else
            begin
              reg868 = reg854[(3'h7):(2'h2)];
              reg871 <= reg854[(3'h7):(3'h7)];
              if ($signed(("pWWopYne" >> reg868)))
                begin
                  for (forvar872 = (1'h0); (forvar872 < (2'h2)); forvar872 = (forvar872 + (1'h1)))
                    begin
                      reg874 = ((((reg809 ? reg683 : reg816) > forvar824) ?
                          $signed((forvar835 ?
                              reg699 : reg889)) : (^~$unsigned(reg683))) - reg718);
                    end
                  reg875 <= $signed(reg781);
                  for (forvar876 = (1'h0); (forvar876 < (1'h0)); forvar876 = (forvar876 + (1'h1)))
                    begin
                      reg878 = $unsigned(((^$signed((8'hb3))) ?
                          ((~^reg665) ?
                              reg732[(4'h8):(3'h7)] : reg709) : ((reg786 ?
                                  (8'hac) : (8'h9c)) ?
                              (|reg673) : (forvar841 ^ (8'ha3)))));
                      reg879 <= $unsigned($signed($signed(wire737)));
                      reg882 <= (forvar835[(4'hf):(4'hc)] * ("q9YUQOBtFKMSc" ?
                          reg784[(1'h0):(1'h0)] : reg665[(1'h0):(1'h0)]));
                      reg885 = (8'hae);
                    end
                  for (forvar886 = (1'h0); (forvar886 < (2'h2)); forvar886 = (forvar886 + (1'h1)))
                    begin
                      reg888 <= reg815[(1'h1):(1'h1)];
                      reg890 <= {reg889};
                    end
                end
              else
                begin
                  for (forvar872 = (1'h0); (forvar872 < (2'h2)); forvar872 = (forvar872 + (1'h1)))
                    begin
                      reg874 = (&($unsigned($unsigned(forvar841)) ?
                          $unsigned($signed(wire737)) : {{reg836}}));
                      reg878 = (&($signed({reg708}) ^~ (~(reg686 ?
                          reg870 : reg857))));
                    end
                  reg880 = {((~|"O1xGGkiET6O") ?
                          reg885[(4'hd):(3'h6)] : reg808)};
                  reg881 = {(-reg890[(1'h0):(1'h0)])};
                  for (forvar882 = (1'h0); (forvar882 < (1'h1)); forvar882 = (forvar882 + (1'h1)))
                    begin
                      reg885 = "t9iR";
                    end
                end
              if ({$signed($signed((reg855 ? reg819 : forvar842)))})
                begin
                  for (forvar891 = (1'h0); (forvar891 < (2'h2)); forvar891 = (forvar891 + (1'h1)))
                    begin
                      reg892 <= $signed(reg662);
                      reg893 = reg689;
                      reg894 = $signed(reg667[(1'h1):(1'h1)]);
                    end
                  for (forvar895 = (1'h0); (forvar895 < (1'h0)); forvar895 = (forvar895 + (1'h1)))
                    begin
                      reg896 = reg821[(2'h2):(1'h1)];
                      reg897 = {$unsigned($signed($unsigned((8'hb6))))};
                      reg898 <= (!({$unsigned(reg859)} ?
                          (~reg754[(4'h8):(3'h4)]) : (8'ha3)));
                      reg899 = reg867[(2'h2):(1'h1)];
                    end
                  for (forvar900 = (1'h0); (forvar900 < (1'h0)); forvar900 = (forvar900 + (1'h1)))
                    begin
                      reg901 = reg887;
                      reg902 <= ($unsigned(($unsigned(reg689) ?
                              $signed((8'ha5)) : $unsigned(forvar837))) ?
                          ({$unsigned(forvar872)} ?
                              {{(8'ha9)}} : "A7zw5T8Ozs") : (&((reg673 ?
                              reg754 : reg667) || ((8'hb9) ?
                              (8'ha9) : reg694))));
                    end
                  for (forvar903 = (1'h0); (forvar903 < (1'h1)); forvar903 = (forvar903 + (1'h1)))
                    begin
                      reg904 = ((~|$unsigned((forvar900 != wire655))) ?
                          "f43X" : reg818);
                      reg905 = ((~reg857) < "6Yw");
                      reg906 = (((~|$unsigned(reg827)) - reg894[(1'h1):(1'h1)]) ?
                          (((|forvar853) ? reg684[(2'h3):(2'h2)] : (~^reg820)) ?
                              ((reg869 ? reg721 : reg833) ?
                                  $signed(reg729) : $unsigned(reg721)) : "O") : reg819[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar891 = (1'h0); (forvar891 < (1'h1)); forvar891 = (forvar891 + (1'h1)))
                    begin
                      reg892 <= reg825;
                      reg895 <= forvar900;
                      reg898 <= reg691[(2'h2):(2'h2)];
                    end
                  reg899 = "Iq2LVRIZ";
                end
            end
        end
      reg907 <= reg843;
      for (forvar908 = (1'h0); (forvar908 < (2'h3)); forvar908 = (forvar908 + (1'h1)))
        begin
          for (forvar909 = (1'h0); (forvar909 < (2'h3)); forvar909 = (forvar909 + (1'h1)))
            begin
              reg910 = reg859;
              reg911 = (forvar810 ?
                  (^~$unsigned(reg901[(3'h4):(3'h4)])) : $unsigned(((|reg661) ?
                      {(8'hae)} : reg827)));
            end
          if ({(reg879[(4'h8):(1'h1)] ^~ ($signed((8'hb4)) ?
                  "HpMc" : ((8'hb0) * reg684)))})
            begin
              reg912 = $unsigned({$unsigned((reg811 ? (8'ha2) : reg673))});
              if ((~|reg842))
                begin
                  for (forvar913 = (1'h0); (forvar913 < (1'h1)); forvar913 = (forvar913 + (1'h1)))
                    begin
                      reg914 <= $signed((^~{(reg864 ? forvar824 : reg704)}));
                      reg915 <= ((8'ha6) ?
                          reg804[(1'h1):(1'h1)] : ("yJPEghrA" ?
                              {reg661} : {$unsigned(reg709)}));
                    end
                  for (forvar916 = (1'h0); (forvar916 < (2'h2)); forvar916 = (forvar916 + (1'h1)))
                    begin
                      reg917 = ($unsigned(((-forvar885) || {reg815})) && (~|reg902));
                      reg918 = $signed($unsigned((~(reg876 < reg813))));
                      reg919 = reg818;
                    end
                  if ({"v0cIwXZe2w2Y674"})
                    begin
                      reg920 = $unsigned(reg878);
                      reg921 <= (8'h9c);
                      reg922 = $unsigned((reg754 ?
                          ((~^reg658) ?
                              $signed(reg825) : (!reg864)) : {reg845[(3'h7):(3'h7)]}));
                      reg923 <= (reg722[(2'h2):(1'h0)] ?
                          reg918 : ("k" ?
                              reg862[(3'h7):(1'h1)] : $unsigned($unsigned(reg848))));
                    end
                  else
                    begin
                      reg921 <= reg685;
                    end
                end
              else
                begin
                  reg913 <= reg839;
                  reg914 <= reg868[(3'h7):(3'h6)];
                  reg916 = (!$signed({$unsigned(reg793)}));
                  reg917 = $unsigned(reg729);
                end
              reg924 <= (reg857 && (+$signed(forvar824)));
              for (forvar925 = (1'h0); (forvar925 < (1'h1)); forvar925 = (forvar925 + (1'h1)))
                begin
                  for (forvar926 = (1'h0); (forvar926 < (2'h3)); forvar926 = (forvar926 + (1'h1)))
                    begin
                      reg927 = $unsigned(($signed(reg912) ?
                          "bMHs7mvfX7Gsk6" : reg899[(4'h8):(2'h2)]));
                      reg928 = reg793[(3'h5):(1'h1)];
                      reg929 <= reg872;
                    end
                  for (forvar930 = (1'h0); (forvar930 < (2'h2)); forvar930 = (forvar930 + (1'h1)))
                    begin
                      reg931 = reg754;
                    end
                  reg932 <= "dS0rkGCal5V";
                end
            end
          else
            begin
              reg913 <= (-(~^($unsigned((8'hb4)) ?
                  (~&(8'haa)) : $unsigned(forvar853))));
            end
          if ((reg894[(1'h1):(1'h0)] > (~^(-(|forvar925)))))
            begin
              reg933 <= reg669[(4'hb):(4'ha)];
              reg934 <= {((-$signed(reg792)) ? reg732 : (!reg809))};
              for (forvar935 = (1'h0); (forvar935 < (2'h3)); forvar935 = (forvar935 + (1'h1)))
                begin
                  reg936 = "usIBtfTWQyo";
                  reg937 <= {(~|reg910)};
                  reg938 = reg794[(4'h9):(3'h6)];
                  reg939 = $unsigned(reg913);
                end
              if ($signed(forvar845))
                begin
                  reg940 = $signed("C");
                  for (forvar941 = (1'h0); (forvar941 < (2'h2)); forvar941 = (forvar941 + (1'h1)))
                    begin
                      reg942 <= ({$signed(forvar853[(4'h8):(4'h8)])} & "w");
                      reg943 <= reg836[(1'h0):(1'h0)];
                      reg944 = reg818[(3'h6):(1'h0)];
                    end
                  reg945 <= {"a"};
                  reg946 = {reg923[(3'h4):(2'h3)]};
                end
              else
                begin
                  reg940 = ((((reg661 + (8'haa)) <= $signed(reg830)) ?
                      $unsigned({forvar882}) : (|reg913[(1'h1):(1'h0)])) == "JT5qeBvQPG");
                  reg941 = $signed((((reg792 ^~ (8'h9f)) ?
                          forvar842[(3'h7):(3'h6)] : reg809) ?
                      (~$signed(reg829)) : $signed((reg784 * (8'hb7)))));
                  if ((~&"6"))
                    begin
                      reg944 = $unsigned(reg831[(1'h0):(1'h0)]);
                      reg946 = (forvar845[(4'hb):(3'h4)] ?
                          reg694[(1'h1):(1'h0)] : reg911);
                    end
                  else
                    begin
                      reg944 = ($signed((|(reg824 <<< reg875))) << $signed(forvar926));
                      reg945 <= "XHTLYKO";
                    end
                  reg947 <= reg847;
                end
            end
          else
            begin
              for (forvar933 = (1'h0); (forvar933 < (1'h0)); forvar933 = (forvar933 + (1'h1)))
                begin
                  if (reg781)
                    begin
                      reg935 = reg875[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg935 = reg696[(4'h8):(2'h2)];
                      reg937 <= $unsigned((8'hb7));
                      reg942 <= (8'h9e);
                    end
                  if ((!$signed(reg815[(2'h2):(1'h0)])))
                    begin
                      reg944 = $signed(reg867[(2'h3):(1'h0)]);
                      reg945 <= "6QL9Db8";
                      reg947 <= $signed(reg941);
                      reg948 = reg850[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg943 <= $signed($signed({(forvar842 > reg927)}));
                      reg945 <= $signed((^~$unsigned({reg914})));
                      reg946 = ({(^{reg878})} ?
                          {"Hq3ICoxEI"} : {((-forvar886) - (~|reg939))});
                      reg948 = $unsigned($signed(reg744[(3'h6):(2'h2)]));
                    end
                  if ($signed(""))
                    begin
                      reg949 = reg936[(3'h5):(1'h0)];
                      reg950 = forvar837[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg951 <= (&("A" & (reg876[(2'h2):(2'h2)] ?
                          (reg939 <= (8'ha0)) : (-reg928))));
                      reg952 = (|$unsigned((+reg881)));
                      reg953 = reg882;
                      reg954 = {$unsigned((~&(8'hac)))};
                    end
                  reg955 = (~^reg848);
                end
              if ($signed($unsigned((~&forvar872))))
                begin
                  reg956 = (~|$unsigned({$unsigned(reg952)}));
                  for (forvar957 = (1'h0); (forvar957 < (2'h2)); forvar957 = (forvar957 + (1'h1)))
                    begin
                      reg958 <= ($signed("yoIAf3QiN250F") ?
                          "uHcIQ7RZu27" : reg870[(2'h2):(2'h2)]);
                    end
                end
              else
                begin
                  if ((((8'haf) == $unsigned((reg941 < forvar903))) ?
                      ($signed($unsigned((8'ha0))) ?
                          reg661[(3'h5):(3'h4)] : $unsigned(((8'haf) == reg936))) : (("lJKQHWD" ?
                          reg755 : (reg924 >> reg665)) < ((&reg704) != reg736))))
                    begin
                      reg957 <= (~^(^$unsigned((reg944 ? forvar872 : reg718))));
                      reg959 = {($signed($unsigned((8'h9c))) ?
                              ($unsigned(reg855) ?
                                  (~|forvar833) : reg696) : (reg917 ?
                                  reg826[(4'ha):(3'h4)] : (~^reg953)))};
                      reg960 = (^~reg812);
                    end
                  else
                    begin
                      reg956 = $signed("olZdIB");
                      reg959 = reg661;
                      reg961 <= (-"cnsd77U82mIL4ic");
                      reg962 = "JqgCpTCmPDM4n";
                    end
                end
              for (forvar963 = (1'h0); (forvar963 < (2'h3)); forvar963 = (forvar963 + (1'h1)))
                begin
                  reg964 = $signed(reg746);
                  if (((-("VHI5dlc8zdqUZ" ?
                          (reg831 ?
                              reg924 : forvar890) : reg792[(4'he):(3'h6)])) ?
                      $unsigned(($unsigned(reg927) ?
                          {reg668} : (reg893 ~^ reg816))) : "hL"))
                    begin
                      reg965 = reg677[(3'h5):(2'h3)];
                      reg966 <= $unsigned((reg934 & $unsigned((!reg879))));
                      reg967 = (~|{($unsigned((8'haf)) && $signed(reg935))});
                      reg968 <= (~^(~|$signed(((8'hb1) + reg825))));
                    end
                  else
                    begin
                      reg965 = ($signed(((reg746 ? reg945 : reg891) < reg917)) ?
                          ("" & forvar933[(3'h5):(3'h5)]) : (reg937 ?
                              $unsigned({reg754}) : $signed((reg677 ?
                                  reg814 : reg843))));
                      reg967 = $signed({reg883});
                      reg968 <= reg879[(4'hd):(4'h8)];
                      reg969 = $signed({(^reg897[(3'h7):(3'h4)])});
                    end
                  for (forvar970 = (1'h0); (forvar970 < (1'h1)); forvar970 = (forvar970 + (1'h1)))
                    begin
                      reg971 <= (reg711[(3'h6):(3'h4)] ?
                          (8'hb9) : ((~|(~reg850)) != (+reg815[(4'hb):(3'h5)])));
                    end
                  for (forvar972 = (1'h0); (forvar972 < (1'h0)); forvar972 = (forvar972 + (1'h1)))
                    begin
                      reg973 = ((((8'hab) ?
                              (~|reg883) : $signed((8'hac))) ^ (wire655 ?
                              $signed(reg686) : $signed(reg876))) ?
                          $unsigned({forvar853[(2'h3):(2'h3)]}) : ((&(reg964 & forvar876)) >> ({reg896} ?
                              (~|reg849) : (reg904 >= (8'h9e)))));
                      reg974 = "2zhhd";
                    end
                end
            end
          reg975 = $signed(reg678);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module624  (y, clk, wire629, wire628, wire627, wire626, wire625);
  output wire [(32'h85):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire629;
  input wire signed [(4'ha):(1'h0)] wire628;
  input wire [(4'hc):(1'h0)] wire627;
  input wire [(4'he):(1'h0)] wire626;
  input wire signed [(3'h7):(1'h0)] wire625;
  wire signed [(4'he):(1'h0)] wire644;
  wire signed [(4'hc):(1'h0)] wire633;
  wire [(4'hc):(1'h0)] wire632;
  wire signed [(2'h2):(1'h0)] wire631;
  wire [(4'ha):(1'h0)] wire630;
  reg signed [(2'h3):(1'h0)] reg641 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg638 = (1'h0);
  reg [(3'h6):(1'h0)] reg635 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg639 = (1'h0);
  reg [(4'hb):(1'h0)] reg643 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg642 = (1'h0);
  reg [(4'hf):(1'h0)] reg640 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar639 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar637 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg636 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar634 = (1'h0);
  assign y = {wire631, reg641, reg638, reg636, (1'h0)};
  assign wire630 = $unsigned((^{(wire626 && wire626)}));
  assign wire631 = (wire627[(4'hc):(3'h5)] ?
                       $signed((&$signed(wire625))) : (wire630 == (+$unsigned((8'ha8)))));
  assign wire632 = $unsigned(wire625);
  assign wire633 = $signed(wire626[(4'h9):(4'h8)]);
  always
    @(posedge clk) begin
      for (forvar634 = (1'h0); (forvar634 < (1'h1)); forvar634 = (forvar634 + (1'h1)))
        begin
          reg635 <= (-wire628);
          reg636 = wire625[(2'h3):(1'h0)];
          for (forvar637 = (1'h0); (forvar637 < (2'h3)); forvar637 = (forvar637 + (1'h1)))
            begin
              reg638 <= $unsigned((+("vNNWaCldSLVFNJ" > "DMcn")));
              if ($signed((($signed(reg635) * "V0") >> forvar637)))
                begin
                  for (forvar639 = (1'h0); (forvar639 < (2'h3)); forvar639 = (forvar639 + (1'h1)))
                    begin
                      reg640 = (|$signed({(~&wire630)}));
                      reg641 <= "GDfummRHCH3JS3f";
                    end
                  reg642 = {wire629[(4'h8):(3'h6)]};
                  reg643 = wire633[(4'hc):(1'h0)];
                end
              else
                begin
                  reg639 = wire630[(3'h7):(2'h3)];
                  reg640 = wire626;
                end
            end
        end
    end
  assign wire644 = ($signed(wire626[(3'h7):(2'h3)]) | {$unsigned($signed(wire633))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1291
#(parameter param1848 = (8'ha6))
(y, clk, wire1292, wire1293, wire1294, wire1295, wire1296);
  output wire [(32'hccc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire1292;
  input wire signed [(2'h3):(1'h0)] wire1293;
  input wire signed [(4'hb):(1'h0)] wire1294;
  input wire [(4'hf):(1'h0)] wire1295;
  input wire signed [(3'h5):(1'h0)] wire1296;
  wire signed [(4'h8):(1'h0)] wire1847;
  wire signed [(3'h4):(1'h0)] wire1663;
  wire signed [(4'hb):(1'h0)] wire1556;
  wire [(3'h4):(1'h0)] wire1297;
  wire [(4'hb):(1'h0)] wire1298;
  wire signed [(3'h5):(1'h0)] wire1299;
  wire signed [(3'h7):(1'h0)] wire1538;
  reg signed [(3'h7):(1'h0)] reg1846 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1842 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1833 = (1'h0);
  reg [(3'h5):(1'h0)] reg1831 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1829 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1827 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1826 = (1'h0);
  reg [(4'he):(1'h0)] reg1820 = (1'h0);
  reg [(4'h8):(1'h0)] reg1812 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1796 = (1'h0);
  reg [(2'h3):(1'h0)] reg1817 = (1'h0);
  reg [(5'h10):(1'h0)] reg1813 = (1'h0);
  reg [(3'h4):(1'h0)] reg1807 = (1'h0);
  reg [(4'ha):(1'h0)] reg1806 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1805 = (1'h0);
  reg [(4'hc):(1'h0)] reg1801 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1803 = (1'h0);
  reg [(4'h9):(1'h0)] reg1802 = (1'h0);
  reg [(4'hf):(1'h0)] reg1721 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1790 = (1'h0);
  reg [(4'h9):(1'h0)] reg1783 = (1'h0);
  reg [(4'hd):(1'h0)] reg1780 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1779 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1773 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1771 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1767 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1763 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1759 = (1'h0);
  reg [(4'hd):(1'h0)] reg1752 = (1'h0);
  reg [(3'h6):(1'h0)] reg1747 = (1'h0);
  reg [(5'h10):(1'h0)] reg1745 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1743 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1734 = (1'h0);
  reg [(4'hf):(1'h0)] reg1729 = (1'h0);
  reg [(4'hd):(1'h0)] reg1728 = (1'h0);
  reg [(2'h2):(1'h0)] reg1726 = (1'h0);
  reg [(4'hd):(1'h0)] reg1725 = (1'h0);
  reg [(3'h7):(1'h0)] reg1724 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1722 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1716 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1708 = (1'h0);
  reg [(4'hc):(1'h0)] reg1703 = (1'h0);
  reg [(2'h3):(1'h0)] reg1701 = (1'h0);
  reg [(3'h5):(1'h0)] reg1697 = (1'h0);
  reg [(4'h8):(1'h0)] reg1694 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1689 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1685 = (1'h0);
  reg [(3'h4):(1'h0)] reg1682 = (1'h0);
  reg [(4'he):(1'h0)] reg1680 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1677 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1673 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1668 = (1'h0);
  reg [(4'hf):(1'h0)] reg1661 = (1'h0);
  reg [(4'ha):(1'h0)] reg1657 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1649 = (1'h0);
  reg [(4'hf):(1'h0)] reg1636 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1645 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1643 = (1'h0);
  reg [(3'h4):(1'h0)] reg1641 = (1'h0);
  reg [(3'h6):(1'h0)] reg1639 = (1'h0);
  reg [(3'h5):(1'h0)] reg1638 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1633 = (1'h0);
  reg [(2'h2):(1'h0)] reg1632 = (1'h0);
  reg [(4'hb):(1'h0)] reg1619 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1614 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1628 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1626 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1625 = (1'h0);
  reg [(2'h3):(1'h0)] reg1623 = (1'h0);
  reg [(4'h9):(1'h0)] reg1608 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1597 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1595 = (1'h0);
  reg [(4'hf):(1'h0)] reg1594 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1589 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1586 = (1'h0);
  reg [(2'h2):(1'h0)] reg1584 = (1'h0);
  reg [(3'h7):(1'h0)] reg1583 = (1'h0);
  reg [(4'hc):(1'h0)] reg1580 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1575 = (1'h0);
  reg [(4'hc):(1'h0)] reg1574 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1572 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1571 = (1'h0);
  reg [(3'h5):(1'h0)] reg1570 = (1'h0);
  reg [(4'ha):(1'h0)] reg1569 = (1'h0);
  reg [(2'h3):(1'h0)] reg1566 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1564 = (1'h0);
  reg [(4'hf):(1'h0)] reg1563 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1560 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1548 = (1'h0);
  reg [(4'he):(1'h0)] reg1555 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1553 = (1'h0);
  reg [(4'hf):(1'h0)] reg1552 = (1'h0);
  reg [(4'hb):(1'h0)] reg1550 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1545 = (1'h0);
  reg [(3'h6):(1'h0)] reg1543 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1821 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1819 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1798 = (1'h0);
  reg [(3'h7):(1'h0)] reg1845 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1844 = (1'h0);
  reg [(2'h2):(1'h0)] reg1843 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1841 = (1'h0);
  reg [(4'hb):(1'h0)] reg1840 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1839 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1838 = (1'h0);
  reg [(4'hf):(1'h0)] reg1837 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1836 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1835 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1834 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1832 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1829 = (1'h0);
  reg [(4'hd):(1'h0)] reg1830 = (1'h0);
  reg [(3'h5):(1'h0)] reg1828 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1825 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1824 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1823 = (1'h0);
  reg [(4'he):(1'h0)] reg1822 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1821 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1819 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1815 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1810 = (1'h0);
  reg [(2'h3):(1'h0)] reg1809 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1808 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1802 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1818 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1814 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1816 = (1'h0);
  reg [(3'h6):(1'h0)] reg1815 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1814 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1812 = (1'h0);
  reg [(3'h5):(1'h0)] reg1811 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1810 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1809 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1808 = (1'h0);
  reg [(4'hc):(1'h0)] reg1804 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1801 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1800 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1799 = (1'h0);
  reg [(3'h7):(1'h0)] reg1798 = (1'h0);
  reg [(4'h9):(1'h0)] reg1797 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1796 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1795 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1722 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1794 = (1'h0);
  reg [(3'h4):(1'h0)] reg1793 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1792 = (1'h0);
  reg [(3'h7):(1'h0)] reg1791 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1789 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1788 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1787 = (1'h0);
  reg [(3'h7):(1'h0)] reg1786 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1785 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1784 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1781 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1784 = (1'h0);
  reg [(4'hf):(1'h0)] reg1782 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1781 = (1'h0);
  reg [(4'hc):(1'h0)] reg1778 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1777 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1776 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1775 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1774 = (1'h0);
  reg [(3'h4):(1'h0)] reg1772 = (1'h0);
  reg [(4'hd):(1'h0)] reg1770 = (1'h0);
  reg [(3'h6):(1'h0)] reg1769 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1768 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1766 = (1'h0);
  reg [(3'h4):(1'h0)] reg1765 = (1'h0);
  reg [(4'he):(1'h0)] forvar1764 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1762 = (1'h0);
  reg [(3'h7):(1'h0)] reg1761 = (1'h0);
  reg [(2'h2):(1'h0)] reg1760 = (1'h0);
  reg [(5'h10):(1'h0)] reg1758 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1757 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1756 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1755 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1754 = (1'h0);
  reg [(3'h5):(1'h0)] reg1753 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1751 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1750 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1749 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1748 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1746 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1744 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1742 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1741 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1740 = (1'h0);
  reg [(4'h9):(1'h0)] reg1739 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1738 = (1'h0);
  reg [(3'h5):(1'h0)] reg1737 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1736 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1735 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1733 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1733 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1723 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1732 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1731 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1730 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1727 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1723 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1721 = (1'h0);
  reg [(2'h2):(1'h0)] reg1720 = (1'h0);
  reg [(4'ha):(1'h0)] reg1713 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1719 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1718 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1717 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1716 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1715 = (1'h0);
  reg [(4'ha):(1'h0)] reg1714 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1713 = (1'h0);
  reg [(3'h5):(1'h0)] reg1712 = (1'h0);
  reg [(3'h4):(1'h0)] reg1711 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1710 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1709 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1707 = (1'h0);
  reg [(4'h8):(1'h0)] reg1706 = (1'h0);
  reg [(3'h5):(1'h0)] reg1705 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1704 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1702 = (1'h0);
  reg [(4'hf):(1'h0)] reg1700 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1699 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1698 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1696 = (1'h0);
  reg [(2'h3):(1'h0)] reg1695 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1693 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1692 = (1'h0);
  reg [(3'h7):(1'h0)] reg1691 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1690 = (1'h0);
  reg [(3'h4):(1'h0)] reg1688 = (1'h0);
  reg [(4'h8):(1'h0)] reg1687 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1686 = (1'h0);
  reg [(4'he):(1'h0)] reg1684 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1683 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1681 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1679 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1678 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1676 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1675 = (1'h0);
  reg [(4'ha):(1'h0)] reg1674 = (1'h0);
  reg [(2'h3):(1'h0)] reg1672 = (1'h0);
  reg [(3'h5):(1'h0)] reg1671 = (1'h0);
  reg [(4'h9):(1'h0)] reg1670 = (1'h0);
  reg [(5'h10):(1'h0)] reg1669 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1667 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1666 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1665 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1664 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1662 = (1'h0);
  reg [(3'h6):(1'h0)] reg1656 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1660 = (1'h0);
  reg [(3'h6):(1'h0)] reg1659 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1658 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1656 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1655 = (1'h0);
  reg [(2'h2):(1'h0)] reg1654 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1653 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1652 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1651 = (1'h0);
  reg [(5'h10):(1'h0)] reg1650 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1648 = (1'h0);
  reg [(4'h9):(1'h0)] reg1647 = (1'h0);
  reg [(3'h6):(1'h0)] reg1646 = (1'h0);
  reg [(4'ha):(1'h0)] reg1644 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1642 = (1'h0);
  reg [(5'h10):(1'h0)] reg1640 = (1'h0);
  reg [(4'hf):(1'h0)] reg1637 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1636 = (1'h0);
  reg [(3'h5):(1'h0)] reg1635 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1634 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1625 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1624 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1620 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1617 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1616 = (1'h0);
  reg [(4'hd):(1'h0)] reg1611 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1610 = (1'h0);
  reg [(4'hc):(1'h0)] reg1631 = (1'h0);
  reg [(4'h8):(1'h0)] reg1630 = (1'h0);
  reg [(4'hc):(1'h0)] reg1629 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1627 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1624 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1622 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1621 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1620 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1619 = (1'h0);
  reg [(4'hb):(1'h0)] reg1618 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1617 = (1'h0);
  reg [(4'hf):(1'h0)] reg1616 = (1'h0);
  reg [(4'hc):(1'h0)] reg1615 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1614 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1613 = (1'h0);
  reg [(4'hf):(1'h0)] reg1612 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1611 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1610 = (1'h0);
  reg [(3'h6):(1'h0)] reg1609 = (1'h0);
  reg [(3'h7):(1'h0)] reg1607 = (1'h0);
  reg [(4'h9):(1'h0)] reg1606 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1605 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1604 = (1'h0);
  reg [(4'ha):(1'h0)] reg1603 = (1'h0);
  reg [(4'ha):(1'h0)] reg1602 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1601 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1600 = (1'h0);
  reg [(4'hd):(1'h0)] reg1599 = (1'h0);
  reg [(3'h7):(1'h0)] reg1588 = (1'h0);
  reg [(4'hc):(1'h0)] reg1598 = (1'h0);
  reg [(5'h10):(1'h0)] reg1596 = (1'h0);
  reg [(3'h5):(1'h0)] reg1593 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1592 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1591 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1590 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1588 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1587 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1585 = (1'h0);
  reg [(3'h5):(1'h0)] reg1582 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1581 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1574 = (1'h0);
  reg [(4'he):(1'h0)] reg1573 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1568 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1562 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1558 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1581 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1580 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1577 = (1'h0);
  reg [(4'he):(1'h0)] forvar1576 = (1'h0);
  reg [(2'h2):(1'h0)] reg1579 = (1'h0);
  reg [(4'hc):(1'h0)] reg1578 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1577 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1576 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1573 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1568 = (1'h0);
  reg [(4'hb):(1'h0)] reg1567 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1565 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1559 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1557 = (1'h0);
  reg [(3'h6):(1'h0)] reg1565 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1562 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1561 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1559 = (1'h0);
  reg [(5'h10):(1'h0)] reg1558 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1557 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1546 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1542 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1554 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1552 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1551 = (1'h0);
  reg [(3'h4):(1'h0)] reg1549 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1548 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1547 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1546 = (1'h0);
  reg [(4'he):(1'h0)] reg1544 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1542 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1541 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1540 = (1'h0);
  assign y = {wire1556,
                 wire1298,
                 reg1842,
                 reg1833,
                 reg1827,
                 reg1812,
                 reg1796,
                 reg1817,
                 reg1813,
                 reg1807,
                 reg1801,
                 reg1721,
                 reg1790,
                 reg1783,
                 reg1780,
                 reg1752,
                 reg1745,
                 reg1728,
                 reg1722,
                 reg1716,
                 reg1708,
                 reg1703,
                 reg1689,
                 reg1668,
                 reg1649,
                 reg1636,
                 reg1643,
                 reg1639,
                 reg1595,
                 reg1586,
                 reg1584,
                 reg1572,
                 reg1569,
                 reg1552,
                 reg1821,
                 forvar1819,
                 forvar1798,
                 reg1843,
                 forvar1839,
                 reg1837,
                 reg1836,
                 forvar1835,
                 forvar1829,
                 forvar1825,
                 reg1819,
                 forvar1815,
                 reg1809,
                 forvar1809,
                 reg1804,
                 forvar1796,
                 reg1795,
                 forvar1722,
                 forvar1792,
                 reg1791,
                 forvar1787,
                 forvar1781,
                 forvar1776,
                 reg1772,
                 reg1757,
                 reg1754,
                 forvar1748,
                 reg1744,
                 reg1742,
                 reg1739,
                 forvar1733,
                 reg1730,
                 forvar1721,
                 reg1715,
                 forvar1713,
                 reg1709,
                 forvar1707,
                 reg1705,
                 forvar1699,
                 reg1688,
                 forvar1686,
                 reg1678,
                 reg1676,
                 reg1674,
                 reg1672,
                 forvar1665,
                 reg1664,
                 reg1662,
                 reg1658,
                 forvar1656,
                 reg1652,
                 forvar1651,
                 forvar1648,
                 reg1647,
                 reg1646,
                 reg1644,
                 forvar1636,
                 reg1635,
                 reg1617,
                 reg1630,
                 forvar1624,
                 reg1621,
                 reg1618,
                 reg1616,
                 reg1615,
                 reg1613,
                 reg1612,
                 reg1604,
                 forvar1601,
                 reg1599,
                 reg1588,
                 reg1598,
                 reg1596,
                 forvar1590,
                 reg1585,
                 forvar1581,
                 forvar1562,
                 forvar1558,
                 reg1581,
                 forvar1577,
                 reg1576,
                 forvar1568,
                 forvar1559,
                 reg1557,
                 reg1565,
                 reg1562,
                 reg1559,
                 forvar1552,
                 forvar1548,
                 forvar1541,
                 forvar1540,
                 (1'h0)};
  assign wire1297 = $unsigned($signed(({wire1295} ?
                        (&wire1293) : (wire1292 ? wire1295 : wire1292))));
  assign wire1298 = wire1293[(2'h2):(1'h0)];
  assign wire1299 = "45JbidzwaItFQ";
  module1300 #() modinst1539 (.wire1302(wire1292), .y(wire1538), .wire1304(wire1295), .wire1303(wire1298), .wire1305(wire1299), .wire1301(wire1296), .clk(clk));
  always
    @(posedge clk) begin
      for (forvar1540 = (1'h0); (forvar1540 < (2'h3)); forvar1540 = (forvar1540 + (1'h1)))
        begin
          if ($unsigned(wire1538[(1'h1):(1'h0)]))
            begin
              for (forvar1541 = (1'h0); (forvar1541 < (2'h3)); forvar1541 = (forvar1541 + (1'h1)))
                begin
                  if (($unsigned(((|wire1538) ?
                      $unsigned(wire1292) : $unsigned(wire1299))) * wire1292[(4'hd):(4'hd)]))
                    begin
                      reg1542 = wire1294[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg1543 <= "ImUoFLKx0wl";
                      reg1544 = "sy";
                      reg1545 <= wire1538[(2'h2):(1'h1)];
                      reg1546 = (-{((wire1297 ?
                              (8'ha3) : wire1299) * forvar1541)});
                    end
                  reg1547 = (-$unsigned(($signed(forvar1541) ?
                      $signed(wire1295) : $signed(wire1297))));
                  for (forvar1548 = (1'h0); (forvar1548 < (1'h1)); forvar1548 = (forvar1548 + (1'h1)))
                    begin
                      reg1549 = (^((~^((8'ha2) - reg1547)) ?
                          ($signed(reg1543) <= $signed(reg1545)) : wire1298[(3'h5):(2'h2)]));
                    end
                end
              if (wire1292[(4'hc):(2'h3)])
                begin
                  reg1550 <= forvar1548;
                  reg1551 = reg1549[(2'h3):(2'h3)];
                  reg1552 <= $signed("r3");
                end
              else
                begin
                  reg1550 <= (~^wire1298[(3'h6):(1'h1)]);
                  reg1551 = "xe5TifRAIEU";
                  for (forvar1552 = (1'h0); (forvar1552 < (1'h1)); forvar1552 = (forvar1552 + (1'h1)))
                    begin
                      reg1553 <= reg1550[(3'h5):(1'h1)];
                      reg1554 = forvar1540[(2'h3):(2'h2)];
                    end
                end
              reg1555 <= "GYXEFs6";
            end
          else
            begin
              for (forvar1541 = (1'h0); (forvar1541 < (2'h3)); forvar1541 = (forvar1541 + (1'h1)))
                begin
                  for (forvar1542 = (1'h0); (forvar1542 < (2'h3)); forvar1542 = (forvar1542 + (1'h1)))
                    begin
                      reg1543 <= $unsigned(wire1292[(4'hd):(3'h7)]);
                      reg1544 = (($unsigned((~&reg1552)) ?
                              reg1543[(3'h4):(2'h2)] : (8'ha3)) ?
                          (^(-$signed(reg1543))) : (^~(|((8'ha5) ?
                              wire1293 : reg1547))));
                    end
                  reg1545 <= reg1550;
                  for (forvar1546 = (1'h0); (forvar1546 < (2'h3)); forvar1546 = (forvar1546 + (1'h1)))
                    begin
                      reg1548 <= (^~{{{forvar1546}}});
                      reg1550 <= (~reg1549);
                    end
                  reg1551 = (8'hb0);
                end
              reg1552 <= $signed((!(-(reg1542 ? wire1298 : reg1549))));
            end
        end
    end
  assign wire1556 = (^~wire1295);
  always
    @(posedge clk) begin
      if ($unsigned((wire1298 ^ (^~"w5yTuECBxBa7RyO"))))
        begin
          if (((reg1552[(4'he):(4'hb)] ?
              $unsigned((~&wire1293)) : (-$unsigned(wire1297))) <= (~$signed((reg1543 <= wire1293)))))
            begin
              for (forvar1557 = (1'h0); (forvar1557 < (2'h3)); forvar1557 = (forvar1557 + (1'h1)))
                begin
                  if (($signed($signed($signed(wire1295))) <<< wire1292[(3'h6):(3'h5)]))
                    begin
                      reg1558 = $unsigned($signed(reg1555[(4'h8):(3'h5)]));
                      reg1559 = wire1556;
                      reg1560 <= (wire1296 ?
                          ($unsigned(wire1556) > {(reg1543 ?
                                  reg1548 : reg1553)}) : $signed(wire1297[(2'h2):(1'h0)]));
                      reg1561 = ($signed(((&(8'ha4)) < (!reg1560))) ?
                          ($signed((8'ha6)) < (wire1292[(4'hf):(4'hf)] ?
                              $signed(wire1299) : {wire1294})) : $unsigned((~(reg1560 ?
                              wire1296 : wire1292))));
                    end
                  else
                    begin
                      reg1558 = (^~$unsigned($signed((wire1556 ?
                          wire1297 : wire1556))));
                      reg1559 = $unsigned((reg1555[(4'h8):(3'h6)] ?
                          (reg1543[(3'h5):(2'h2)] > reg1560[(4'h9):(1'h0)]) : reg1555));
                    end
                  if ((|reg1552[(3'h7):(3'h6)]))
                    begin
                      reg1562 = $unsigned((~|$signed(wire1295[(3'h7):(2'h3)])));
                    end
                  else
                    begin
                      reg1563 <= $unsigned(wire1556[(4'h9):(4'h8)]);
                    end
                  reg1564 <= $signed($unsigned("TmkpfFMhihWgzPi"));
                  reg1565 = (~reg1559);
                end
              reg1566 <= (reg1560 ?
                  wire1297[(2'h3):(1'h0)] : ($signed({wire1297}) || {$signed(wire1292)}));
            end
          else
            begin
              if ($signed(wire1556))
                begin
                  reg1557 = reg1561[(2'h3):(1'h0)];
                end
              else
                begin
                  if ({(reg1550 << "26nKZ")})
                    begin
                      reg1557 = forvar1557;
                      reg1558 = (!wire1556);
                    end
                  else
                    begin
                      reg1557 = (^(reg1555[(1'h1):(1'h1)] || $signed(reg1550[(2'h2):(1'h0)])));
                      reg1558 = "8ICk2KXwX";
                    end
                  for (forvar1559 = (1'h0); (forvar1559 < (2'h2)); forvar1559 = (forvar1559 + (1'h1)))
                    begin
                      reg1560 <= wire1294[(4'ha):(1'h1)];
                      reg1561 = (~^$signed(((^wire1297) ?
                          {reg1553} : $signed(forvar1557))));
                      reg1563 <= $unsigned("5");
                      reg1564 <= $unsigned(($signed(((8'hb0) ?
                          reg1566 : (8'hb4))) >> "uPv1DoUk1R3h3nC"));
                    end
                end
              for (forvar1565 = (1'h0); (forvar1565 < (1'h1)); forvar1565 = (forvar1565 + (1'h1)))
                begin
                  reg1567 = wire1295[(4'hc):(4'hc)];
                  for (forvar1568 = (1'h0); (forvar1568 < (1'h1)); forvar1568 = (forvar1568 + (1'h1)))
                    begin
                      reg1569 <= "82Rrs";
                      reg1570 <= ($signed(($signed(reg1562) ?
                          reg1559[(1'h0):(1'h0)] : wire1556)) >= $signed($unsigned((&forvar1559))));
                      reg1571 <= ((&($signed(forvar1565) >= (-(8'ha1)))) ?
                          (forvar1568 ?
                              (^~reg1552[(4'hd):(3'h6)]) : "voE") : ({(reg1543 != reg1567)} ?
                              ((~&forvar1557) ?
                                  (reg1565 > reg1560) : {reg1543}) : (~&forvar1565)));
                      reg1572 <= (reg1561 ?
                          $unsigned((+"bfsTdAxf0iFccK3")) : (reg1567[(3'h5):(3'h4)] ?
                              (8'ha5) : ((wire1299 >= reg1565) ?
                                  $unsigned(wire1293) : ((8'haa) <<< reg1571))));
                    end
                  for (forvar1573 = (1'h0); (forvar1573 < (2'h3)); forvar1573 = (forvar1573 + (1'h1)))
                    begin
                      reg1574 <= ($unsigned("bTbfaILe") > wire1297[(3'h4):(2'h2)]);
                    end
                end
              reg1575 <= "fm7A5uXi7u";
              if (((!$unsigned("vva4CICL3WQS")) ?
                  ((-(~&reg1570)) ?
                      reg1560[(1'h1):(1'h1)] : ((~|reg1555) + {reg1565})) : ("T7QDvw" <<< (reg1548 ?
                      $signed(wire1298) : reg1572[(3'h5):(1'h1)]))))
                begin
                  reg1576 = wire1293[(1'h1):(1'h1)];
                  for (forvar1577 = (1'h0); (forvar1577 < (2'h3)); forvar1577 = (forvar1577 + (1'h1)))
                    begin
                      reg1578 = "fK";
                      reg1579 = {wire1292[(3'h6):(2'h2)]};
                    end
                  reg1580 <= {((+$signed(reg1553)) > ({reg1555} < {reg1550}))};
                end
              else
                begin
                  for (forvar1576 = (1'h0); (forvar1576 < (2'h3)); forvar1576 = (forvar1576 + (1'h1)))
                    begin
                      reg1577 = $unsigned($unsigned($signed(reg1545)));
                      reg1578 = (~^forvar1559[(3'h5):(1'h1)]);
                    end
                  reg1579 = "P7gMZmxo9JkPQ1Y";
                  for (forvar1580 = (1'h0); (forvar1580 < (1'h1)); forvar1580 = (forvar1580 + (1'h1)))
                    begin
                      reg1581 = $unsigned((~(((8'hac) <<< reg1569) ?
                          $unsigned(reg1560) : wire1556[(3'h5):(2'h3)])));
                    end
                end
            end
        end
      else
        begin
          if ((8'h9e))
            begin
              for (forvar1557 = (1'h0); (forvar1557 < (1'h1)); forvar1557 = (forvar1557 + (1'h1)))
                begin
                  for (forvar1558 = (1'h0); (forvar1558 < (2'h3)); forvar1558 = (forvar1558 + (1'h1)))
                    begin
                      reg1559 = {$signed($unsigned({reg1571}))};
                      reg1561 = $signed(("fFyMNvYc" ?
                          (forvar1573 | $signed(reg1562)) : reg1559[(1'h0):(1'h0)]));
                    end
                end
              for (forvar1562 = (1'h0); (forvar1562 < (2'h2)); forvar1562 = (forvar1562 + (1'h1)))
                begin
                  if ("niIsWKk")
                    begin
                      reg1563 <= (-("" ?
                          $unsigned((reg1550 ?
                              reg1577 : forvar1562)) : (|wire1299[(3'h4):(3'h4)])));
                      reg1565 = reg1550;
                    end
                  else
                    begin
                      reg1565 = $unsigned({("HkzPcsv6" != (reg1572 ?
                              reg1569 : reg1569))});
                      reg1567 = $unsigned((-reg1575));
                      reg1568 = ({$signed(reg1553[(1'h0):(1'h0)])} ?
                          ({reg1560} ? reg1581 : "O4z") : "DgOraxfeWuxApqu");
                      reg1573 = ((!({forvar1562} || (~^reg1569))) ?
                          $signed($unsigned($signed(wire1297))) : $signed(($unsigned(reg1553) ?
                              reg1577[(1'h0):(1'h0)] : wire1292[(1'h0):(1'h0)])));
                    end
                  for (forvar1574 = (1'h0); (forvar1574 < (1'h1)); forvar1574 = (forvar1574 + (1'h1)))
                    begin
                      reg1575 <= $signed((-reg1555[(3'h7):(3'h7)]));
                      reg1576 = $signed(((8'hba) > $unsigned(reg1570)));
                      reg1577 = (($unsigned(wire1556) ?
                              ((reg1578 ? reg1550 : reg1545) ?
                                  (reg1566 <= forvar1558) : $unsigned(reg1568)) : (reg1563[(3'h6):(3'h4)] >> {reg1576})) ?
                          $signed("GQV") : {$unsigned((wire1292 + reg1562))});
                      reg1580 <= $unsigned((-$unsigned((forvar1557 + reg1572))));
                    end
                  for (forvar1581 = (1'h0); (forvar1581 < (2'h3)); forvar1581 = (forvar1581 + (1'h1)))
                    begin
                      reg1582 = ("SIz7HAU7GeX" + $signed(("yo0g" <= $signed(reg1575))));
                      reg1583 <= $unsigned((~reg1577));
                      reg1584 <= $unsigned(forvar1562[(1'h1):(1'h0)]);
                    end
                end
              reg1585 = ("OOD3" ^ wire1294[(4'ha):(2'h3)]);
              reg1586 <= $signed($unsigned({$unsigned(reg1558)}));
            end
          else
            begin
              for (forvar1557 = (1'h0); (forvar1557 < (2'h3)); forvar1557 = (forvar1557 + (1'h1)))
                begin
                  for (forvar1558 = (1'h0); (forvar1558 < (1'h1)); forvar1558 = (forvar1558 + (1'h1)))
                    begin
                      reg1559 = "kn";
                      reg1561 = $signed(reg1550);
                      reg1562 = reg1582;
                    end
                  reg1565 = (~(^$unsigned($signed(forvar1557))));
                end
              reg1567 = (8'ha6);
            end
          for (forvar1587 = (1'h0); (forvar1587 < (2'h2)); forvar1587 = (forvar1587 + (1'h1)))
            begin
              if ((~^reg1561[(1'h1):(1'h0)]))
                begin
                  for (forvar1588 = (1'h0); (forvar1588 < (1'h1)); forvar1588 = (forvar1588 + (1'h1)))
                    begin
                      reg1589 <= $unsigned({$signed($unsigned((8'h9f)))});
                    end
                  for (forvar1590 = (1'h0); (forvar1590 < (1'h1)); forvar1590 = (forvar1590 + (1'h1)))
                    begin
                      reg1591 = reg1584;
                      reg1592 = forvar1587;
                      reg1593 = (|reg1550[(1'h0):(1'h0)]);
                      reg1594 <= $signed(reg1561);
                    end
                  if (((8'hb6) ?
                      (!$unsigned(reg1557[(2'h2):(2'h2)])) : (({reg1559} == $signed(reg1574)) || "P6b2eS")))
                    begin
                      reg1595 <= reg1576;
                      reg1596 = $signed(reg1577);
                    end
                  else
                    begin
                      reg1596 = $signed(reg1559[(3'h6):(3'h5)]);
                      reg1597 <= $unsigned(reg1578);
                      reg1598 = $unsigned(forvar1577);
                    end
                end
              else
                begin
                  reg1588 = (8'ha8);
                  reg1589 <= (~&"E27O");
                end
              reg1599 = "";
              for (forvar1600 = (1'h0); (forvar1600 < (1'h0)); forvar1600 = (forvar1600 + (1'h1)))
                begin
                  for (forvar1601 = (1'h0); (forvar1601 < (1'h0)); forvar1601 = (forvar1601 + (1'h1)))
                    begin
                      reg1602 = ($signed({(+reg1580)}) ?
                          forvar1562 : $unsigned(($signed(reg1561) <= {(8'ha2)})));
                      reg1603 = forvar1600;
                      reg1604 = (((~^forvar1558) && $unsigned($unsigned(reg1570))) - "");
                    end
                  for (forvar1605 = (1'h0); (forvar1605 < (2'h3)); forvar1605 = (forvar1605 + (1'h1)))
                    begin
                      reg1606 = reg1555;
                      reg1607 = $unsigned(({$signed(reg1561)} ?
                          $unsigned(reg1564[(3'h6):(3'h5)]) : (~^(+reg1586))));
                      reg1608 <= (|{reg1603});
                    end
                end
            end
          reg1609 = $signed($unsigned((^(reg1559 ? reg1581 : forvar1577))));
          if ($unsigned("wdVdEZd"))
            begin
              for (forvar1610 = (1'h0); (forvar1610 < (1'h1)); forvar1610 = (forvar1610 + (1'h1)))
                begin
                  for (forvar1611 = (1'h0); (forvar1611 < (2'h3)); forvar1611 = (forvar1611 + (1'h1)))
                    begin
                      reg1612 = $unsigned($signed(forvar1576));
                      reg1613 = $signed($signed({$signed(reg1603)}));
                    end
                  for (forvar1614 = (1'h0); (forvar1614 < (1'h1)); forvar1614 = (forvar1614 + (1'h1)))
                    begin
                      reg1615 = (-(!(^(~reg1576))));
                      reg1616 = "1Zs";
                    end
                end
              for (forvar1617 = (1'h0); (forvar1617 < (2'h3)); forvar1617 = (forvar1617 + (1'h1)))
                begin
                  reg1618 = forvar1574[(1'h0):(1'h0)];
                end
              for (forvar1619 = (1'h0); (forvar1619 < (2'h3)); forvar1619 = (forvar1619 + (1'h1)))
                begin
                  for (forvar1620 = (1'h0); (forvar1620 < (1'h1)); forvar1620 = (forvar1620 + (1'h1)))
                    begin
                      reg1621 = "1G";
                      reg1622 = $unsigned(({reg1577[(2'h2):(1'h1)]} * forvar1611[(4'hc):(2'h3)]));
                      reg1623 <= (-{(~&$signed(reg1604))});
                    end
                  for (forvar1624 = (1'h0); (forvar1624 < (1'h1)); forvar1624 = (forvar1624 + (1'h1)))
                    begin
                      reg1625 <= ("2O8WCVe9VZz" - $signed($unsigned(reg1567)));
                      reg1626 <= {((8'hb9) ?
                              $unsigned($signed(reg1592)) : ($signed((8'hb4)) ?
                                  {(8'h9e)} : (^~reg1545)))};
                    end
                  if ((((!$unsigned(forvar1587)) ?
                      $unsigned($unsigned(reg1584)) : $unsigned({reg1553})) || $signed(reg1608[(1'h0):(1'h0)])))
                    begin
                      reg1627 = reg1612[(4'hd):(3'h7)];
                    end
                  else
                    begin
                      reg1628 <= "qeUyDuw8wFZR";
                      reg1629 = $signed((forvar1565[(3'h6):(2'h3)] ?
                          ("PPt" ?
                              $unsigned((8'h9f)) : $unsigned(reg1564)) : $unsigned($unsigned(reg1586))));
                    end
                  reg1630 = (("OqgV" <= (&wire1556)) ?
                      (^~({forvar1573} ?
                          (reg1582 ?
                              reg1545 : reg1623) : reg1609[(3'h5):(1'h1)])) : $signed((~&reg1618[(3'h7):(3'h6)])));
                end
              reg1631 = ((^~$signed(reg1565)) ?
                  (reg1621 & ({reg1558} ~^ (reg1565 ?
                      forvar1617 : (8'ha3)))) : (+(8'ha2)));
            end
          else
            begin
              if (forvar1559)
                begin
                  if (reg1562)
                    begin
                      reg1610 = $signed((!$unsigned($signed((8'ha0)))));
                      reg1611 = (|"bFDSiQ8K3D");
                      reg1612 = (^(^~$signed($signed(reg1552))));
                    end
                  else
                    begin
                      reg1610 = (reg1557 ?
                          ((8'haf) ?
                              (+wire1295[(4'ha):(2'h3)]) : reg1626[(1'h0):(1'h0)]) : wire1295);
                      reg1611 = ("oOKDfqYEHDb7EUe" - ($signed({(8'ha9)}) * $signed($signed((8'hb9)))));
                      reg1614 <= $signed(reg1559);
                      reg1615 = reg1575[(1'h1):(1'h1)];
                    end
                  for (forvar1616 = (1'h0); (forvar1616 < (2'h3)); forvar1616 = (forvar1616 + (1'h1)))
                    begin
                      reg1617 = (!forvar1617[(5'h10):(4'hd)]);
                      reg1619 <= reg1577[(1'h0):(1'h0)];
                      reg1620 = ($signed("okEyeDMUx") ?
                          reg1618[(2'h2):(1'h0)] : forvar1568[(2'h3):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar1610 = (1'h0); (forvar1610 < (1'h0)); forvar1610 = (forvar1610 + (1'h1)))
                    begin
                      reg1614 <= $signed(((forvar1576[(1'h0):(1'h0)] ?
                          {reg1609} : forvar1562) - (~^"Yzi6XZPvAqQ9F98")));
                      reg1619 <= forvar1580;
                    end
                  for (forvar1620 = (1'h0); (forvar1620 < (2'h3)); forvar1620 = (forvar1620 + (1'h1)))
                    begin
                      reg1623 <= ({("iLeuDt" >> (-reg1612))} ^ (forvar1605 + forvar1588[(2'h2):(1'h1)]));
                      reg1624 = (forvar1617[(4'hd):(3'h5)] & wire1298);
                    end
                  for (forvar1625 = (1'h0); (forvar1625 < (1'h0)); forvar1625 = (forvar1625 + (1'h1)))
                    begin
                      reg1627 = $signed(($unsigned($unsigned((8'ha2))) & (+wire1293)));
                      reg1629 = $unsigned((reg1561[(1'h0):(1'h0)] ?
                          forvar1577[(1'h0):(1'h0)] : $signed($unsigned(reg1624))));
                    end
                  if ($unsigned("Hnifw7"))
                    begin
                      reg1632 <= "1MP8ZxwduwJ";
                      reg1633 <= ((~|(|(reg1578 ? reg1604 : reg1591))) ?
                          {reg1579[(1'h0):(1'h0)]} : ((reg1585[(1'h0):(1'h0)] == ((8'ha0) ?
                              wire1292 : reg1625)) || (((8'hb2) ?
                                  (8'had) : reg1552) ?
                              (&(8'h9c)) : reg1566)));
                      reg1634 = (-(-$signed(forvar1565)));
                      reg1635 = ({((reg1557 ?
                              forvar1590 : reg1621) <= ((8'hb2) ?
                              reg1550 : reg1555))} == {reg1591[(3'h4):(1'h1)]});
                    end
                  else
                    begin
                      reg1632 <= "wOIr6Wuioilzo6";
                      reg1633 <= "B0HXdVg5kfY";
                      reg1634 = (~&reg1626[(2'h2):(1'h0)]);
                      reg1635 = reg1575;
                    end
                end
              if ((($unsigned($signed(reg1595)) ?
                      $unsigned($unsigned(reg1577)) : reg1624) ?
                  $signed(((^~reg1597) ?
                      (reg1631 ?
                          reg1565 : (8'hba)) : $signed(reg1607))) : ({(reg1614 != reg1626)} < reg1557)))
                begin
                  for (forvar1636 = (1'h0); (forvar1636 < (2'h2)); forvar1636 = (forvar1636 + (1'h1)))
                    begin
                      reg1637 = (&(forvar1576[(3'h7):(3'h5)] >> $unsigned(reg1564[(2'h2):(2'h2)])));
                      reg1638 <= reg1604;
                      reg1639 <= $signed(($signed(reg1570) <= $signed((8'ha9))));
                    end
                  reg1640 = $unsigned(reg1585[(1'h0):(1'h0)]);
                  reg1641 <= {$signed($unsigned($unsigned(reg1629)))};
                  if (reg1620[(1'h0):(1'h0)])
                    begin
                      reg1642 = (({reg1588} ?
                              (~^(reg1596 ?
                                  wire1296 : reg1620)) : $signed(reg1578)) ?
                          $unsigned({{forvar1588}}) : reg1559);
                      reg1643 <= "UFCxgu";
                      reg1644 = $unsigned($signed($signed((reg1562 ?
                          reg1578 : forvar1619))));
                      reg1645 <= $unsigned({$unsigned(reg1622)});
                    end
                  else
                    begin
                      reg1642 = (^~($signed("YbEEe") > $unsigned($signed(reg1611))));
                    end
                end
              else
                begin
                  if (reg1619)
                    begin
                      reg1636 <= {({"Q3pxhkGilO"} ?
                              ($signed(forvar1562) != $unsigned(reg1645)) : ((reg1563 ?
                                  (8'h9f) : wire1292) ^~ reg1602))};
                      reg1637 = $signed(reg1571[(3'h7):(3'h7)]);
                      reg1640 = forvar1577[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1637 = $unsigned("GA13OUTwoso");
                      reg1640 = (+$signed(((reg1569 ?
                          reg1639 : reg1560) >> $signed((8'hb5)))));
                    end
                  if (reg1638[(3'h4):(3'h4)])
                    begin
                      reg1642 = $unsigned((((reg1543 ^ reg1575) > (&(8'haf))) ?
                          $unsigned($unsigned(reg1640)) : reg1568[(3'h4):(1'h0)]));
                      reg1643 <= {$unsigned((reg1576 ?
                              reg1580[(4'hc):(3'h6)] : reg1588[(3'h7):(3'h5)]))};
                      reg1645 <= ((((forvar1601 ? reg1627 : forvar1617) ?
                              $unsigned(reg1617) : reg1597) ~^ (reg1550 ?
                              $unsigned(wire1299) : forvar1574[(2'h3):(1'h0)])) ?
                          $unsigned($unsigned({(8'hb1)})) : wire1294);
                      reg1646 = reg1584[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1642 = (&(~$unsigned($signed(reg1561))));
                      reg1644 = "d0ZM4LZtrR";
                      reg1646 = reg1557;
                      reg1647 = (($unsigned((reg1586 ?
                          reg1593 : (8'haa))) >>> "WRv8wHWWyEL5s") * reg1573);
                    end
                  for (forvar1648 = (1'h0); (forvar1648 < (1'h1)); forvar1648 = (forvar1648 + (1'h1)))
                    begin
                      reg1649 <= reg1543;
                      reg1650 = $unsigned(("OsP56H3If0qVJ" & $signed((&reg1592))));
                    end
                  for (forvar1651 = (1'h0); (forvar1651 < (1'h1)); forvar1651 = (forvar1651 + (1'h1)))
                    begin
                      reg1652 = "XElciEqaRFcsO";
                      reg1653 = (~(reg1562 >> {(8'hab)}));
                      reg1654 = {$signed($unsigned(reg1653))};
                      reg1655 = reg1564[(4'h8):(4'h8)];
                    end
                end
              if ($signed(reg1567[(4'hb):(2'h3)]))
                begin
                  for (forvar1656 = (1'h0); (forvar1656 < (1'h0)); forvar1656 = (forvar1656 + (1'h1)))
                    begin
                      reg1657 <= (~|($signed(wire1556[(2'h2):(1'h0)]) & (|forvar1565)));
                      reg1658 = ($signed((forvar1573[(1'h1):(1'h1)] ?
                          (^wire1294) : reg1625)) <<< ($unsigned((reg1602 - reg1571)) ?
                          ($signed(reg1610) ?
                              (reg1569 ?
                                  forvar1590 : reg1607) : "RGWrmBJ68HEIRM") : "fYyykEKap"));
                    end
                  if (("fCHHIxq0o6M" > (~&(~{reg1641}))))
                    begin
                      reg1659 = $unsigned(reg1558);
                      reg1660 = (((^(reg1557 ^ forvar1590)) || reg1602[(3'h5):(3'h5)]) | (8'hba));
                    end
                  else
                    begin
                      reg1659 = ($unsigned((~$unsigned(reg1585))) < $unsigned((~forvar1574[(3'h6):(1'h0)])));
                      reg1661 <= $unsigned(($unsigned((!forvar1577)) ?
                          {$unsigned(reg1643)} : ((~^reg1658) != forvar1580[(1'h0):(1'h0)])));
                    end
                end
              else
                begin
                  if ((8'ha1))
                    begin
                      reg1656 = $signed("GLnI");
                      reg1657 <= {forvar1620[(1'h0):(1'h0)]};
                      reg1658 = reg1638[(1'h0):(1'h0)];
                      reg1659 = reg1613[(3'h7):(1'h1)];
                    end
                  else
                    begin
                      reg1656 = {(8'ha7)};
                    end
                end
            end
        end
      reg1662 = (reg1550 ?
          $signed((forvar1614[(4'hb):(3'h4)] >= reg1627[(3'h7):(3'h4)])) : (((reg1580 == reg1655) ?
                  (reg1611 ? wire1292 : reg1657) : reg1656[(1'h0):(1'h0)]) ?
              ($signed((8'hb4)) ?
                  $unsigned(reg1631) : {reg1564}) : ($signed(forvar1651) ?
                  (+(8'ha0)) : reg1560)));
    end
  assign wire1663 = (&"iGMHGrRFSn");
  always
    @(posedge clk) begin
      reg1664 = $unsigned(($unsigned((&reg1619)) + reg1633));
      for (forvar1665 = (1'h0); (forvar1665 < (1'h1)); forvar1665 = (forvar1665 + (1'h1)))
        begin
          for (forvar1666 = (1'h0); (forvar1666 < (1'h1)); forvar1666 = (forvar1666 + (1'h1)))
            begin
              for (forvar1667 = (1'h0); (forvar1667 < (1'h0)); forvar1667 = (forvar1667 + (1'h1)))
                begin
                  reg1668 <= (wire1298 ?
                      reg1628[(3'h6):(3'h4)] : ((reg1586[(2'h3):(2'h2)] >>> (+reg1564)) ?
                          ("sUWLY0ghiQvn4" && reg1643) : ((-reg1594) <= (reg1636 ?
                              (8'hab) : reg1543))));
                  if (($signed(reg1566) + ((reg1623 * {reg1555}) ?
                      "IPvPES8w" : ((reg1560 >>> reg1639) ?
                          (forvar1666 ? reg1664 : (8'ha7)) : (8'hb5)))))
                    begin
                      reg1669 = $unsigned((-reg1575[(3'h5):(2'h2)]));
                      reg1670 = $unsigned(reg1571[(4'h9):(4'h8)]);
                      reg1671 = "YRr9Dfd7XTcEz9W";
                      reg1672 = ({wire1556} <<< reg1569[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg1669 = reg1594[(2'h3):(2'h2)];
                      reg1673 <= (wire1299 * {reg1608[(3'h4):(2'h2)]});
                      reg1674 = wire1295;
                    end
                  for (forvar1675 = (1'h0); (forvar1675 < (1'h1)); forvar1675 = (forvar1675 + (1'h1)))
                    begin
                      reg1676 = $unsigned({(&(reg1625 == (8'hac)))});
                      reg1677 <= {(~|"p7ACqw0A5Wvs")};
                    end
                  reg1678 = reg1574;
                end
            end
          for (forvar1679 = (1'h0); (forvar1679 < (1'h0)); forvar1679 = (forvar1679 + (1'h1)))
            begin
              reg1680 <= (+$signed($signed((~&reg1560))));
              for (forvar1681 = (1'h0); (forvar1681 < (2'h3)); forvar1681 = (forvar1681 + (1'h1)))
                begin
                  if ($unsigned(reg1645[(2'h2):(2'h2)]))
                    begin
                      reg1682 <= ("RLnOD6" < (((-forvar1666) ?
                              (reg1574 ? wire1295 : wire1294) : (reg1641 ?
                                  reg1589 : reg1548)) ?
                          forvar1665 : $signed((reg1664 >> reg1649))));
                    end
                  else
                    begin
                      reg1683 = reg1677[(4'h8):(3'h6)];
                      reg1684 = "FlL8FU9GSPnV";
                      reg1685 <= "f7psra9HgJKR";
                    end
                end
            end
          for (forvar1686 = (1'h0); (forvar1686 < (2'h2)); forvar1686 = (forvar1686 + (1'h1)))
            begin
              reg1687 = (reg1643[(1'h1):(1'h1)] ?
                  {($signed(forvar1681) | (reg1676 ?
                          forvar1665 : reg1570))} : (~&{reg1641}));
              reg1688 = (~^"pwIY4Kv");
              reg1689 <= ($signed(((!reg1571) <<< $signed((8'ha5)))) != ($unsigned({reg1672}) ?
                  ($signed(wire1293) <= (~|reg1684)) : $signed("ZpP4vsIXYENyDqy")));
            end
          for (forvar1690 = (1'h0); (forvar1690 < (1'h0)); forvar1690 = (forvar1690 + (1'h1)))
            begin
              reg1691 = $unsigned({(reg1597 ?
                      (reg1608 && reg1673) : (reg1560 | reg1575))});
              for (forvar1692 = (1'h0); (forvar1692 < (2'h3)); forvar1692 = (forvar1692 + (1'h1)))
                begin
                  if (reg1673[(2'h2):(1'h0)])
                    begin
                      reg1693 = reg1555[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg1693 = (wire1538[(2'h3):(2'h2)] >= $signed(($signed(reg1657) > $signed(reg1678))));
                      reg1694 <= reg1564[(2'h3):(2'h3)];
                      reg1695 = "G72RShx8";
                    end
                  for (forvar1696 = (1'h0); (forvar1696 < (2'h2)); forvar1696 = (forvar1696 + (1'h1)))
                    begin
                      reg1697 <= (reg1575 >>> $unsigned($unsigned((~|(8'hb3)))));
                    end
                end
              for (forvar1698 = (1'h0); (forvar1698 < (1'h1)); forvar1698 = (forvar1698 + (1'h1)))
                begin
                  for (forvar1699 = (1'h0); (forvar1699 < (1'h0)); forvar1699 = (forvar1699 + (1'h1)))
                    begin
                      reg1700 = (((~reg1580) > (reg1584[(1'h1):(1'h1)] || (reg1550 - (8'haa)))) ^~ (8'h9f));
                      reg1701 <= (reg1670[(3'h4):(2'h2)] >= "Y3a0XtT0YF");
                      reg1702 = ($unsigned(reg1701) < (8'ha6));
                    end
                  if (reg1633[(1'h1):(1'h0)])
                    begin
                      reg1703 <= $signed(("PTQzIFXvp6L0db" ?
                          ((reg1645 ?
                              reg1694 : reg1574) > forvar1690[(1'h1):(1'h0)]) : "o0nmeZdV"));
                      reg1704 = {(&($signed(reg1614) ?
                              $signed(reg1575) : (^~reg1619)))};
                      reg1705 = ((^$signed((reg1583 ^ reg1682))) ?
                          $signed(forvar1679) : (wire1292[(4'hb):(3'h5)] ?
                              {$signed(forvar1665)} : reg1676[(1'h0):(1'h0)]));
                      reg1706 = ($signed(forvar1666[(1'h1):(1'h0)]) || ($signed($signed(forvar1665)) <<< (^~(~^reg1580))));
                    end
                  else
                    begin
                      reg1704 = reg1695;
                      reg1705 = (&reg1626[(1'h0):(1'h0)]);
                    end
                  for (forvar1707 = (1'h0); (forvar1707 < (2'h3)); forvar1707 = (forvar1707 + (1'h1)))
                    begin
                      reg1708 <= reg1672[(1'h1):(1'h0)];
                      reg1709 = reg1608;
                      reg1710 = $unsigned(((^(~^(8'hb7))) + {(wire1296 >= reg1560)}));
                      reg1711 = $unsigned(reg1632);
                    end
                  reg1712 = reg1693[(1'h0):(1'h0)];
                end
              if (reg1623)
                begin
                  for (forvar1713 = (1'h0); (forvar1713 < (1'h0)); forvar1713 = (forvar1713 + (1'h1)))
                    begin
                      reg1714 = ($unsigned(($unsigned(reg1597) || (forvar1675 >> reg1626))) >>> $unsigned(((reg1682 >> reg1705) ?
                          "tByGXT4sev" : (wire1663 ? reg1688 : (8'hba)))));
                      reg1715 = $unsigned((&(+forvar1692[(1'h0):(1'h0)])));
                    end
                  for (forvar1716 = (1'h0); (forvar1716 < (2'h3)); forvar1716 = (forvar1716 + (1'h1)))
                    begin
                      reg1717 = "5bcplbd3RY";
                    end
                  for (forvar1718 = (1'h0); (forvar1718 < (2'h3)); forvar1718 = (forvar1718 + (1'h1)))
                    begin
                      reg1719 = (reg1677[(1'h1):(1'h0)] ?
                          $signed({(reg1715 ?
                                  reg1614 : reg1572)}) : (!(^~$unsigned(forvar1690))));
                    end
                end
              else
                begin
                  reg1713 = ($signed((|reg1709[(2'h2):(1'h0)])) ?
                      reg1673[(3'h4):(2'h2)] : {reg1580[(3'h4):(3'h4)]});
                  reg1714 = $signed(((-$unsigned(reg1608)) ?
                      ({reg1628} ?
                          (reg1697 << (8'hb1)) : $unsigned(reg1682)) : $unsigned((reg1545 >>> (8'ha0)))));
                  if ($signed($signed($signed((~forvar1679)))))
                    begin
                      reg1715 = $signed((wire1292[(3'h5):(3'h4)] <= reg1641));
                    end
                  else
                    begin
                      reg1715 = ($signed($signed(reg1713)) ?
                          wire1293[(1'h1):(1'h1)] : "eblAW");
                      reg1716 <= (~^$signed(reg1669[(4'h9):(2'h3)]));
                    end
                end
            end
        end
      if (reg1548)
        begin
          reg1720 = {$signed(((+reg1569) - reg1563[(4'hd):(3'h6)]))};
          for (forvar1721 = (1'h0); (forvar1721 < (2'h3)); forvar1721 = (forvar1721 + (1'h1)))
            begin
              reg1722 <= reg1643;
              if ($unsigned(forvar1686[(4'h8):(2'h3)]))
                begin
                  for (forvar1723 = (1'h0); (forvar1723 < (2'h2)); forvar1723 = (forvar1723 + (1'h1)))
                    begin
                      reg1724 <= (~$unsigned($signed($unsigned(reg1710))));
                      reg1725 <= $unsigned(("a5VE" ^ "X3MlGX"));
                    end
                  if (reg1626)
                    begin
                      reg1726 <= $unsigned("CSFhn9");
                      reg1727 = $signed($unsigned({"gx"}));
                      reg1728 <= (!reg1657);
                      reg1729 <= "M";
                    end
                  else
                    begin
                      reg1727 = $unsigned((^~{(reg1625 >> reg1716)}));
                      reg1730 = $signed(reg1726);
                      reg1731 = ($signed("Y") <= reg1548[(3'h4):(1'h0)]);
                    end
                  reg1732 = $unsigned(reg1708[(4'hb):(1'h0)]);
                end
              else
                begin
                  reg1723 = (~^$unsigned(reg1687[(1'h1):(1'h1)]));
                  if ((8'ha1))
                    begin
                      reg1727 = reg1583[(2'h2):(1'h1)];
                      reg1730 = ((wire1538[(3'h6):(1'h1)] ?
                          forvar1690 : reg1674) * reg1703);
                      reg1731 = (+$unsigned("mVZi"));
                    end
                  else
                    begin
                      reg1724 <= reg1682[(1'h1):(1'h0)];
                      reg1727 = $signed($signed($signed(((8'hb3) ?
                          forvar1692 : reg1726))));
                      reg1730 = (forvar1721 ?
                          "CJB7hfG" : (reg1580[(3'h7):(3'h7)] ?
                              wire1556 : {reg1710}));
                    end
                end
              if (reg1555[(1'h1):(1'h1)])
                begin
                  reg1733 = reg1710[(1'h1):(1'h1)];
                end
              else
                begin
                  for (forvar1733 = (1'h0); (forvar1733 < (2'h2)); forvar1733 = (forvar1733 + (1'h1)))
                    begin
                      reg1734 <= (reg1614 >>> $unsigned("x"));
                      reg1735 = (~(~&{(~&(8'h9f))}));
                      reg1736 = (&($signed($unsigned(reg1682)) ?
                          ($signed(reg1705) ?
                              reg1614[(2'h3):(2'h2)] : (!reg1545)) : (~^(+forvar1690))));
                      reg1737 = $unsigned(("ZK8ixP0Lpr6T0" && (~^(~|reg1566))));
                    end
                  for (forvar1738 = (1'h0); (forvar1738 < (1'h0)); forvar1738 = (forvar1738 + (1'h1)))
                    begin
                      reg1739 = (reg1552 ^~ (reg1574 ?
                          reg1545 : ({forvar1738} >= $signed(reg1669))));
                    end
                end
              for (forvar1740 = (1'h0); (forvar1740 < (2'h3)); forvar1740 = (forvar1740 + (1'h1)))
                begin
                  if ($unsigned(reg1680))
                    begin
                      reg1741 = forvar1707[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg1741 = "A6mT";
                      reg1742 = "nSqzwI";
                      reg1743 <= forvar1707[(1'h0):(1'h0)];
                      reg1744 = {"d3wXQUNRI"};
                    end
                  reg1745 <= $signed((-{((8'h9f) ~^ (8'ha4))}));
                  for (forvar1746 = (1'h0); (forvar1746 < (2'h2)); forvar1746 = (forvar1746 + (1'h1)))
                    begin
                      reg1747 <= ({(~"VgCx1Q9OlQf2ep")} < reg1735);
                    end
                end
            end
          for (forvar1748 = (1'h0); (forvar1748 < (1'h0)); forvar1748 = (forvar1748 + (1'h1)))
            begin
              for (forvar1749 = (1'h0); (forvar1749 < (1'h1)); forvar1749 = (forvar1749 + (1'h1)))
                begin
                  reg1750 = "wDoE8Q8YALkTl";
                  if ((8'ha4))
                    begin
                      reg1751 = $signed(($unsigned("kI6mMn") ?
                          forvar1679[(1'h1):(1'h1)] : ({(8'hb3)} & reg1623[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg1752 <= ($signed($unsigned((reg1704 ?
                              (8'haa) : (8'hb5)))) ?
                          $unsigned($unsigned($unsigned(reg1625))) : reg1741[(4'h9):(1'h0)]);
                      reg1753 = reg1745;
                      reg1754 = {$unsigned((|$unsigned((8'ha4))))};
                      reg1755 = $unsigned(reg1560[(4'ha):(3'h6)]);
                    end
                  for (forvar1756 = (1'h0); (forvar1756 < (2'h2)); forvar1756 = (forvar1756 + (1'h1)))
                    begin
                      reg1757 = reg1628;
                      reg1758 = reg1757[(1'h1):(1'h1)];
                      reg1759 <= ($unsigned(reg1669[(2'h3):(2'h3)]) ?
                          $signed("4Ktu") : (reg1672 ?
                              ((reg1742 << reg1639) ?
                                  forvar1698[(3'h4):(2'h3)] : "h6xfPgpL9Spr") : reg1742));
                      reg1760 = ($signed($signed(reg1672[(2'h3):(2'h3)])) ?
                          {(-((8'hab) - reg1553))} : reg1614[(1'h0):(1'h0)]);
                    end
                  reg1761 = $unsigned((((+(8'h9f)) << {reg1726}) >> $signed("4nwiL")));
                end
              reg1762 = {reg1564};
              reg1763 <= reg1683;
            end
          if ((~^reg1754[(1'h1):(1'h1)]))
            begin
              for (forvar1764 = (1'h0); (forvar1764 < (2'h3)); forvar1764 = (forvar1764 + (1'h1)))
                begin
                  if ((&{$unsigned($unsigned(reg1589))}))
                    begin
                      reg1765 = $signed(("3oM0rhoWe1" ?
                          reg1739[(1'h0):(1'h0)] : (~|"8J2OeKsO8Ph")));
                      reg1766 = forvar1681[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1767 <= (forvar1721 ?
                          "BEWwEfQIyXDwYVz" : (reg1751 & ("" ?
                              (wire1298 <<< (8'haa)) : (reg1701 ?
                                  reg1711 : (8'hab)))));
                      reg1768 = $signed(((+$signed((8'hb1))) << reg1731[(4'h8):(3'h6)]));
                      reg1769 = ($unsigned(((forvar1675 ?
                                  forvar1723 : reg1729) ?
                              reg1726[(1'h1):(1'h1)] : (reg1673 && wire1663))) ?
                          reg1668[(3'h4):(1'h0)] : {reg1768});
                      reg1770 = ((((~forvar1696) ?
                          {reg1685} : "iWNfBZJekL2wN") && ((reg1726 ?
                          (8'hb6) : reg1714) || (reg1737 ~^ (8'ha2)))) >>> $unsigned(reg1595));
                    end
                  reg1771 <= (forvar1746 ?
                      $unsigned($signed($signed(reg1770))) : $signed(((reg1671 ?
                              reg1691 : forvar1746) ?
                          "iSien1kIL" : (reg1553 <<< reg1754))));
                end
              if (reg1752)
                begin
                  if ($signed($unsigned(reg1768)))
                    begin
                      reg1772 = reg1750[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg1773 <= wire1296[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  reg1772 = wire1297;
                  reg1773 <= reg1742;
                  reg1774 = $signed(reg1566);
                end
              for (forvar1775 = (1'h0); (forvar1775 < (1'h1)); forvar1775 = (forvar1775 + (1'h1)))
                begin
                  for (forvar1776 = (1'h0); (forvar1776 < (2'h2)); forvar1776 = (forvar1776 + (1'h1)))
                    begin
                      reg1777 = $unsigned((!($signed(reg1687) > (~^reg1710))));
                      reg1778 = ($signed(($unsigned(reg1720) <= $unsigned(reg1710))) ?
                          reg1773[(1'h1):(1'h0)] : {reg1693[(2'h2):(1'h1)]});
                      reg1779 <= ((reg1734[(4'hd):(4'hc)] ^~ {$signed(reg1755)}) ?
                          ({forvar1713} ?
                              $signed((&reg1682)) : $unsigned({reg1726})) : (8'had));
                      reg1780 <= (8'haf);
                    end
                end
              for (forvar1781 = (1'h0); (forvar1781 < (2'h2)); forvar1781 = (forvar1781 + (1'h1)))
                begin
                  reg1782 = (8'ha2);
                  reg1783 <= (^reg1586);
                  reg1784 = (reg1545 ^~ $unsigned(((reg1688 << reg1760) ?
                      wire1663[(1'h1):(1'h1)] : (&reg1689))));
                end
            end
          else
            begin
              if (reg1636)
                begin
                  for (forvar1764 = (1'h0); (forvar1764 < (1'h0)); forvar1764 = (forvar1764 + (1'h1)))
                    begin
                      reg1767 <= $signed(("O" ?
                          (-(&reg1676)) : ($signed(reg1769) - $unsigned(reg1638))));
                      reg1771 <= ((&reg1569[(3'h5):(3'h4)]) & {(reg1729 ?
                              reg1674 : $signed(reg1771))});
                      reg1772 = $signed(($unsigned($signed(wire1295)) >>> ($signed(forvar1713) <= (~|(8'hba)))));
                      reg1774 = reg1743[(3'h4):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar1764 = (1'h0); (forvar1764 < (2'h2)); forvar1764 = (forvar1764 + (1'h1)))
                    begin
                      reg1767 <= $unsigned($signed(reg1773[(3'h7):(1'h0)]));
                    end
                  if ($signed({(8'hb9)}))
                    begin
                      reg1768 = forvar1713[(1'h0):(1'h0)];
                      reg1771 <= (^~$signed((!$unsigned(reg1683))));
                      reg1773 <= {{$unsigned((~^forvar1696))}};
                    end
                  else
                    begin
                      reg1771 <= $signed(($signed($signed(reg1641)) ~^ $unsigned((^(8'hb6)))));
                      reg1772 = ($unsigned($signed(reg1762)) ?
                          reg1755 : (reg1757[(2'h2):(2'h2)] ?
                              (reg1727 != reg1626[(1'h1):(1'h0)]) : $signed((-reg1782))));
                    end
                end
              for (forvar1775 = (1'h0); (forvar1775 < (2'h2)); forvar1775 = (forvar1775 + (1'h1)))
                begin
                  for (forvar1776 = (1'h0); (forvar1776 < (2'h2)); forvar1776 = (forvar1776 + (1'h1)))
                    begin
                      reg1779 <= (~&(-($signed((8'hb5)) <<< {(8'h9d)})));
                      reg1781 = reg1771[(4'h9):(4'h8)];
                      reg1783 <= $signed({(&{reg1703})});
                    end
                  for (forvar1784 = (1'h0); (forvar1784 < (1'h0)); forvar1784 = (forvar1784 + (1'h1)))
                    begin
                      reg1785 = (reg1709[(4'hb):(1'h1)] >= $signed(((~|reg1676) ?
                          $unsigned((8'ha0)) : {forvar1699})));
                    end
                  reg1786 = ((($unsigned((8'hb6)) << reg1550) - ("U3Fux1MFm" == wire1293[(1'h1):(1'h0)])) ?
                      (8'hb8) : reg1673[(2'h2):(1'h0)]);
                  for (forvar1787 = (1'h0); (forvar1787 < (1'h1)); forvar1787 = (forvar1787 + (1'h1)))
                    begin
                      reg1788 = "2Iu5";
                      reg1789 = ({$signed($signed((8'ha3)))} ?
                          (~|(|(8'hb9))) : wire1296);
                      reg1790 <= forvar1746[(2'h3):(2'h3)];
                      reg1791 = $unsigned($signed($unsigned(forvar1707[(3'h6):(2'h3)])));
                    end
                end
              for (forvar1792 = (1'h0); (forvar1792 < (1'h0)); forvar1792 = (forvar1792 + (1'h1)))
                begin
                  reg1793 = reg1762;
                  reg1794 = $signed(forvar1784);
                end
            end
        end
      else
        begin
          reg1721 <= ("V" + "thJ");
          for (forvar1722 = (1'h0); (forvar1722 < (2'h2)); forvar1722 = (forvar1722 + (1'h1)))
            begin
              for (forvar1723 = (1'h0); (forvar1723 < (1'h0)); forvar1723 = (forvar1723 + (1'h1)))
                begin
                  reg1727 = reg1641;
                end
            end
        end
      if ((&$unsigned((+(reg1589 ? reg1745 : forvar1781)))))
        begin
          reg1795 = ($signed(($unsigned(reg1717) - (^~(8'hb1)))) ?
              $unsigned(reg1661) : forvar1692);
          if (($signed(reg1583[(3'h5):(3'h4)]) ?
              reg1639 : $signed($signed(reg1545))))
            begin
              if ($unsigned($unsigned(reg1678)))
                begin
                  for (forvar1796 = (1'h0); (forvar1796 < (2'h2)); forvar1796 = (forvar1796 + (1'h1)))
                    begin
                      reg1797 = reg1753[(2'h2):(1'h1)];
                      reg1798 = {reg1700[(3'h6):(3'h5)]};
                    end
                  reg1799 = (8'hb3);
                  reg1800 = {($signed(((8'hae) ?
                          forvar1698 : reg1725)) && reg1758[(4'he):(4'h8)])};
                  for (forvar1801 = (1'h0); (forvar1801 < (2'h3)); forvar1801 = (forvar1801 + (1'h1)))
                    begin
                      reg1802 <= ($signed(reg1701[(2'h3):(2'h2)]) ?
                          reg1625[(1'h0):(1'h0)] : reg1784);
                      reg1803 <= $signed((("1mfQlBf" ?
                          (|forvar1723) : {reg1778}) != $unsigned($unsigned(reg1668))));
                    end
                end
              else
                begin
                  for (forvar1796 = (1'h0); (forvar1796 < (1'h0)); forvar1796 = (forvar1796 + (1'h1)))
                    begin
                      reg1801 <= forvar1698;
                      reg1804 = reg1555;
                      reg1805 <= $signed(reg1614[(1'h0):(1'h0)]);
                      reg1806 <= $signed(reg1641[(1'h1):(1'h1)]);
                    end
                  reg1807 <= reg1677[(4'hd):(4'ha)];
                end
              for (forvar1808 = (1'h0); (forvar1808 < (1'h1)); forvar1808 = (forvar1808 + (1'h1)))
                begin
                  for (forvar1809 = (1'h0); (forvar1809 < (2'h2)); forvar1809 = (forvar1809 + (1'h1)))
                    begin
                      reg1810 = "Gf";
                    end
                  reg1811 = $unsigned("HfdhHZzaD7boRt");
                  for (forvar1812 = (1'h0); (forvar1812 < (2'h2)); forvar1812 = (forvar1812 + (1'h1)))
                    begin
                      reg1813 <= (forvar1746 ? reg1580 : wire1556);
                    end
                end
              if (reg1574)
                begin
                  for (forvar1814 = (1'h0); (forvar1814 < (1'h1)); forvar1814 = (forvar1814 + (1'h1)))
                    begin
                      reg1815 = (^~reg1717[(2'h2):(2'h2)]);
                      reg1816 = wire1296;
                    end
                end
              else
                begin
                  reg1814 = (|$unsigned(((^reg1771) < $unsigned(reg1759))));
                  if (reg1720[(2'h2):(2'h2)])
                    begin
                      reg1817 <= reg1777[(4'h9):(3'h7)];
                    end
                  else
                    begin
                      reg1815 = $unsigned((reg1645[(3'h4):(3'h4)] ?
                          ({reg1638} > (forvar1740 >= reg1589)) : (8'ha6)));
                      reg1816 = ($signed((8'hb3)) ?
                          reg1790[(3'h5):(1'h1)] : $unsigned(forvar1781[(1'h1):(1'h0)]));
                      reg1817 <= reg1638[(3'h5):(3'h4)];
                    end
                end
              reg1818 = ($unsigned(reg1608) ?
                  forvar1707 : $signed($unsigned("FbsUM7BhB1GHp")));
            end
          else
            begin
              reg1796 <= $signed(forvar1718);
              if ((+$unsigned((&"98B7m5M3e0w"))))
                begin
                  if ($unsigned("V0GMmiQ"))
                    begin
                      reg1797 = reg1709;
                      reg1798 = $unsigned((!{forvar1721[(4'he):(4'hb)]}));
                      reg1799 = reg1711;
                    end
                  else
                    begin
                      reg1797 = $unsigned($unsigned(("AJ5k5Y7GFz6" * (reg1795 ?
                          reg1645 : reg1811))));
                      reg1801 <= $signed($unsigned((^reg1639[(1'h1):(1'h0)])));
                    end
                end
              else
                begin
                  reg1797 = forvar1699;
                end
              for (forvar1802 = (1'h0); (forvar1802 < (1'h0)); forvar1802 = (forvar1802 + (1'h1)))
                begin
                  reg1803 <= (^~reg1802);
                  reg1804 = (8'h9d);
                  if (reg1569)
                    begin
                      reg1805 <= ((!$unsigned((|reg1762))) + "DZKp4inb");
                      reg1806 <= $signed({"itvQs3v78qM"});
                      reg1807 <= reg1733[(4'ha):(4'ha)];
                      reg1808 = ({{(reg1797 ?
                                  reg1797 : reg1552)}} ^ "zI8OgK763zesvL");
                    end
                  else
                    begin
                      reg1805 <= ((reg1731[(3'h7):(2'h3)] ?
                          (|(reg1628 ^ reg1553)) : $signed(reg1688[(2'h3):(2'h2)])) ^~ reg1583[(2'h3):(1'h1)]);
                      reg1806 <= {"SzbubPHhBDLW"};
                    end
                end
              if ((&(|(~reg1670))))
                begin
                  if ($signed("rITJi8"))
                    begin
                      reg1809 = ("FPqaqG" & $signed($signed(reg1811)));
                      reg1810 = ($signed($unsigned((reg1575 || reg1779))) ?
                          $unsigned($unsigned(wire1294[(3'h7):(1'h0)])) : (!(8'hb2)));
                      reg1811 = (reg1702 ?
                          reg1684[(2'h2):(1'h0)] : reg1623[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1809 = reg1790[(3'h6):(3'h4)];
                      reg1810 = forvar1679[(1'h1):(1'h1)];
                    end
                  reg1812 <= ($unsigned($unsigned((reg1736 ?
                          (8'ha3) : reg1682))) ?
                      $unsigned("eWrkFflkHFv") : (~^$signed(reg1784[(2'h2):(1'h1)])));
                  reg1814 = (~^forvar1781);
                end
              else
                begin
                  reg1809 = "A";
                  for (forvar1810 = (1'h0); (forvar1810 < (2'h2)); forvar1810 = (forvar1810 + (1'h1)))
                    begin
                      reg1812 <= $unsigned(({(reg1683 < (8'hba))} ?
                          "Sn" : {(^reg1731)}));
                      reg1814 = $signed(reg1763);
                    end
                  for (forvar1815 = (1'h0); (forvar1815 < (1'h1)); forvar1815 = (forvar1815 + (1'h1)))
                    begin
                      reg1816 = reg1695[(1'h1):(1'h0)];
                      reg1818 = "kqlyvLGad3uDxmN";
                      reg1819 = $unsigned((reg1810[(1'h1):(1'h1)] ?
                          (^"z0tXXk") : $unsigned($unsigned(forvar1746))));
                      reg1820 <= (((^reg1572) || "EeRbIhDv7W") < (($signed((8'hb6)) < "FMFkfpYx41i") == (~$signed(reg1813))));
                    end
                  for (forvar1821 = (1'h0); (forvar1821 < (2'h2)); forvar1821 = (forvar1821 + (1'h1)))
                    begin
                      reg1822 = {reg1584};
                    end
                end
            end
          for (forvar1823 = (1'h0); (forvar1823 < (2'h3)); forvar1823 = (forvar1823 + (1'h1)))
            begin
              for (forvar1824 = (1'h0); (forvar1824 < (1'h1)); forvar1824 = (forvar1824 + (1'h1)))
                begin
                  for (forvar1825 = (1'h0); (forvar1825 < (1'h1)); forvar1825 = (forvar1825 + (1'h1)))
                    begin
                      reg1826 <= forvar1721[(2'h2):(1'h1)];
                      reg1827 <= (-(8'ha0));
                      reg1828 = $signed("LaLA4a7Om");
                    end
                end
            end
          if (reg1799[(2'h3):(2'h3)])
            begin
              reg1829 <= reg1814[(4'h8):(3'h6)];
              reg1830 = $signed(reg1750);
            end
          else
            begin
              for (forvar1829 = (1'h0); (forvar1829 < (2'h3)); forvar1829 = (forvar1829 + (1'h1)))
                begin
                  reg1831 <= (8'hb8);
                  for (forvar1832 = (1'h0); (forvar1832 < (2'h2)); forvar1832 = (forvar1832 + (1'h1)))
                    begin
                      reg1833 <= forvar1690;
                      reg1834 = forvar1825[(1'h0):(1'h0)];
                    end
                  for (forvar1835 = (1'h0); (forvar1835 < (1'h0)); forvar1835 = (forvar1835 + (1'h1)))
                    begin
                      reg1836 = $signed({wire1299});
                    end
                  reg1837 = reg1830[(1'h0):(1'h0)];
                end
              reg1838 = $unsigned("KqJy9vh");
              for (forvar1839 = (1'h0); (forvar1839 < (2'h3)); forvar1839 = (forvar1839 + (1'h1)))
                begin
                  reg1840 = $signed((8'haa));
                  for (forvar1841 = (1'h0); (forvar1841 < (1'h1)); forvar1841 = (forvar1841 + (1'h1)))
                    begin
                      reg1842 <= {(reg1768 ?
                              {{reg1765}} : {$unsigned(reg1723)})};
                    end
                  if (($unsigned((~|$unsigned(reg1668))) || (8'hb8)))
                    begin
                      reg1843 = {(-(~&$unsigned(reg1694)))};
                      reg1844 = reg1702[(4'hd):(4'h9)];
                      reg1845 = ($unsigned(reg1683[(3'h5):(2'h3)]) + (reg1550[(3'h7):(3'h5)] ?
                          (forvar1748[(2'h3):(2'h3)] ?
                              reg1757 : $signed(reg1804)) : $signed($unsigned((8'ha2)))));
                      reg1846 <= "";
                    end
                  else
                    begin
                      reg1843 = (-((forvar1764 ?
                              $signed(reg1722) : ((8'had) ?
                                  forvar1781 : forvar1721)) ?
                          "xefwHGSXu5t" : reg1641));
                      reg1846 <= $signed(reg1649);
                    end
                end
            end
        end
      else
        begin
          reg1796 <= (reg1643 ?
              (+(8'ha5)) : (reg1712[(3'h5):(1'h1)] << (forvar1699 ?
                  $unsigned(reg1755) : {reg1767})));
          if (($unsigned((forvar1810[(4'hd):(1'h0)] ~^ (~^reg1774))) ?
              reg1566 : "Ia9U66MsJJpVTn"))
            begin
              reg1797 = reg1677[(3'h6):(3'h6)];
              for (forvar1798 = (1'h0); (forvar1798 < (1'h1)); forvar1798 = (forvar1798 + (1'h1)))
                begin
                  reg1801 <= (($signed($signed(reg1705)) ?
                      $unsigned(((8'hb1) ?
                          (8'haa) : reg1552)) : "yie") * $unsigned(reg1842));
                  if ((~((+forvar1748) <= reg1793[(2'h2):(1'h1)])))
                    begin
                      reg1804 = {forvar1722[(3'h5):(1'h1)]};
                    end
                  else
                    begin
                      reg1804 = reg1687;
                      reg1805 <= $signed(((forvar1666[(3'h4):(1'h1)] >> reg1809) - ({reg1830} ?
                          reg1688[(1'h1):(1'h1)] : $signed(reg1543))));
                    end
                  reg1808 = ($unsigned("XDdL2x6N4tlbJ") ?
                      "U" : (($unsigned((8'haa)) >> (reg1619 - reg1639)) | ($unsigned(reg1703) ?
                          "f7d" : $signed(reg1632))));
                  reg1812 <= $signed("eUGc1");
                end
            end
          else
            begin
              if ((8'hb7))
                begin
                  reg1797 = (~{$unsigned(reg1589[(3'h6):(2'h3)])});
                  if ($signed(($unsigned({(8'hb0)}) & (|(^reg1623)))))
                    begin
                      reg1798 = ("9aPhZ" ?
                          reg1834 : ($signed(reg1751) <<< reg1571[(4'ha):(3'h7)]));
                      reg1801 <= reg1703[(2'h3):(2'h3)];
                      reg1804 = (({(&forvar1776)} ?
                              ((|reg1765) ?
                                  $unsigned(reg1569) : $signed(forvar1679)) : {{forvar1784}}) ?
                          reg1799 : ((&"0N0DP") ^~ (!((8'haa) ?
                              wire1663 : reg1769))));
                    end
                  else
                    begin
                      reg1801 <= (reg1694 << $signed(forvar1749[(3'h6):(1'h0)]));
                      reg1804 = ((^reg1815[(2'h2):(2'h2)]) < $signed(reg1771[(4'h9):(3'h7)]));
                      reg1808 = $unsigned(forvar1740);
                      reg1809 = "";
                    end
                end
              else
                begin
                  reg1801 <= (^($signed((^reg1733)) <<< reg1836));
                end
              if ((^~(($signed(reg1837) <= reg1550) | $signed(reg1735))))
                begin
                  reg1810 = $signed($signed(forvar1679[(2'h3):(2'h3)]));
                  reg1811 = "";
                  if (wire1292[(2'h3):(2'h2)])
                    begin
                      reg1814 = forvar1781[(1'h0):(1'h0)];
                      reg1815 = $unsigned((~^(((8'ha5) - (8'ha5)) ?
                          (8'hb9) : $unsigned(reg1608))));
                      reg1816 = forvar1740[(3'h4):(2'h3)];
                      reg1817 <= "9I4tCENU3ROZVa";
                    end
                  else
                    begin
                      reg1814 = $unsigned(({{reg1706}} ?
                          reg1636 : ((reg1702 && reg1649) ^~ (8'ha6))));
                      reg1815 = $signed(($unsigned((reg1717 - (8'ha7))) ?
                          ($unsigned(reg1715) ?
                              (reg1819 && forvar1787) : (-reg1797)) : "aAXurVm2YIkh3k"));
                      reg1816 = forvar1841;
                      reg1818 = (~|{((wire1296 >> forvar1686) ?
                              "5s" : $unsigned(reg1574))});
                    end
                end
              else
                begin
                  reg1810 = $signed((((|reg1560) ?
                          $signed(forvar1699) : (^~reg1570)) ?
                      forvar1824 : reg1768));
                  if ("y7o")
                    begin
                      reg1812 <= "H1GlDiPr51M";
                    end
                  else
                    begin
                      reg1811 = ({$signed(reg1595)} && (~&reg1834[(3'h5):(2'h2)]));
                      reg1814 = reg1763;
                      reg1817 <= (($unsigned($unsigned(reg1728)) <= reg1702) ?
                          (+($unsigned(forvar1835) ?
                              {reg1626} : reg1830)) : reg1751[(3'h6):(2'h3)]);
                    end
                end
            end
          for (forvar1819 = (1'h0); (forvar1819 < (2'h3)); forvar1819 = (forvar1819 + (1'h1)))
            begin
              reg1821 = forvar1666;
            end
        end
    end
  assign wire1847 = reg1661[(4'hd):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1300  (y, clk, wire1305, wire1304, wire1303, wire1302, wire1301);
  output wire [(32'h955):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire1305;
  input wire [(4'hf):(1'h0)] wire1304;
  input wire signed [(4'hb):(1'h0)] wire1303;
  input wire signed [(4'hf):(1'h0)] wire1302;
  input wire [(3'h5):(1'h0)] wire1301;
  wire signed [(4'h9):(1'h0)] wire1498;
  wire [(4'h8):(1'h0)] wire1497;
  wire [(4'he):(1'h0)] wire1496;
  wire signed [(3'h4):(1'h0)] wire1371;
  wire [(4'he):(1'h0)] wire1347;
  wire signed [(3'h4):(1'h0)] wire1307;
  wire [(2'h2):(1'h0)] wire1306;
  reg signed [(3'h4):(1'h0)] reg1535 = (1'h0);
  reg [(4'he):(1'h0)] reg1532 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1530 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1526 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1521 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1520 = (1'h0);
  reg [(5'h10):(1'h0)] reg1519 = (1'h0);
  reg [(4'hb):(1'h0)] reg1513 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1511 = (1'h0);
  reg [(3'h5):(1'h0)] reg1506 = (1'h0);
  reg [(2'h2):(1'h0)] reg1505 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1503 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1492 = (1'h0);
  reg [(4'ha):(1'h0)] reg1490 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1489 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1479 = (1'h0);
  reg [(3'h7):(1'h0)] reg1477 = (1'h0);
  reg [(4'h9):(1'h0)] reg1474 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1467 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1457 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1438 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1460 = (1'h0);
  reg [(2'h3):(1'h0)] reg1453 = (1'h0);
  reg [(4'hf):(1'h0)] reg1447 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1444 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1436 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1432 = (1'h0);
  reg [(4'h9):(1'h0)] reg1430 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1423 = (1'h0);
  reg [(4'hc):(1'h0)] reg1421 = (1'h0);
  reg [(4'hd):(1'h0)] reg1418 = (1'h0);
  reg [(4'h8):(1'h0)] reg1415 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1412 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1406 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1404 = (1'h0);
  reg [(4'hc):(1'h0)] reg1401 = (1'h0);
  reg [(3'h7):(1'h0)] reg1400 = (1'h0);
  reg [(4'ha):(1'h0)] reg1399 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1396 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1391 = (1'h0);
  reg [(4'he):(1'h0)] reg1390 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1385 = (1'h0);
  reg [(2'h2):(1'h0)] reg1378 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1374 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1368 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1365 = (1'h0);
  reg [(3'h4):(1'h0)] reg1363 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1358 = (1'h0);
  reg [(4'he):(1'h0)] reg1361 = (1'h0);
  reg [(3'h6):(1'h0)] reg1359 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1354 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1352 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1351 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1342 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1340 = (1'h0);
  reg [(4'he):(1'h0)] reg1339 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1337 = (1'h0);
  reg [(3'h5):(1'h0)] reg1332 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1327 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1324 = (1'h0);
  reg [(4'hb):(1'h0)] reg1323 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1319 = (1'h0);
  reg [(4'he):(1'h0)] reg1315 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1310 = (1'h0);
  reg [(3'h4):(1'h0)] reg1312 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1309 = (1'h0);
  reg [(4'hd):(1'h0)] reg1537 = (1'h0);
  reg [(4'hf):(1'h0)] reg1536 = (1'h0);
  reg [(2'h2):(1'h0)] reg1534 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1533 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1531 = (1'h0);
  reg [(3'h5):(1'h0)] reg1529 = (1'h0);
  reg [(4'hd):(1'h0)] reg1528 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1527 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1516 = (1'h0);
  reg [(2'h2):(1'h0)] reg1525 = (1'h0);
  reg [(4'h9):(1'h0)] reg1524 = (1'h0);
  reg [(4'he):(1'h0)] reg1523 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1522 = (1'h0);
  reg [(4'hd):(1'h0)] reg1518 = (1'h0);
  reg [(4'hb):(1'h0)] reg1517 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1516 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1515 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1514 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1512 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1510 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1509 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1508 = (1'h0);
  reg [(4'hf):(1'h0)] reg1507 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1504 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1502 = (1'h0);
  reg [(3'h4):(1'h0)] reg1501 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1500 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1499 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1495 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1494 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1493 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1491 = (1'h0);
  reg [(4'hd):(1'h0)] reg1488 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1487 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1486 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1485 = (1'h0);
  reg [(4'hc):(1'h0)] reg1484 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1483 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1482 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1481 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1480 = (1'h0);
  reg [(5'h10):(1'h0)] reg1478 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1475 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1473 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1471 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1476 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1475 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1473 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1472 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1471 = (1'h0);
  reg [(4'h8):(1'h0)] reg1470 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1469 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1468 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1466 = (1'h0);
  reg [(3'h5):(1'h0)] reg1465 = (1'h0);
  reg [(4'ha):(1'h0)] reg1464 = (1'h0);
  reg [(4'he):(1'h0)] forvar1463 = (1'h0);
  reg [(4'he):(1'h0)] forvar1456 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1458 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1452 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1446 = (1'h0);
  reg [(4'he):(1'h0)] forvar1445 = (1'h0);
  reg [(4'hd):(1'h0)] reg1439 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1440 = (1'h0);
  reg [(4'hd):(1'h0)] reg1463 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1462 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1461 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1459 = (1'h0);
  reg [(4'hf):(1'h0)] reg1458 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1457 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1456 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1455 = (1'h0);
  reg [(3'h6):(1'h0)] reg1454 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1452 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1451 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1450 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1449 = (1'h0);
  reg [(4'hd):(1'h0)] reg1448 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1446 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1445 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1443 = (1'h0);
  reg [(4'ha):(1'h0)] reg1442 = (1'h0);
  reg [(4'h9):(1'h0)] reg1441 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1440 = (1'h0);
  reg [(4'he):(1'h0)] forvar1439 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1438 = (1'h0);
  reg [(4'hc):(1'h0)] reg1437 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1435 = (1'h0);
  reg [(4'hf):(1'h0)] reg1434 = (1'h0);
  reg [(2'h3):(1'h0)] reg1433 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1431 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1429 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1428 = (1'h0);
  reg [(2'h2):(1'h0)] reg1427 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1426 = (1'h0);
  reg [(3'h5):(1'h0)] reg1425 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1423 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1424 = (1'h0);
  reg [(3'h6):(1'h0)] reg1422 = (1'h0);
  reg [(4'h8):(1'h0)] reg1420 = (1'h0);
  reg [(4'hc):(1'h0)] reg1419 = (1'h0);
  reg [(2'h3):(1'h0)] reg1417 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1416 = (1'h0);
  reg [(4'h9):(1'h0)] reg1414 = (1'h0);
  reg [(3'h5):(1'h0)] reg1413 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1411 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1411 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1410 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1409 = (1'h0);
  reg [(4'h8):(1'h0)] reg1408 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1397 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1393 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1407 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1405 = (1'h0);
  reg [(3'h7):(1'h0)] reg1403 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1402 = (1'h0);
  reg [(3'h4):(1'h0)] reg1398 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1397 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1395 = (1'h0);
  reg [(4'hc):(1'h0)] reg1394 = (1'h0);
  reg [(4'hd):(1'h0)] reg1393 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1392 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1389 = (1'h0);
  reg [(2'h3):(1'h0)] reg1388 = (1'h0);
  reg [(4'hc):(1'h0)] reg1387 = (1'h0);
  reg [(4'h9):(1'h0)] reg1386 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1384 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1383 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1382 = (1'h0);
  reg [(4'he):(1'h0)] forvar1381 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1380 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1379 = (1'h0);
  reg [(4'he):(1'h0)] reg1377 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1376 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1375 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1373 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1372 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1370 = (1'h0);
  reg [(5'h10):(1'h0)] reg1369 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1367 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1366 = (1'h0);
  reg [(3'h5):(1'h0)] reg1364 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1361 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1354 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1353 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1352 = (1'h0);
  reg [(4'h9):(1'h0)] reg1362 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1360 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1358 = (1'h0);
  reg [(3'h6):(1'h0)] reg1348 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1357 = (1'h0);
  reg [(2'h2):(1'h0)] reg1356 = (1'h0);
  reg [(4'he):(1'h0)] reg1355 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1353 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1350 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1349 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1348 = (1'h0);
  reg [(3'h6):(1'h0)] reg1343 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1342 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1341 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1346 = (1'h0);
  reg [(4'ha):(1'h0)] reg1345 = (1'h0);
  reg [(3'h4):(1'h0)] reg1344 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1343 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1341 = (1'h0);
  reg [(5'h10):(1'h0)] reg1338 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1336 = (1'h0);
  reg [(4'hd):(1'h0)] reg1335 = (1'h0);
  reg [(3'h4):(1'h0)] reg1334 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1333 = (1'h0);
  reg [(4'hb):(1'h0)] reg1331 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1330 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1326 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1320 = (1'h0);
  reg [(4'he):(1'h0)] reg1317 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1329 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1328 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1327 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1326 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1325 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1322 = (1'h0);
  reg [(4'hf):(1'h0)] reg1321 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1320 = (1'h0);
  reg [(3'h5):(1'h0)] reg1318 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1317 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1316 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1311 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1314 = (1'h0);
  reg [(2'h3):(1'h0)] reg1313 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1311 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1310 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1308 = (1'h0);
  assign y = {wire1496,
                 wire1371,
                 wire1347,
                 wire1307,
                 reg1530,
                 reg1526,
                 reg1519,
                 reg1511,
                 reg1505,
                 reg1503,
                 reg1489,
                 reg1479,
                 reg1457,
                 reg1460,
                 reg1453,
                 reg1432,
                 reg1412,
                 reg1400,
                 reg1396,
                 reg1390,
                 reg1385,
                 reg1374,
                 reg1368,
                 reg1363,
                 reg1358,
                 reg1361,
                 reg1359,
                 reg1351,
                 reg1342,
                 reg1332,
                 reg1323,
                 reg1310,
                 reg1536,
                 forvar1531,
                 reg1529,
                 forvar1516,
                 reg1518,
                 forvar1515,
                 reg1514,
                 forvar1510,
                 forvar1504,
                 forvar1502,
                 reg1495,
                 forvar1482,
                 reg1481,
                 forvar1475,
                 reg1475,
                 reg1472,
                 reg1470,
                 forvar1469,
                 forvar1468,
                 reg1466,
                 reg1464,
                 forvar1458,
                 reg1458,
                 forvar1457,
                 reg1456,
                 reg1454,
                 forvar1452,
                 reg1449,
                 reg1448,
                 forvar1439,
                 reg1434,
                 reg1433,
                 forvar1423,
                 reg1424,
                 reg1422,
                 reg1420,
                 reg1419,
                 reg1417,
                 reg1414,
                 reg1413,
                 forvar1411,
                 reg1411,
                 forvar1409,
                 reg1408,
                 reg1397,
                 forvar1392,
                 forvar1381,
                 reg1380,
                 forvar1376,
                 forvar1375,
                 forvar1372,
                 reg1348,
                 forvar1353,
                 forvar1341,
                 reg1335,
                 reg1334,
                 forvar1333,
                 reg1331,
                 reg1317,
                 reg1328,
                 reg1326,
                 reg1325,
                 reg1320,
                 reg1318,
                 reg1316,
                 reg1314,
                 (1'h0)};
  assign wire1306 = (wire1305 && $unsigned(({wire1303} ?
                        wire1305[(2'h2):(1'h1)] : $signed(wire1302))));
  assign wire1307 = (~^$signed($unsigned((wire1303 ? wire1302 : (8'hb7)))));
  always
    @(posedge clk) begin
      for (forvar1308 = (1'h0); (forvar1308 < (1'h0)); forvar1308 = (forvar1308 + (1'h1)))
        begin
          if ((~forvar1308))
            begin
              reg1309 <= ((^wire1303[(3'h4):(2'h2)]) >> ($signed((forvar1308 ?
                  wire1301 : wire1301)) >= ((wire1302 ?
                      forvar1308 : forvar1308) ?
                  (8'ha6) : $signed(wire1304))));
              if ((~wire1301[(3'h5):(3'h5)]))
                begin
                  for (forvar1310 = (1'h0); (forvar1310 < (2'h3)); forvar1310 = (forvar1310 + (1'h1)))
                    begin
                      reg1311 = (wire1302[(1'h1):(1'h0)] ?
                          (8'ha4) : $unsigned($signed((|reg1309))));
                      reg1312 <= $signed($unsigned(wire1301));
                      reg1313 = wire1301[(3'h5):(3'h4)];
                      reg1314 = wire1302;
                    end
                end
              else
                begin
                  reg1310 <= (-($unsigned($unsigned((8'hba))) ^~ reg1312[(2'h3):(2'h3)]));
                  for (forvar1311 = (1'h0); (forvar1311 < (2'h2)); forvar1311 = (forvar1311 + (1'h1)))
                    begin
                      reg1313 = "M";
                      reg1314 = {{$unsigned($unsigned(forvar1308))}};
                      reg1315 <= $signed((^wire1301[(2'h3):(1'h1)]));
                    end
                end
              reg1316 = $signed((wire1304[(3'h5):(1'h1)] ^ wire1301[(1'h0):(1'h0)]));
              for (forvar1317 = (1'h0); (forvar1317 < (1'h0)); forvar1317 = (forvar1317 + (1'h1)))
                begin
                  reg1318 = reg1313[(2'h2):(1'h1)];
                  if ($unsigned(("CbyA5fFdYR" >= (-(-forvar1311)))))
                    begin
                      reg1319 <= $signed($signed($signed(reg1312)));
                      reg1320 = $unsigned($unsigned({wire1306[(1'h0):(1'h0)]}));
                      reg1321 = "g9JYSAp5Lw";
                    end
                  else
                    begin
                      reg1319 <= forvar1310;
                      reg1320 = ("rLo2zx1vIU4T" ?
                          (reg1310[(4'hc):(4'h8)] || (&$signed(reg1315))) : $signed((+$signed(reg1309))));
                    end
                  if (reg1315)
                    begin
                      reg1322 = $signed((((wire1304 ? forvar1317 : reg1321) ?
                          wire1307[(1'h1):(1'h1)] : $unsigned(reg1316)) >> ("0Bxiz5BdEh" ?
                          $unsigned(wire1307) : reg1315[(2'h3):(1'h0)])));
                      reg1323 <= (^((&wire1304[(4'hd):(4'hc)]) ?
                          (wire1301[(3'h5):(3'h4)] ?
                              (reg1321 ?
                                  wire1301 : reg1322) : (wire1302 || reg1312)) : (8'ha2)));
                      reg1324 <= ((8'hb4) * ($unsigned((~|(8'h9e))) ?
                          (reg1311 <<< reg1312[(2'h2):(1'h0)]) : ((&forvar1317) ?
                              ((8'ha0) == wire1305) : (wire1301 | wire1306))));
                    end
                  else
                    begin
                      reg1323 <= (((+{reg1315}) ?
                          $signed($signed(wire1305)) : "QXW") ^~ reg1318[(1'h1):(1'h0)]);
                      reg1325 = reg1324[(1'h1):(1'h1)];
                      reg1326 = $signed($unsigned(wire1304));
                    end
                  for (forvar1327 = (1'h0); (forvar1327 < (1'h0)); forvar1327 = (forvar1327 + (1'h1)))
                    begin
                      reg1328 = forvar1327;
                      reg1329 = $signed({wire1301});
                    end
                end
            end
          else
            begin
              reg1309 <= (forvar1317 ^ ($signed((reg1318 ?
                  reg1326 : (8'had))) ~^ reg1328[(2'h2):(1'h0)]));
              for (forvar1310 = (1'h0); (forvar1310 < (2'h3)); forvar1310 = (forvar1310 + (1'h1)))
                begin
                  reg1311 = ((-{"2oxRZtI46"}) ?
                      $signed(({reg1328} ?
                          $unsigned(forvar1308) : ((8'hb1) ^ reg1321))) : reg1313);
                end
              if ((reg1314 ?
                  reg1309[(1'h0):(1'h0)] : (((reg1311 ? reg1318 : forvar1327) ?
                          $unsigned(reg1314) : (8'hae)) ?
                      reg1316[(1'h0):(1'h0)] : "RxoqtZDAeW")))
                begin
                  if ("")
                    begin
                      reg1312 <= $unsigned(reg1323);
                      reg1315 <= $unsigned(({(reg1320 ? reg1326 : wire1302)} ?
                          $signed((wire1301 ?
                              reg1319 : reg1321)) : $signed("Q4yYIhnt2KK")));
                      reg1316 = "";
                      reg1317 = reg1311;
                    end
                  else
                    begin
                      reg1312 <= (~|$signed($unsigned((&forvar1308))));
                      reg1315 <= ((8'hae) ? reg1312[(1'h0):(1'h0)] : reg1326);
                      reg1319 <= ((wire1301 ?
                              reg1326[(2'h3):(2'h2)] : $unsigned($signed(reg1329))) ?
                          ((-(forvar1317 >> wire1304)) ?
                              (((8'hb3) + wire1305) - forvar1327) : (^reg1324)) : $unsigned(($unsigned(reg1325) ?
                              $signed(reg1310) : reg1319[(4'ha):(4'h9)])));
                    end
                  for (forvar1320 = (1'h0); (forvar1320 < (1'h0)); forvar1320 = (forvar1320 + (1'h1)))
                    begin
                      reg1321 = (8'ha4);
                    end
                  reg1323 <= $signed((-reg1323[(1'h0):(1'h0)]));
                end
              else
                begin
                  if ((~^(({wire1307} == forvar1310) ?
                      "4n8" : "TTDF6ymg3fMsRu")))
                    begin
                      reg1313 = "NKfC";
                    end
                  else
                    begin
                      reg1313 = reg1312[(1'h1):(1'h1)];
                    end
                  reg1315 <= $unsigned({reg1326[(4'h9):(4'h8)]});
                  if (((~wire1307[(3'h4):(1'h1)]) ?
                      $unsigned({{(8'hba)}}) : $unsigned((8'hb2))))
                    begin
                      reg1316 = (^~(8'hb7));
                      reg1319 <= $unsigned({reg1323});
                      reg1320 = (+(forvar1317 * {(reg1323 ?
                              wire1307 : (8'h9d))}));
                    end
                  else
                    begin
                      reg1319 <= reg1324;
                      reg1323 <= $unsigned((|forvar1327));
                      reg1325 = (~^"BwCcXewuC");
                    end
                  for (forvar1326 = (1'h0); (forvar1326 < (2'h2)); forvar1326 = (forvar1326 + (1'h1)))
                    begin
                      reg1327 <= $signed($signed((^~(reg1323 > forvar1320))));
                      reg1328 = reg1312[(1'h1):(1'h1)];
                      reg1329 = $unsigned({($signed(reg1322) ?
                              (forvar1320 & reg1318) : {wire1306})});
                    end
                end
            end
          for (forvar1330 = (1'h0); (forvar1330 < (1'h0)); forvar1330 = (forvar1330 + (1'h1)))
            begin
              reg1331 = reg1322[(3'h7):(3'h7)];
              reg1332 <= (-reg1313);
              for (forvar1333 = (1'h0); (forvar1333 < (2'h2)); forvar1333 = (forvar1333 + (1'h1)))
                begin
                  if (({((~&reg1332) && (wire1302 > reg1326))} ?
                      wire1303 : reg1315[(3'h5):(3'h4)]))
                    begin
                      reg1334 = $unsigned({($signed((8'ha6)) >= reg1312[(3'h4):(1'h1)])});
                    end
                  else
                    begin
                      reg1334 = $signed(wire1302[(3'h4):(3'h4)]);
                      reg1335 = reg1321[(1'h0):(1'h0)];
                      reg1336 = ({$unsigned($unsigned(wire1304))} == reg1331[(2'h3):(2'h3)]);
                    end
                  reg1337 <= wire1307[(1'h1):(1'h0)];
                end
            end
          if ($unsigned(""))
            begin
              reg1338 = {($unsigned((reg1336 >> reg1318)) ?
                      reg1311 : (reg1322 <<< $unsigned(wire1307)))};
            end
          else
            begin
              if (({(~&reg1334[(2'h3):(2'h2)])} ?
                  {$unsigned(reg1325)} : {(((8'hb4) >= forvar1317) < $unsigned(wire1302))}))
                begin
                  if ((reg1317 | ("LVn1TCpiItDvid" ? "6" : reg1318)))
                    begin
                      reg1339 <= reg1335;
                      reg1340 <= ((("s" != ((8'hb9) < forvar1320)) || {(reg1318 >> wire1307)}) < {(~^(-forvar1327))});
                    end
                  else
                    begin
                      reg1338 = ($signed($signed((reg1335 > (8'ha3)))) ?
                          ("L5dOZvZC" ?
                              ((8'ha1) ?
                                  (reg1326 ? forvar1330 : reg1309) : (reg1339 ?
                                      reg1310 : reg1329)) : "a96v") : "xJdSJ2vIkfbMJd7");
                    end
                  for (forvar1341 = (1'h0); (forvar1341 < (2'h3)); forvar1341 = (forvar1341 + (1'h1)))
                    begin
                      reg1342 <= "JFk";
                    end
                  for (forvar1343 = (1'h0); (forvar1343 < (2'h2)); forvar1343 = (forvar1343 + (1'h1)))
                    begin
                      reg1344 = $unsigned(("TsRZX4H" * (reg1318 ?
                          (|reg1332) : reg1340[(4'h9):(2'h2)])));
                      reg1345 = $signed("Ko");
                      reg1346 = (((|(|(8'hb8))) ?
                          $signed((forvar1308 ?
                              reg1329 : reg1324)) : ((&reg1334) ?
                              $unsigned(forvar1341) : (wire1305 > (8'haf)))) != {forvar1317});
                    end
                end
              else
                begin
                  reg1338 = $unsigned((reg1326[(1'h1):(1'h1)] && {(forvar1343 != wire1302)}));
                  reg1341 = ((((reg1331 ^~ forvar1341) < (reg1331 ?
                      forvar1333 : reg1338)) ~^ ((-reg1336) ?
                      forvar1311[(1'h1):(1'h1)] : (forvar1311 && wire1304))) ^~ (((reg1323 + forvar1311) < (!reg1332)) ?
                      forvar1317[(3'h5):(3'h4)] : $signed((reg1316 ?
                          reg1319 : reg1310))));
                  for (forvar1342 = (1'h0); (forvar1342 < (2'h3)); forvar1342 = (forvar1342 + (1'h1)))
                    begin
                      reg1343 = reg1325[(2'h3):(2'h2)];
                    end
                  reg1344 = ("sMzze" ?
                      forvar1326 : $unsigned(((reg1342 ?
                          (8'haa) : wire1306) != reg1329)));
                end
            end
        end
    end
  assign wire1347 = "CyBVpyQYEP";
  always
    @(posedge clk) begin
      if ({{$unsigned(reg1312[(3'h4):(2'h3)])}})
        begin
          for (forvar1348 = (1'h0); (forvar1348 < (1'h0)); forvar1348 = (forvar1348 + (1'h1)))
            begin
              reg1349 = $signed(wire1301);
              reg1350 = reg1324[(4'h9):(3'h5)];
            end
        end
      else
        begin
          if (wire1347)
            begin
              if (wire1347)
                begin
                  for (forvar1348 = (1'h0); (forvar1348 < (2'h3)); forvar1348 = (forvar1348 + (1'h1)))
                    begin
                      reg1351 <= ((8'hb6) | $unsigned({(8'ha0)}));
                      reg1352 <= (8'hb4);
                    end
                  for (forvar1353 = (1'h0); (forvar1353 < (1'h1)); forvar1353 = (forvar1353 + (1'h1)))
                    begin
                      reg1354 <= reg1352[(4'ha):(2'h3)];
                      reg1355 = (($unsigned($unsigned(reg1351)) ^~ ((!wire1306) ?
                              ((8'had) ? reg1342 : reg1351) : {wire1305})) ?
                          reg1350[(3'h6):(2'h3)] : $signed(("mHw53A5OyrdfBd" ~^ {(8'ha8)})));
                      reg1356 = (~($unsigned($signed((8'ha3))) != (~|(reg1354 + (8'ha9)))));
                      reg1357 = $unsigned("miEQWplwJs");
                    end
                end
              else
                begin
                  reg1348 = "UAW0qdeAPpli8";
                  reg1349 = reg1323[(2'h3):(2'h2)];
                end
              for (forvar1358 = (1'h0); (forvar1358 < (1'h0)); forvar1358 = (forvar1358 + (1'h1)))
                begin
                  if ($signed($unsigned($signed(reg1350))))
                    begin
                      reg1359 <= wire1307[(1'h0):(1'h0)];
                      reg1360 = "kIdCLPTRcHHUfY";
                    end
                  else
                    begin
                      reg1359 <= (|($unsigned({reg1337}) >> {reg1348[(3'h6):(2'h3)]}));
                      reg1361 <= $unsigned($signed(reg1355));
                    end
                end
              reg1362 = forvar1358[(3'h6):(1'h0)];
            end
          else
            begin
              reg1351 <= $unsigned(reg1356[(2'h2):(2'h2)]);
              for (forvar1352 = (1'h0); (forvar1352 < (1'h1)); forvar1352 = (forvar1352 + (1'h1)))
                begin
                  reg1353 = $unsigned((8'ha2));
                  for (forvar1354 = (1'h0); (forvar1354 < (2'h3)); forvar1354 = (forvar1354 + (1'h1)))
                    begin
                      reg1358 <= $unsigned(("XE" ?
                          "s958HeJ6IXk7aP" : {$signed(wire1305)}));
                    end
                  reg1360 = (reg1319[(4'hf):(4'h9)] | (8'hac));
                  for (forvar1361 = (1'h0); (forvar1361 < (2'h2)); forvar1361 = (forvar1361 + (1'h1)))
                    begin
                      reg1363 <= ($signed(reg1319[(3'h4):(1'h0)]) != $signed(""));
                      reg1364 = $unsigned(reg1352[(4'h8):(3'h7)]);
                      reg1365 <= ((reg1332[(3'h4):(2'h2)] > $unsigned(reg1351[(2'h3):(2'h2)])) < $unsigned($unsigned((reg1312 ?
                          wire1302 : reg1323))));
                      reg1366 = ((~^$unsigned((|wire1303))) > (&(~&$unsigned(wire1302))));
                    end
                end
              reg1367 = (+reg1361[(4'hb):(1'h1)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg1368 <= ("56AV" && reg1324[(1'h0):(1'h0)]);
      reg1369 = wire1347;
      reg1370 = $signed((!((reg1323 ? reg1319 : reg1319) ?
          (reg1312 < reg1319) : $signed(wire1304))));
    end
  assign wire1371 = reg1354[(2'h3):(2'h3)];
  always
    @(posedge clk) begin
      for (forvar1372 = (1'h0); (forvar1372 < (1'h0)); forvar1372 = (forvar1372 + (1'h1)))
        begin
          for (forvar1373 = (1'h0); (forvar1373 < (2'h2)); forvar1373 = (forvar1373 + (1'h1)))
            begin
              reg1374 <= ((((~reg1312) <= reg1323) ?
                  ((forvar1372 ? reg1340 : (8'had)) ?
                      (forvar1373 && reg1354) : wire1305[(3'h5):(2'h3)]) : (|"NKH")) | $signed(({reg1361} | (^wire1305))));
              for (forvar1375 = (1'h0); (forvar1375 < (1'h1)); forvar1375 = (forvar1375 + (1'h1)))
                begin
                  for (forvar1376 = (1'h0); (forvar1376 < (2'h2)); forvar1376 = (forvar1376 + (1'h1)))
                    begin
                      reg1377 = reg1319;
                      reg1378 <= forvar1372[(4'h8):(1'h0)];
                      reg1379 = {(~(wire1303 ?
                              $unsigned(reg1354) : $signed(wire1303)))};
                    end
                  reg1380 = ((8'ha4) < $unsigned($unsigned((!reg1323))));
                end
              for (forvar1381 = (1'h0); (forvar1381 < (1'h1)); forvar1381 = (forvar1381 + (1'h1)))
                begin
                  for (forvar1382 = (1'h0); (forvar1382 < (1'h0)); forvar1382 = (forvar1382 + (1'h1)))
                    begin
                      reg1383 = reg1363;
                    end
                end
              for (forvar1384 = (1'h0); (forvar1384 < (2'h3)); forvar1384 = (forvar1384 + (1'h1)))
                begin
                  if ((8'hb9))
                    begin
                      reg1385 <= $unsigned($signed({$unsigned(forvar1372)}));
                      reg1386 = {$unsigned({(reg1324 <= reg1380)})};
                    end
                  else
                    begin
                      reg1386 = reg1337[(4'hf):(4'h9)];
                      reg1387 = ($unsigned(reg1359) > (~&((wire1347 & (8'hb9)) ?
                          reg1309 : reg1310[(3'h4):(1'h1)])));
                      reg1388 = "0MJNg7dcboPCtxH";
                    end
                  reg1389 = {{reg1337[(4'h9):(4'h9)]}};
                end
            end
        end
      reg1390 <= (!(8'hab));
      reg1391 <= {reg1378};
    end
  always
    @(posedge clk) begin
      if (((wire1304 - $signed((reg1368 ? reg1374 : reg1319))) ?
          (~^(((8'ha6) ? reg1332 : reg1358) ?
              wire1305[(1'h1):(1'h0)] : wire1303[(3'h7):(3'h4)])) : $unsigned($unsigned((|reg1315)))))
        begin
          for (forvar1392 = (1'h0); (forvar1392 < (2'h2)); forvar1392 = (forvar1392 + (1'h1)))
            begin
              if (reg1342)
                begin
                  reg1393 = (~&reg1323);
                  if ({((~^$signed(reg1363)) ?
                          reg1337[(3'h4):(3'h4)] : $unsigned((forvar1392 ?
                              reg1363 : (8'ha8))))})
                    begin
                      reg1394 = (&($unsigned({wire1371}) >= (^~(!wire1347))));
                    end
                  else
                    begin
                      reg1394 = ("WQx1k4xmMCc" ?
                          ($signed((reg1374 >>> reg1332)) || "d5kaatv6x") : (wire1302 > ((&(8'hb4)) ?
                              $signed(wire1301) : "qeCvwMskw76zYz4")));
                      reg1395 = $unsigned(($unsigned((&wire1347)) ?
                          $unsigned("VkviOq2eaatg2") : $signed((reg1315 >> reg1385))));
                      reg1396 <= "xqr9zZkUZt9W8";
                    end
                  for (forvar1397 = (1'h0); (forvar1397 < (2'h3)); forvar1397 = (forvar1397 + (1'h1)))
                    begin
                      reg1398 = (8'ha8);
                      reg1399 <= {(reg1390[(4'he):(3'h6)] ^~ (reg1374 ^~ "8xliQ8"))};
                      reg1400 <= $signed($unsigned(reg1339[(2'h3):(1'h1)]));
                      reg1401 <= "Ewc";
                    end
                  if ((reg1399[(3'h6):(3'h6)] ?
                      ($signed((8'ha5)) ?
                          (!(forvar1397 || reg1400)) : (reg1312 ?
                              (8'hba) : (reg1390 < wire1301))) : {$signed(((8'hac) & reg1332))}))
                    begin
                      reg1402 = (($unsigned((forvar1397 ?
                          wire1371 : reg1315)) < reg1401[(1'h1):(1'h0)]) >= "ZsNG");
                      reg1403 = (forvar1397 * $signed($unsigned("LVb")));
                    end
                  else
                    begin
                      reg1404 <= "UytPhpnt6";
                    end
                end
              else
                begin
                  reg1393 = reg1312;
                  reg1394 = "bB474i";
                end
              reg1405 = (reg1378 ?
                  $unsigned(reg1398[(1'h0):(1'h0)]) : ({$unsigned((8'hb5))} ?
                      {reg1354} : $unsigned($signed((8'haf)))));
              reg1406 <= wire1306[(1'h0):(1'h0)];
            end
          reg1407 = reg1398;
        end
      else
        begin
          for (forvar1392 = (1'h0); (forvar1392 < (2'h2)); forvar1392 = (forvar1392 + (1'h1)))
            begin
              if ("SmqnFkaq0wd9kX")
                begin
                  for (forvar1393 = (1'h0); (forvar1393 < (1'h1)); forvar1393 = (forvar1393 + (1'h1)))
                    begin
                      reg1394 = (+"mapXxtEPvah");
                      reg1396 <= (~|(reg1399 ?
                          ((|reg1323) == (reg1406 ?
                              reg1339 : (8'ha0))) : $signed(reg1339)));
                      reg1397 = $unsigned({(~|$signed(reg1394))});
                    end
                  reg1398 = $signed("0dJZKa4Wf4QK");
                end
              else
                begin
                  for (forvar1393 = (1'h0); (forvar1393 < (2'h3)); forvar1393 = (forvar1393 + (1'h1)))
                    begin
                      reg1396 <= $unsigned((((|reg1368) ^ "bshCOeQs4AumV") ?
                          (reg1394 ?
                              $unsigned(reg1354) : (!reg1315)) : {reg1319[(4'hf):(3'h4)]}));
                      reg1397 = {{(!$unsigned(wire1303))}};
                      reg1399 <= ($signed($unsigned({wire1347})) >> $signed(reg1354));
                      reg1400 <= $unsigned(((&reg1405) < (~^$signed((8'hb6)))));
                    end
                  reg1402 = wire1371[(1'h1):(1'h1)];
                  reg1403 = {(({reg1396} ? $unsigned(reg1358) : {wire1306}) ?
                          reg1398[(2'h3):(2'h3)] : $signed((reg1312 != reg1394)))};
                end
            end
        end
      reg1408 = (8'hb1);
      for (forvar1409 = (1'h0); (forvar1409 < (2'h3)); forvar1409 = (forvar1409 + (1'h1)))
        begin
          for (forvar1410 = (1'h0); (forvar1410 < (1'h0)); forvar1410 = (forvar1410 + (1'h1)))
            begin
              if ((~&$unsigned(wire1304)))
                begin
                  reg1411 = reg1315;
                  reg1412 <= ($signed((|reg1363[(1'h0):(1'h0)])) > (!wire1347));
                end
              else
                begin
                  for (forvar1411 = (1'h0); (forvar1411 < (1'h0)); forvar1411 = (forvar1411 + (1'h1)))
                    begin
                      reg1413 = ($unsigned((((8'hb2) ?
                              (8'hb2) : wire1304) && (reg1339 ~^ reg1332))) ?
                          "" : reg1396[(2'h2):(1'h0)]);
                      reg1414 = $signed(reg1319);
                      reg1415 <= (reg1402[(3'h6):(3'h5)] * (~^$unsigned(reg1337[(3'h5):(1'h0)])));
                    end
                  for (forvar1416 = (1'h0); (forvar1416 < (1'h1)); forvar1416 = (forvar1416 + (1'h1)))
                    begin
                      reg1417 = $unsigned({{$unsigned(reg1385)}});
                      reg1418 <= $unsigned({(^~$signed(reg1339))});
                      reg1419 = ($unsigned(($signed(reg1358) ?
                              $unsigned(reg1401) : $signed(reg1400))) ?
                          $signed(((8'h9c) >> {forvar1393})) : (8'ha0));
                      reg1420 = $unsigned((reg1406[(3'h4):(2'h2)] ^ $signed($unsigned(forvar1409))));
                    end
                  reg1421 <= wire1307[(1'h1):(1'h0)];
                end
              reg1422 = reg1339[(3'h6):(3'h6)];
              if ($signed({$signed($signed(forvar1392))}))
                begin
                  reg1423 <= (!({wire1306[(2'h2):(1'h0)]} ?
                      ((reg1361 + reg1395) & (reg1327 ?
                          reg1413 : wire1302)) : {"3htY7XtGlzavk"}));
                  reg1424 = (^~(8'hb2));
                end
              else
                begin
                  for (forvar1423 = (1'h0); (forvar1423 < (1'h0)); forvar1423 = (forvar1423 + (1'h1)))
                    begin
                      reg1424 = $unsigned(reg1354[(4'hf):(4'hf)]);
                      reg1425 = ((|{{reg1315}}) ?
                          $unsigned({$signed(reg1309)}) : reg1411);
                    end
                  for (forvar1426 = (1'h0); (forvar1426 < (1'h0)); forvar1426 = (forvar1426 + (1'h1)))
                    begin
                      reg1427 = "4Po";
                    end
                  if (($signed($signed($signed(reg1397))) ?
                      wire1306[(1'h1):(1'h1)] : (~^{"kNAG"})))
                    begin
                      reg1428 = $signed(("GJd384aKUPr" * ((wire1307 ^ wire1371) ?
                          (reg1339 & reg1398) : forvar1423)));
                      reg1429 = (~&reg1374[(4'h9):(3'h7)]);
                      reg1430 <= reg1394;
                    end
                  else
                    begin
                      reg1428 = reg1354;
                    end
                  for (forvar1431 = (1'h0); (forvar1431 < (1'h1)); forvar1431 = (forvar1431 + (1'h1)))
                    begin
                      reg1432 <= ((8'hb0) + {$signed(((8'h9d) ?
                              reg1407 : (8'hb0)))});
                      reg1433 = ($unsigned(reg1419[(2'h2):(1'h0)]) ?
                          ($signed((forvar1409 << reg1327)) | "XJCHT") : (((8'ha3) ?
                              "9Ug2k8" : (+reg1413)) <<< $unsigned((^(8'hab)))));
                      reg1434 = reg1411;
                      reg1435 = (reg1351 ?
                          "o1Dsban" : $unsigned(reg1433[(1'h0):(1'h0)]));
                    end
                end
            end
          reg1436 <= $signed((!reg1413[(1'h0):(1'h0)]));
        end
      if (("DloJTsLOZ" ? (reg1363 <<< "75i1") : reg1436))
        begin
          reg1437 = {$signed((8'ha0))};
          for (forvar1438 = (1'h0); (forvar1438 < (2'h3)); forvar1438 = (forvar1438 + (1'h1)))
            begin
              for (forvar1439 = (1'h0); (forvar1439 < (2'h2)); forvar1439 = (forvar1439 + (1'h1)))
                begin
                  for (forvar1440 = (1'h0); (forvar1440 < (1'h1)); forvar1440 = (forvar1440 + (1'h1)))
                    begin
                      reg1441 = reg1342[(4'hd):(2'h2)];
                      reg1442 = ({$signed($signed((8'ha0)))} - ($signed((reg1441 ?
                          reg1368 : (8'hb3))) + $signed(reg1411)));
                      reg1443 = reg1406;
                      reg1444 <= $unsigned(($unsigned(((8'hb2) ^ reg1396)) ?
                          "hzvwDCEd1v" : reg1407));
                    end
                  reg1445 = $signed((($unsigned((8'hb4)) ^~ $signed(reg1324)) ?
                      reg1419[(1'h1):(1'h1)] : (^"FOa20Rg8WVAR")));
                  for (forvar1446 = (1'h0); (forvar1446 < (2'h2)); forvar1446 = (forvar1446 + (1'h1)))
                    begin
                      reg1447 <= $signed({((~reg1411) - $signed(reg1390))});
                      reg1448 = forvar1416;
                      reg1449 = forvar1416;
                      reg1450 = $unsigned($signed(forvar1397));
                    end
                end
              for (forvar1451 = (1'h0); (forvar1451 < (1'h0)); forvar1451 = (forvar1451 + (1'h1)))
                begin
                  for (forvar1452 = (1'h0); (forvar1452 < (2'h2)); forvar1452 = (forvar1452 + (1'h1)))
                    begin
                      reg1453 <= {$signed((~|(+reg1449)))};
                      reg1454 = reg1450[(1'h1):(1'h1)];
                      reg1455 = $unsigned($unsigned(reg1324));
                      reg1456 = reg1408;
                    end
                  for (forvar1457 = (1'h0); (forvar1457 < (2'h2)); forvar1457 = (forvar1457 + (1'h1)))
                    begin
                      reg1458 = reg1312[(2'h3):(2'h2)];
                      reg1459 = ((~|{(reg1414 <<< reg1448)}) < ($unsigned(forvar1411) ?
                          ((reg1404 ?
                              reg1361 : (8'hb7)) > reg1397) : {{(8'ha0)}}));
                      reg1460 <= wire1303[(4'h9):(2'h2)];
                      reg1461 = ("LVcQ" == (reg1415 & ((forvar1451 <= forvar1397) != reg1453[(2'h3):(2'h3)])));
                    end
                  reg1462 = {(8'hae)};
                  reg1463 = "nQ8RDSo";
                end
            end
        end
      else
        begin
          reg1438 <= reg1403[(2'h3):(1'h1)];
          if ({$signed($signed(reg1339))})
            begin
              if (reg1352)
                begin
                  for (forvar1439 = (1'h0); (forvar1439 < (2'h3)); forvar1439 = (forvar1439 + (1'h1)))
                    begin
                      reg1440 = ((forvar1438 ?
                          ((-forvar1392) ?
                              reg1401[(2'h2):(2'h2)] : reg1453) : ($signed(reg1332) & {reg1395})) - forvar1397[(1'h1):(1'h1)]);
                      reg1444 <= {($signed(forvar1452[(1'h1):(1'h1)]) ?
                              "4Aszs7GeHKqKMX4" : "N8TOI")};
                    end
                end
              else
                begin
                  reg1439 = (forvar1409 ?
                      $signed(wire1371[(1'h1):(1'h1)]) : $unsigned((reg1441[(1'h0):(1'h0)] ?
                          forvar1446[(3'h7):(1'h0)] : (+reg1428))));
                end
              for (forvar1445 = (1'h0); (forvar1445 < (1'h1)); forvar1445 = (forvar1445 + (1'h1)))
                begin
                  for (forvar1446 = (1'h0); (forvar1446 < (2'h2)); forvar1446 = (forvar1446 + (1'h1)))
                    begin
                      reg1447 <= $signed("Tkwtk5MI");
                      reg1448 = reg1433[(1'h1):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar1439 = (1'h0); (forvar1439 < (2'h3)); forvar1439 = (forvar1439 + (1'h1)))
                begin
                  if ("QxNTssP")
                    begin
                      reg1440 = wire1307[(2'h2):(1'h1)];
                      reg1441 = $unsigned((~&(|(+forvar1426))));
                      reg1444 <= {(8'h9c)};
                    end
                  else
                    begin
                      reg1444 <= ((~^(~|forvar1438)) ?
                          reg1450 : ("x1ugbr8nd" && (|reg1342[(2'h3):(1'h1)])));
                      reg1445 = {(~$signed((reg1418 ? reg1437 : reg1450)))};
                    end
                  if ($signed($signed(reg1448[(4'h8):(3'h5)])))
                    begin
                      reg1446 = $unsigned(($unsigned((reg1385 || reg1418)) ?
                          $signed(reg1458[(4'hf):(4'hd)]) : "GWUHI71EtxXv"));
                      reg1448 = $unsigned(reg1403);
                      reg1449 = $signed("QglQ9CwY");
                    end
                  else
                    begin
                      reg1447 <= reg1436;
                    end
                  reg1450 = $unsigned(((!reg1390) ?
                      $unsigned(reg1461[(4'h8):(2'h3)]) : forvar1446[(1'h1):(1'h0)]));
                  for (forvar1451 = (1'h0); (forvar1451 < (1'h1)); forvar1451 = (forvar1451 + (1'h1)))
                    begin
                      reg1452 = (~&($unsigned($signed(reg1365)) ^ (|$unsigned((8'hb5)))));
                      reg1453 <= (&reg1440[(2'h2):(2'h2)]);
                    end
                end
              reg1454 = (reg1454[(1'h0):(1'h0)] == (($signed(reg1455) >= reg1455) ?
                  wire1303 : (~reg1444[(2'h2):(1'h1)])));
              reg1455 = reg1414[(3'h5):(3'h5)];
            end
          if (($unsigned(((+forvar1410) || {reg1453})) <= reg1450))
            begin
              reg1456 = $unsigned({$unsigned($unsigned(reg1452))});
              for (forvar1457 = (1'h0); (forvar1457 < (2'h2)); forvar1457 = (forvar1457 + (1'h1)))
                begin
                  for (forvar1458 = (1'h0); (forvar1458 < (1'h0)); forvar1458 = (forvar1458 + (1'h1)))
                    begin
                      reg1459 = "4SkycWVF";
                    end
                  reg1461 = $signed(reg1446);
                end
            end
          else
            begin
              for (forvar1456 = (1'h0); (forvar1456 < (1'h0)); forvar1456 = (forvar1456 + (1'h1)))
                begin
                  if (($signed(($signed(reg1391) - (^~reg1361))) ?
                      reg1340 : ($unsigned((reg1327 ?
                          (8'h9f) : reg1436)) && (~|"NIksahVUfz70"))))
                    begin
                      reg1457 <= (|forvar1426[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg1458 = $signed(forvar1438);
                    end
                  if (($signed($unsigned("lQK4B2UJ")) ^ ($unsigned($signed(forvar1397)) >>> ($unsigned(forvar1457) ?
                      ((8'had) << reg1363) : reg1457[(1'h1):(1'h1)]))))
                    begin
                      reg1459 = (reg1390 | reg1455[(4'hc):(2'h2)]);
                    end
                  else
                    begin
                      reg1459 = reg1428[(4'hc):(3'h5)];
                      reg1460 <= $unsigned(((reg1460[(2'h3):(1'h1)] ^ $unsigned(reg1352)) | (~^$signed((8'hb4)))));
                      reg1461 = "n1DIMZxZLlUR1";
                      reg1462 = $unsigned(((-{reg1448}) ^~ (~&$signed(reg1428))));
                    end
                  for (forvar1463 = (1'h0); (forvar1463 < (2'h2)); forvar1463 = (forvar1463 + (1'h1)))
                    begin
                      reg1464 = $signed(reg1323[(4'h8):(1'h0)]);
                      reg1465 = $unsigned($unsigned($signed((reg1407 ?
                          (8'ha7) : reg1417))));
                      reg1466 = (~|reg1352);
                      reg1467 <= reg1323[(4'ha):(2'h3)];
                    end
                end
            end
          if ($signed($signed($signed({reg1447}))))
            begin
              for (forvar1468 = (1'h0); (forvar1468 < (2'h2)); forvar1468 = (forvar1468 + (1'h1)))
                begin
                  for (forvar1469 = (1'h0); (forvar1469 < (2'h2)); forvar1469 = (forvar1469 + (1'h1)))
                    begin
                      reg1470 = ("5Y1" * $signed($unsigned(reg1433[(2'h2):(2'h2)])));
                    end
                end
              if ((~^(({reg1327} >= (reg1457 - reg1399)) || $signed(reg1407))))
                begin
                  for (forvar1471 = (1'h0); (forvar1471 < (2'h3)); forvar1471 = (forvar1471 + (1'h1)))
                    begin
                      reg1472 = (&{$unsigned($signed(reg1400))});
                    end
                  reg1473 = (~^($unsigned(forvar1471) || reg1434));
                  if ((($signed((reg1324 <= (8'ha2))) ?
                          $signed((reg1441 + reg1455)) : ((reg1462 ?
                              forvar1423 : reg1432) >>> $signed(reg1401))) ?
                      (8'h9e) : $signed($unsigned((reg1437 ?
                          reg1319 : reg1394)))))
                    begin
                      reg1474 <= ((~^$unsigned((^~reg1342))) < reg1465[(2'h3):(1'h0)]);
                      reg1475 = forvar1416[(3'h7):(1'h0)];
                      reg1476 = {("wP9Xvamv" ?
                              (^~reg1430[(1'h0):(1'h0)]) : reg1417[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg1474 <= (8'hb8);
                      reg1475 = forvar1457;
                    end
                end
              else
                begin
                  reg1471 = (reg1401[(2'h2):(1'h1)] ?
                      $signed($signed($signed((8'hb7)))) : ($unsigned($unsigned(reg1358)) - $signed((reg1415 | reg1475))));
                  reg1472 = reg1467[(3'h5):(1'h0)];
                  for (forvar1473 = (1'h0); (forvar1473 < (1'h1)); forvar1473 = (forvar1473 + (1'h1)))
                    begin
                      reg1475 = (reg1438 != $unsigned((!(wire1347 > forvar1468))));
                    end
                  reg1476 = reg1475[(2'h2):(1'h1)];
                end
            end
          else
            begin
              for (forvar1468 = (1'h0); (forvar1468 < (1'h0)); forvar1468 = (forvar1468 + (1'h1)))
                begin
                  for (forvar1469 = (1'h0); (forvar1469 < (1'h0)); forvar1469 = (forvar1469 + (1'h1)))
                    begin
                      reg1474 <= (^~(reg1385[(3'h4):(2'h3)] + ($signed(reg1441) >= "kd3PQ")));
                    end
                  for (forvar1475 = (1'h0); (forvar1475 < (1'h0)); forvar1475 = (forvar1475 + (1'h1)))
                    begin
                      reg1477 <= "SEmfBU";
                      reg1478 = {$unsigned({(reg1446 ? reg1407 : reg1352)})};
                      reg1479 <= (reg1478 <<< forvar1458);
                    end
                  for (forvar1480 = (1'h0); (forvar1480 < (2'h2)); forvar1480 = (forvar1480 + (1'h1)))
                    begin
                      reg1481 = {{reg1446[(4'hc):(1'h0)]}};
                    end
                  for (forvar1482 = (1'h0); (forvar1482 < (2'h2)); forvar1482 = (forvar1482 + (1'h1)))
                    begin
                      reg1483 = {wire1347[(4'hb):(4'h8)]};
                      reg1484 = reg1434;
                    end
                end
              for (forvar1485 = (1'h0); (forvar1485 < (1'h0)); forvar1485 = (forvar1485 + (1'h1)))
                begin
                  if (({((forvar1397 + forvar1409) - {wire1301})} ?
                      $signed(((reg1432 >> reg1414) ?
                          reg1481 : (reg1473 ?
                              reg1393 : reg1359))) : (reg1406[(3'h5):(1'h1)] * $signed($unsigned(reg1363)))))
                    begin
                      reg1486 = reg1459;
                      reg1487 = $unsigned((reg1419[(3'h4):(2'h3)] <<< $unsigned(((8'haa) >> reg1449))));
                      reg1488 = reg1452;
                    end
                  else
                    begin
                      reg1486 = (~&$unsigned((~^reg1351)));
                      reg1489 <= ("1HXB0ct3mc48" ?
                          $unsigned(((~(8'ha6)) ?
                              reg1319[(3'h4):(2'h3)] : reg1358)) : ($unsigned($signed((8'hab))) ^~ ($signed((8'ha1)) + $unsigned(reg1374))));
                      reg1490 <= "Yz9W";
                    end
                  if ($signed($signed($unsigned((reg1457 ?
                      (8'ha5) : wire1301)))))
                    begin
                      reg1491 = reg1403[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg1492 <= forvar1440;
                      reg1493 = $signed($signed({(~&reg1458)}));
                    end
                  for (forvar1494 = (1'h0); (forvar1494 < (1'h0)); forvar1494 = (forvar1494 + (1'h1)))
                    begin
                      reg1495 = ($unsigned(wire1304) ?
                          (reg1422[(2'h2):(1'h1)] >>> (forvar1480 ?
                              $unsigned(reg1474) : "hCLBrVGxke")) : (~&$unsigned($unsigned(reg1432))));
                    end
                end
            end
        end
    end
  assign wire1496 = reg1310;
  assign wire1497 = $signed((^$signed((reg1361 ? wire1301 : (8'ha5)))));
  assign wire1498 = reg1490[(3'h5):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar1499 = (1'h0); (forvar1499 < (2'h2)); forvar1499 = (forvar1499 + (1'h1)))
        begin
          for (forvar1500 = (1'h0); (forvar1500 < (2'h3)); forvar1500 = (forvar1500 + (1'h1)))
            begin
              reg1501 = $signed((8'hb9));
              for (forvar1502 = (1'h0); (forvar1502 < (2'h3)); forvar1502 = (forvar1502 + (1'h1)))
                begin
                  reg1503 <= reg1312;
                  for (forvar1504 = (1'h0); (forvar1504 < (1'h1)); forvar1504 = (forvar1504 + (1'h1)))
                    begin
                      reg1505 <= (+$unsigned({reg1368}));
                      reg1506 <= reg1492;
                      reg1507 = {(wire1303 != reg1319)};
                      reg1508 = reg1312;
                    end
                end
              for (forvar1509 = (1'h0); (forvar1509 < (2'h2)); forvar1509 = (forvar1509 + (1'h1)))
                begin
                  for (forvar1510 = (1'h0); (forvar1510 < (1'h1)); forvar1510 = (forvar1510 + (1'h1)))
                    begin
                      reg1511 <= reg1436[(3'h7):(1'h0)];
                    end
                  for (forvar1512 = (1'h0); (forvar1512 < (2'h2)); forvar1512 = (forvar1512 + (1'h1)))
                    begin
                      reg1513 <= $signed("LXWXcIH6QeaoJaf");
                      reg1514 = (~|(~("qA" & $signed(reg1354))));
                    end
                end
            end
          for (forvar1515 = (1'h0); (forvar1515 < (2'h2)); forvar1515 = (forvar1515 + (1'h1)))
            begin
              if (($signed((8'hb7)) ? (~|(-reg1506)) : ""))
                begin
                  reg1516 = wire1305;
                  if ($unsigned($signed({{reg1514}})))
                    begin
                      reg1517 = ("xZYCA6p9ky2f" ?
                          $signed(reg1516[(2'h3):(1'h1)]) : ("1" ^~ reg1516));
                    end
                  else
                    begin
                      reg1517 = ((~^$unsigned(reg1453[(1'h1):(1'h0)])) | ((~&(&(8'h9d))) && ("WNY" ?
                          "bk" : reg1399[(4'ha):(4'h8)])));
                      reg1518 = reg1489[(3'h5):(2'h3)];
                      reg1519 <= (8'ha5);
                    end
                  if (wire1302)
                    begin
                      reg1520 <= {((~reg1351[(2'h2):(1'h1)]) ?
                              ((forvar1512 ~^ (8'h9f)) <<< wire1498) : $unsigned((^~(8'ha5))))};
                    end
                  else
                    begin
                      reg1520 <= (((reg1310[(2'h3):(1'h1)] << $unsigned((8'hb8))) * {(|(8'hb7))}) - wire1304[(4'hd):(3'h6)]);
                      reg1521 <= $unsigned((+(|(~&reg1332))));
                      reg1522 = ((~&"xTA2h1WYI") ?
                          reg1323[(3'h6):(3'h4)] : $signed(((reg1518 != reg1385) + $unsigned(reg1324))));
                    end
                  if ({((~|(8'h9c)) && reg1327[(4'h9):(2'h3)])})
                    begin
                      reg1523 = ((8'ha8) != "Tr9xcTdYob");
                      reg1524 = $signed((^$unsigned($signed(reg1522))));
                    end
                  else
                    begin
                      reg1523 = (-reg1516);
                      reg1524 = reg1310[(4'hb):(4'h9)];
                      reg1525 = reg1352;
                    end
                end
              else
                begin
                  for (forvar1516 = (1'h0); (forvar1516 < (2'h3)); forvar1516 = (forvar1516 + (1'h1)))
                    begin
                      reg1519 <= ($unsigned((~&$unsigned((8'ha8)))) & (reg1490 ?
                          reg1412[(3'h5):(1'h0)] : wire1304[(4'hc):(4'h9)]));
                      reg1522 = {(~$signed(reg1489))};
                      reg1526 <= wire1305;
                    end
                  for (forvar1527 = (1'h0); (forvar1527 < (1'h0)); forvar1527 = (forvar1527 + (1'h1)))
                    begin
                      reg1528 = reg1415;
                      reg1529 = (^~$unsigned((^{reg1368})));
                      reg1530 <= ((reg1517 ?
                          reg1374[(4'h9):(2'h2)] : $signed(reg1342)) * reg1342);
                    end
                  for (forvar1531 = (1'h0); (forvar1531 < (2'h3)); forvar1531 = (forvar1531 + (1'h1)))
                    begin
                      reg1532 <= $unsigned($unsigned(((reg1444 >> wire1302) << {forvar1502})));
                    end
                  for (forvar1533 = (1'h0); (forvar1533 < (2'h3)); forvar1533 = (forvar1533 + (1'h1)))
                    begin
                      reg1534 = (~({(-reg1516)} ?
                          $unsigned((forvar1499 <= reg1351)) : reg1368[(1'h0):(1'h0)]));
                      reg1535 <= $signed($signed($unsigned((wire1307 ?
                          reg1514 : (8'ha2)))));
                      reg1536 = $unsigned({(+(reg1390 * reg1535))});
                    end
                end
            end
          reg1537 = ((((reg1457 ? reg1518 : forvar1499) ?
                  ((8'h9f) ? (8'ha9) : reg1339) : ((8'hb2) ?
                      (8'ha4) : reg1479)) <= "93RS") ?
              reg1529 : (~&((reg1529 != reg1525) ? wire1307 : "kokWuK9Xx")));
        end
    end
endmodule