(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'he4d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire0;
  input wire signed [(4'hb):(1'h0)] wire1;
  input wire signed [(4'he):(1'h0)] wire2;
  input wire signed [(4'h8):(1'h0)] wire3;
  input wire signed [(3'h6):(1'h0)] wire4;
  wire [(4'h9):(1'h0)] wire1906;
  wire signed [(3'h7):(1'h0)] wire1905;
  wire [(4'hf):(1'h0)] wire1904;
  wire [(2'h2):(1'h0)] wire1903;
  wire [(4'h9):(1'h0)] wire1902;
  wire signed [(3'h6):(1'h0)] wire1822;
  wire [(3'h7):(1'h0)] wire1821;
  wire signed [(3'h7):(1'h0)] wire1753;
  wire [(3'h6):(1'h0)] wire1088;
  wire signed [(3'h5):(1'h0)] wire1086;
  wire signed [(4'he):(1'h0)] wire632;
  wire [(4'h9):(1'h0)] wire631;
  wire [(3'h7):(1'h0)] wire629;
  reg [(3'h5):(1'h0)] reg1901 = (1'h0);
  reg [(4'hf):(1'h0)] reg1900 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1899 = (1'h0);
  reg [(4'ha):(1'h0)] reg1898 = (1'h0);
  reg [(3'h4):(1'h0)] reg1897 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1896 = (1'h0);
  reg [(2'h2):(1'h0)] reg1895 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1893 = (1'h0);
  reg [(4'hb):(1'h0)] reg1891 = (1'h0);
  reg [(4'h9):(1'h0)] reg1889 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1887 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1886 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1885 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1884 = (1'h0);
  reg [(3'h6):(1'h0)] reg1823 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1879 = (1'h0);
  reg [(4'h8):(1'h0)] reg1878 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1877 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1876 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1875 = (1'h0);
  reg [(3'h6):(1'h0)] reg1874 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1873 = (1'h0);
  reg [(3'h7):(1'h0)] reg1872 = (1'h0);
  reg [(4'hb):(1'h0)] reg1871 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1869 = (1'h0);
  reg [(3'h4):(1'h0)] reg1868 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1867 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1866 = (1'h0);
  reg [(4'ha):(1'h0)] reg1865 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1863 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1862 = (1'h0);
  reg [(4'hd):(1'h0)] reg1861 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1860 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1859 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1858 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1857 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1855 = (1'h0);
  reg [(4'h9):(1'h0)] reg1856 = (1'h0);
  reg [(4'he):(1'h0)] reg1854 = (1'h0);
  reg [(5'h10):(1'h0)] reg1853 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1852 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1851 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1849 = (1'h0);
  reg [(4'ha):(1'h0)] reg1848 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1846 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1845 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1844 = (1'h0);
  reg [(3'h5):(1'h0)] reg1842 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1841 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1840 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1828 = (1'h0);
  reg [(4'h9):(1'h0)] reg1838 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1837 = (1'h0);
  reg [(4'hd):(1'h0)] reg1836 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1835 = (1'h0);
  reg [(3'h5):(1'h0)] reg1834 = (1'h0);
  reg [(4'hc):(1'h0)] reg1832 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1831 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1830 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1829 = (1'h0);
  reg [(3'h4):(1'h0)] reg1827 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1826 = (1'h0);
  reg [(4'ha):(1'h0)] reg1825 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1824 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1820 = (1'h0);
  reg [(4'hf):(1'h0)] reg1819 = (1'h0);
  reg [(3'h5):(1'h0)] reg1818 = (1'h0);
  reg [(4'h9):(1'h0)] reg1816 = (1'h0);
  reg [(4'hc):(1'h0)] reg1815 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1814 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1811 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1809 = (1'h0);
  reg [(3'h4):(1'h0)] reg1808 = (1'h0);
  reg [(3'h7):(1'h0)] reg1807 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1806 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1805 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1804 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1803 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1801 = (1'h0);
  reg [(4'ha):(1'h0)] reg1799 = (1'h0);
  reg [(4'h9):(1'h0)] reg1798 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1796 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1795 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1794 = (1'h0);
  reg [(4'hf):(1'h0)] reg1793 = (1'h0);
  reg [(2'h2):(1'h0)] reg1792 = (1'h0);
  reg [(4'he):(1'h0)] reg1791 = (1'h0);
  reg [(3'h7):(1'h0)] reg1789 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1788 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1787 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1785 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1784 = (1'h0);
  reg [(3'h4):(1'h0)] reg1783 = (1'h0);
  reg [(4'hc):(1'h0)] reg1782 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1781 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1780 = (1'h0);
  reg [(5'h10):(1'h0)] reg1779 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1778 = (1'h0);
  reg [(4'h8):(1'h0)] reg1777 = (1'h0);
  reg [(3'h7):(1'h0)] reg1776 = (1'h0);
  reg [(4'h8):(1'h0)] reg1768 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1759 = (1'h0);
  reg [(2'h2):(1'h0)] reg1775 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1774 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1773 = (1'h0);
  reg [(3'h7):(1'h0)] reg1772 = (1'h0);
  reg [(3'h5):(1'h0)] reg1771 = (1'h0);
  reg [(3'h5):(1'h0)] reg1762 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1770 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1769 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1767 = (1'h0);
  reg [(4'ha):(1'h0)] reg1766 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1765 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1764 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1763 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1761 = (1'h0);
  reg [(4'hc):(1'h0)] reg1760 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1758 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1757 = (1'h0);
  reg [(4'h8):(1'h0)] reg635 = (1'h0);
  reg [(4'hc):(1'h0)] reg636 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg638 = (1'h0);
  reg [(5'h10):(1'h0)] reg639 = (1'h0);
  reg [(4'he):(1'h0)] reg640 = (1'h0);
  reg [(4'hf):(1'h0)] reg641 = (1'h0);
  reg [(3'h5):(1'h0)] reg644 = (1'h0);
  reg [(3'h4):(1'h0)] reg645 = (1'h0);
  reg [(3'h4):(1'h0)] reg646 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg648 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg649 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg652 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg653 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg654 = (1'h0);
  reg [(4'h9):(1'h0)] reg655 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg656 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg657 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg658 = (1'h0);
  reg [(2'h2):(1'h0)] reg660 = (1'h0);
  reg [(4'h9):(1'h0)] reg661 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg662 = (1'h0);
  reg [(4'hc):(1'h0)] reg664 = (1'h0);
  reg [(4'hd):(1'h0)] reg665 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg666 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg634 = (1'h0);
  reg [(3'h7):(1'h0)] reg637 = (1'h0);
  reg signed [(4'he):(1'h0)] reg643 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg647 = (1'h0);
  reg [(4'hb):(1'h0)] reg650 = (1'h0);
  reg signed [(4'he):(1'h0)] reg651 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg659 = (1'h0);
  reg [(3'h7):(1'h0)] reg642 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg663 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg667 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg668 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg669 = (1'h0);
  reg [(4'hf):(1'h0)] reg670 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg671 = (1'h0);
  reg [(4'hf):(1'h0)] reg674 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg675 = (1'h0);
  reg [(2'h3):(1'h0)] reg676 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg677 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg678 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg679 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg680 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg681 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg683 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg684 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg685 = (1'h0);
  reg [(3'h5):(1'h0)] reg687 = (1'h0);
  reg [(2'h2):(1'h0)] reg688 = (1'h0);
  reg [(4'hf):(1'h0)] reg689 = (1'h0);
  reg [(2'h2):(1'h0)] reg691 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg692 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg693 = (1'h0);
  reg [(4'hd):(1'h0)] reg694 = (1'h0);
  reg [(4'h8):(1'h0)] reg695 = (1'h0);
  reg [(4'hb):(1'h0)] reg697 = (1'h0);
  reg signed [(4'he):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg699 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg702 = (1'h0);
  reg signed [(4'he):(1'h0)] reg704 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg705 = (1'h0);
  reg [(3'h4):(1'h0)] reg706 = (1'h0);
  reg [(3'h6):(1'h0)] reg707 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg708 = (1'h0);
  reg [(3'h5):(1'h0)] reg711 = (1'h0);
  reg [(4'hf):(1'h0)] reg712 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg713 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg714 = (1'h0);
  reg [(4'ha):(1'h0)] reg715 = (1'h0);
  reg [(5'h10):(1'h0)] reg716 = (1'h0);
  reg [(3'h7):(1'h0)] reg717 = (1'h0);
  reg [(3'h4):(1'h0)] reg718 = (1'h0);
  reg [(4'h8):(1'h0)] reg690 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg720 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg721 = (1'h0);
  reg [(4'ha):(1'h0)] reg724 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg726 = (1'h0);
  reg [(5'h10):(1'h0)] reg727 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg728 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg729 = (1'h0);
  reg [(3'h4):(1'h0)] reg701 = (1'h0);
  reg [(4'he):(1'h0)] reg703 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg709 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg696 = (1'h0);
  reg [(3'h6):(1'h0)] reg719 = (1'h0);
  reg [(2'h3):(1'h0)] reg722 = (1'h0);
  reg [(2'h2):(1'h0)] reg723 = (1'h0);
  reg [(4'h9):(1'h0)] reg725 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg730 = (1'h0);
  reg [(2'h2):(1'h0)] reg731 = (1'h0);
  reg [(4'ha):(1'h0)] reg732 = (1'h0);
  reg [(4'he):(1'h0)] reg733 = (1'h0);
  reg [(4'h8):(1'h0)] reg734 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg736 = (1'h0);
  reg [(4'hd):(1'h0)] reg737 = (1'h0);
  reg [(4'hf):(1'h0)] reg738 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1089 = (1'h0);
  reg [(4'hc):(1'h0)] reg1090 = (1'h0);
  reg [(4'hd):(1'h0)] reg1092 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1093 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1095 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1096 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1097 = (1'h0);
  reg [(4'hc):(1'h0)] reg1098 = (1'h0);
  reg [(5'h10):(1'h0)] reg1100 = (1'h0);
  reg [(5'h10):(1'h0)] reg1091 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1094 = (1'h0);
  reg [(4'hd):(1'h0)] reg1099 = (1'h0);
  reg [(4'hf):(1'h0)] reg1101 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1102 = (1'h0);
  reg [(3'h5):(1'h0)] reg1103 = (1'h0);
  reg [(2'h2):(1'h0)] reg1104 = (1'h0);
  reg [(4'hb):(1'h0)] reg1105 = (1'h0);
  reg [(5'h10):(1'h0)] reg1106 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1107 = (1'h0);
  reg [(4'he):(1'h0)] reg1108 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1109 = (1'h0);
  reg [(4'h8):(1'h0)] reg1110 = (1'h0);
  reg [(4'hf):(1'h0)] reg1111 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1112 = (1'h0);
  reg [(3'h4):(1'h0)] reg1113 = (1'h0);
  reg [(4'hb):(1'h0)] reg1114 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1116 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1117 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1118 = (1'h0);
  reg [(3'h7):(1'h0)] reg1119 = (1'h0);
  reg [(4'h8):(1'h0)] reg1121 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1122 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1123 = (1'h0);
  reg [(2'h2):(1'h0)] reg1124 = (1'h0);
  reg [(5'h10):(1'h0)] reg1125 = (1'h0);
  reg [(3'h6):(1'h0)] reg1126 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1120 = (1'h0);
  reg [(4'hb):(1'h0)] reg1127 = (1'h0);
  reg [(4'he):(1'h0)] reg1115 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1128 = (1'h0);
  reg [(4'he):(1'h0)] reg1130 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1131 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1132 = (1'h0);
  reg [(4'h8):(1'h0)] reg1134 = (1'h0);
  reg [(4'he):(1'h0)] reg1135 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1136 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1140 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1142 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1143 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1144 = (1'h0);
  reg [(2'h2):(1'h0)] reg1146 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1147 = (1'h0);
  reg [(3'h5):(1'h0)] reg1148 = (1'h0);
  reg [(4'he):(1'h0)] reg1149 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1151 = (1'h0);
  reg [(3'h4):(1'h0)] reg1152 = (1'h0);
  reg [(3'h6):(1'h0)] reg1153 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1154 = (1'h0);
  reg [(4'h9):(1'h0)] reg1158 = (1'h0);
  reg [(2'h2):(1'h0)] reg1159 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1160 = (1'h0);
  reg [(4'ha):(1'h0)] reg1161 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1165 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1166 = (1'h0);
  reg [(5'h10):(1'h0)] reg1167 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1168 = (1'h0);
  reg [(4'he):(1'h0)] reg1170 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1894 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1892 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1890 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1888 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1883 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1882 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1881 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1880 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1824 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1870 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1864 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1852 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1855 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1850 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1847 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1843 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1839 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1835 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1827 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1833 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1828 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1823 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1817 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1813 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1812 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1810 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1802 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1800 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1797 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1790 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1786 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1778 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1770 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1765 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1757 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1768 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1762 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1759 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1756 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1755 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1169 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1164 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1163 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1162 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1157 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1156 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1155 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1150 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1145 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1141 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1139 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1138 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1137 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1133 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1129 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1126 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1121 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1112 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1110 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1089 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1122 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1120 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1115 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1108 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1107 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1103 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1102 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1090 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1099 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1094 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1091 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar721 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar735 = (1'h0);
  reg [(4'h9):(1'h0)] forvar733 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar726 = (1'h0);
  reg [(4'h9):(1'h0)] forvar716 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar692 = (1'h0);
  reg [(4'ha):(1'h0)] forvar708 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar704 = (1'h0);
  reg [(4'he):(1'h0)] forvar695 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar693 = (1'h0);
  reg [(4'h9):(1'h0)] forvar725 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar723 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar722 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar719 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar687 = (1'h0);
  reg [(4'h8):(1'h0)] forvar710 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar709 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar703 = (1'h0);
  reg [(4'hb):(1'h0)] forvar701 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar700 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar696 = (1'h0);
  reg [(4'hb):(1'h0)] forvar690 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar686 = (1'h0);
  reg [(4'he):(1'h0)] forvar682 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar673 = (1'h0);
  reg [(2'h3):(1'h0)] forvar672 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar661 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar653 = (1'h0);
  reg [(4'hb):(1'h0)] forvar638 = (1'h0);
  reg [(4'h8):(1'h0)] forvar657 = (1'h0);
  reg [(3'h4):(1'h0)] forvar652 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar648 = (1'h0);
  reg [(3'h6):(1'h0)] forvar644 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar636 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar663 = (1'h0);
  reg [(4'he):(1'h0)] forvar659 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar651 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar650 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar647 = (1'h0);
  reg [(4'h8):(1'h0)] forvar643 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar642 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar637 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar634 = (1'h0);
  reg [(2'h2):(1'h0)] forvar633 = (1'h0);
  assign y = {wire1906,
                 wire1905,
                 wire1904,
                 wire1903,
                 wire1902,
                 wire1822,
                 wire1821,
                 wire1753,
                 wire1088,
                 wire1086,
                 wire632,
                 wire631,
                 wire629,
                 reg1901,
                 reg1900,
                 reg1899,
                 reg1898,
                 reg1897,
                 reg1896,
                 reg1895,
                 reg1893,
                 reg1891,
                 reg1889,
                 reg1887,
                 reg1886,
                 reg1885,
                 reg1884,
                 reg1823,
                 reg1879,
                 reg1878,
                 reg1877,
                 reg1876,
                 reg1875,
                 reg1874,
                 reg1873,
                 reg1872,
                 reg1871,
                 reg1869,
                 reg1868,
                 reg1867,
                 reg1866,
                 reg1865,
                 reg1863,
                 reg1862,
                 reg1861,
                 reg1860,
                 reg1859,
                 reg1858,
                 reg1857,
                 reg1855,
                 reg1856,
                 reg1854,
                 reg1853,
                 reg1852,
                 reg1851,
                 reg1849,
                 reg1848,
                 reg1846,
                 reg1845,
                 reg1844,
                 reg1842,
                 reg1841,
                 reg1840,
                 reg1828,
                 reg1838,
                 reg1837,
                 reg1836,
                 reg1835,
                 reg1834,
                 reg1832,
                 reg1831,
                 reg1830,
                 reg1829,
                 reg1827,
                 reg1826,
                 reg1825,
                 reg1824,
                 reg1820,
                 reg1819,
                 reg1818,
                 reg1816,
                 reg1815,
                 reg1814,
                 reg1811,
                 reg1809,
                 reg1808,
                 reg1807,
                 reg1806,
                 reg1805,
                 reg1804,
                 reg1803,
                 reg1801,
                 reg1799,
                 reg1798,
                 reg1796,
                 reg1795,
                 reg1794,
                 reg1793,
                 reg1792,
                 reg1791,
                 reg1789,
                 reg1788,
                 reg1787,
                 reg1785,
                 reg1784,
                 reg1783,
                 reg1782,
                 reg1781,
                 reg1780,
                 reg1779,
                 reg1778,
                 reg1777,
                 reg1776,
                 reg1768,
                 reg1759,
                 reg1775,
                 reg1774,
                 reg1773,
                 reg1772,
                 reg1771,
                 reg1762,
                 reg1770,
                 reg1769,
                 reg1767,
                 reg1766,
                 reg1765,
                 reg1764,
                 reg1763,
                 reg1761,
                 reg1760,
                 reg1758,
                 reg1757,
                 reg635,
                 reg636,
                 reg638,
                 reg639,
                 reg640,
                 reg641,
                 reg644,
                 reg645,
                 reg646,
                 reg648,
                 reg649,
                 reg652,
                 reg653,
                 reg654,
                 reg655,
                 reg656,
                 reg657,
                 reg658,
                 reg660,
                 reg661,
                 reg662,
                 reg664,
                 reg665,
                 reg666,
                 reg634,
                 reg637,
                 reg643,
                 reg647,
                 reg650,
                 reg651,
                 reg659,
                 reg642,
                 reg663,
                 reg667,
                 reg668,
                 reg669,
                 reg670,
                 reg671,
                 reg674,
                 reg675,
                 reg676,
                 reg677,
                 reg678,
                 reg679,
                 reg680,
                 reg681,
                 reg683,
                 reg684,
                 reg685,
                 reg687,
                 reg688,
                 reg689,
                 reg691,
                 reg692,
                 reg693,
                 reg694,
                 reg695,
                 reg697,
                 reg698,
                 reg699,
                 reg702,
                 reg704,
                 reg705,
                 reg706,
                 reg707,
                 reg708,
                 reg711,
                 reg712,
                 reg713,
                 reg714,
                 reg715,
                 reg716,
                 reg717,
                 reg718,
                 reg690,
                 reg720,
                 reg721,
                 reg724,
                 reg726,
                 reg727,
                 reg728,
                 reg729,
                 reg701,
                 reg703,
                 reg709,
                 reg696,
                 reg719,
                 reg722,
                 reg723,
                 reg725,
                 reg730,
                 reg731,
                 reg732,
                 reg733,
                 reg734,
                 reg736,
                 reg737,
                 reg738,
                 reg1089,
                 reg1090,
                 reg1092,
                 reg1093,
                 reg1095,
                 reg1096,
                 reg1097,
                 reg1098,
                 reg1100,
                 reg1091,
                 reg1094,
                 reg1099,
                 reg1101,
                 reg1102,
                 reg1103,
                 reg1104,
                 reg1105,
                 reg1106,
                 reg1107,
                 reg1108,
                 reg1109,
                 reg1110,
                 reg1111,
                 reg1112,
                 reg1113,
                 reg1114,
                 reg1116,
                 reg1117,
                 reg1118,
                 reg1119,
                 reg1121,
                 reg1122,
                 reg1123,
                 reg1124,
                 reg1125,
                 reg1126,
                 reg1120,
                 reg1127,
                 reg1115,
                 reg1128,
                 reg1130,
                 reg1131,
                 reg1132,
                 reg1134,
                 reg1135,
                 reg1136,
                 reg1140,
                 reg1142,
                 reg1143,
                 reg1144,
                 reg1146,
                 reg1147,
                 reg1148,
                 reg1149,
                 reg1151,
                 reg1152,
                 reg1153,
                 reg1154,
                 reg1158,
                 reg1159,
                 reg1160,
                 reg1161,
                 reg1165,
                 reg1166,
                 reg1167,
                 reg1168,
                 reg1170,
                 forvar1894,
                 forvar1892,
                 forvar1890,
                 forvar1888,
                 forvar1883,
                 forvar1882,
                 forvar1881,
                 forvar1880,
                 forvar1824,
                 forvar1870,
                 forvar1864,
                 forvar1852,
                 forvar1855,
                 forvar1850,
                 forvar1847,
                 forvar1843,
                 forvar1839,
                 forvar1835,
                 forvar1827,
                 forvar1833,
                 forvar1828,
                 forvar1823,
                 forvar1817,
                 forvar1813,
                 forvar1812,
                 forvar1810,
                 forvar1802,
                 forvar1800,
                 forvar1797,
                 forvar1790,
                 forvar1786,
                 forvar1778,
                 forvar1770,
                 forvar1765,
                 forvar1757,
                 forvar1768,
                 forvar1762,
                 forvar1759,
                 forvar1756,
                 forvar1755,
                 forvar1169,
                 forvar1164,
                 forvar1163,
                 forvar1162,
                 forvar1157,
                 forvar1156,
                 forvar1155,
                 forvar1150,
                 forvar1145,
                 forvar1141,
                 forvar1139,
                 forvar1138,
                 forvar1137,
                 forvar1133,
                 forvar1129,
                 forvar1126,
                 forvar1121,
                 forvar1112,
                 forvar1110,
                 forvar1089,
                 forvar1122,
                 forvar1120,
                 forvar1115,
                 forvar1108,
                 forvar1107,
                 forvar1103,
                 forvar1102,
                 forvar1090,
                 forvar1099,
                 forvar1094,
                 forvar1091,
                 forvar721,
                 forvar735,
                 forvar733,
                 forvar726,
                 forvar716,
                 forvar692,
                 forvar708,
                 forvar704,
                 forvar695,
                 forvar693,
                 forvar725,
                 forvar723,
                 forvar722,
                 forvar719,
                 forvar687,
                 forvar710,
                 forvar709,
                 forvar703,
                 forvar701,
                 forvar700,
                 forvar696,
                 forvar690,
                 forvar686,
                 forvar682,
                 forvar673,
                 forvar672,
                 forvar661,
                 forvar653,
                 forvar638,
                 forvar657,
                 forvar652,
                 forvar648,
                 forvar644,
                 forvar636,
                 forvar663,
                 forvar659,
                 forvar651,
                 forvar650,
                 forvar647,
                 forvar643,
                 forvar642,
                 forvar637,
                 forvar634,
                 forvar633,
                 (1'h0)};
  module5 #() modinst630 (.clk(clk), .wire8(wire0), .wire7(wire2), .wire6(wire1), .wire10(wire3), .wire9(wire4), .y(wire629));
  assign wire631 = $unsigned($unsigned((^~{wire3})));
  assign wire632 = $signed($signed(wire4[(2'h2):(1'h0)]));
  always
    @(posedge clk) begin
      if ($unsigned($signed($unsigned(wire2))))
        begin
          for (forvar633 = (1'h0); (forvar633 < (1'h0)); forvar633 = (forvar633 + (1'h1)))
            begin
              for (forvar634 = (1'h0); (forvar634 < (2'h3)); forvar634 = (forvar634 + (1'h1)))
                begin
                  reg635 <= (~({$unsigned(forvar633)} ?
                      (wire2 ? wire2 : $signed(wire4)) : (|$signed(wire629))));
                  reg636 <= $signed($unsigned((forvar634[(2'h3):(2'h2)] ?
                      forvar634[(3'h7):(3'h7)] : wire631[(1'h1):(1'h1)])));
                  for (forvar637 = (1'h0); (forvar637 < (2'h2)); forvar637 = (forvar637 + (1'h1)))
                    begin
                      reg638 <= {$unsigned(wire0)};
                      reg639 <= ($signed(($unsigned((8'ha5)) >= reg638)) <<< wire0);
                      reg640 <= wire2;
                      reg641 <= ((8'ha1) <= $unsigned(wire1));
                    end
                end
              for (forvar642 = (1'h0); (forvar642 < (1'h1)); forvar642 = (forvar642 + (1'h1)))
                begin
                  for (forvar643 = (1'h0); (forvar643 < (1'h0)); forvar643 = (forvar643 + (1'h1)))
                    begin
                      reg644 <= forvar634[(3'h7):(3'h5)];
                      reg645 <= $signed((($unsigned(wire3) >> wire4[(2'h3):(2'h2)]) ?
                          ((-forvar642) <<< (reg635 ?
                              (8'hb4) : forvar634)) : ($unsigned(reg641) ?
                              forvar634[(2'h2):(2'h2)] : ((8'hb7) ?
                                  (8'hba) : forvar637))));
                      reg646 <= ((~|$signed((reg635 & forvar637))) ?
                          ((8'hb3) ?
                              (((8'h9d) ?
                                  reg635 : wire4) < wire631) : (-reg635[(3'h4):(3'h4)])) : $signed((wire4 || $unsigned((8'ha9)))));
                    end
                  for (forvar647 = (1'h0); (forvar647 < (2'h2)); forvar647 = (forvar647 + (1'h1)))
                    begin
                      reg648 <= (+(^~reg635[(3'h5):(3'h4)]));
                      reg649 <= forvar637;
                    end
                end
            end
          for (forvar650 = (1'h0); (forvar650 < (2'h3)); forvar650 = (forvar650 + (1'h1)))
            begin
              for (forvar651 = (1'h0); (forvar651 < (2'h3)); forvar651 = (forvar651 + (1'h1)))
                begin
                  if (reg648[(3'h6):(1'h1)])
                    begin
                      reg652 <= ((wire631 ~^ ($unsigned(reg639) ?
                          forvar650 : forvar633[(1'h1):(1'h1)])) ^ reg638);
                      reg653 <= $unsigned(forvar647);
                      reg654 <= {$unsigned((forvar633[(1'h0):(1'h0)] ?
                              (reg653 ? (8'ha3) : reg636) : (forvar643 ?
                                  forvar642 : reg639)))};
                    end
                  else
                    begin
                      reg652 <= forvar647;
                      reg653 <= $unsigned(((!{reg652}) | (|$signed(wire632))));
                    end
                  if ((8'hb9))
                    begin
                      reg655 <= $signed(((~$unsigned(reg638)) + wire632));
                    end
                  else
                    begin
                      reg655 <= forvar650[(1'h1):(1'h1)];
                      reg656 <= $unsigned($signed(wire1[(3'h4):(1'h1)]));
                      reg657 <= (^~reg656[(4'h9):(1'h0)]);
                      reg658 <= forvar634;
                    end
                  for (forvar659 = (1'h0); (forvar659 < (2'h3)); forvar659 = (forvar659 + (1'h1)))
                    begin
                      reg660 <= wire3;
                      reg661 <= (~(^~($signed((8'had)) * (wire632 ?
                          reg652 : wire1))));
                      reg662 <= (~^(^~$signed(((8'ha1) >= (8'ha3)))));
                    end
                end
              for (forvar663 = (1'h0); (forvar663 < (2'h2)); forvar663 = (forvar663 + (1'h1)))
                begin
                  if (wire629)
                    begin
                      reg664 <= {({$unsigned(reg644)} ?
                              ((reg653 ? reg652 : forvar647) ?
                                  (reg639 ?
                                      reg636 : reg638) : (!reg656)) : reg638)};
                      reg665 <= $signed($unsigned($signed(((8'ha0) >= wire1))));
                      reg666 <= (reg662 == $unsigned(reg661));
                    end
                  else
                    begin
                      reg664 <= wire3[(3'h4):(3'h4)];
                    end
                end
            end
        end
      else
        begin
          if (({$signed({reg658})} <= (((8'hb3) >>> forvar643[(4'h8):(2'h2)]) * {(reg648 ?
                  forvar633 : forvar650)})))
            begin
              for (forvar633 = (1'h0); (forvar633 < (1'h1)); forvar633 = (forvar633 + (1'h1)))
                begin
                  if ($unsigned(reg649))
                    begin
                      reg634 <= $signed((reg661 || ((forvar634 ?
                          reg639 : reg649) <<< ((8'ha0) ^ reg645))));
                    end
                  else
                    begin
                      reg634 <= ((($signed((8'ha8)) ?
                                  (forvar633 <<< forvar643) : (reg646 ?
                                      (8'ha8) : wire2)) ?
                              forvar634 : reg652) ?
                          (((reg635 == reg654) ~^ $signed(forvar651)) ?
                              ($unsigned(reg662) ?
                                  (|reg662) : (~reg662)) : wire1) : (~&($unsigned(forvar637) ~^ reg657)));
                      reg635 <= $signed((reg638[(2'h3):(2'h2)] != $signed((reg664 || (8'hb2)))));
                    end
                  for (forvar636 = (1'h0); (forvar636 < (2'h2)); forvar636 = (forvar636 + (1'h1)))
                    begin
                      reg637 <= ((reg653[(3'h5):(2'h3)] ?
                              ((reg635 >>> reg639) ?
                                  reg645[(1'h0):(1'h0)] : (reg636 ?
                                      forvar633 : wire2)) : (~^{reg665})) ?
                          ((~|(forvar659 >>> forvar633)) ?
                              forvar650[(2'h2):(2'h2)] : reg653) : (^~forvar642[(3'h5):(2'h2)]));
                      reg638 <= (forvar634 >= {reg640[(1'h1):(1'h0)]});
                      reg639 <= forvar636;
                    end
                  reg640 <= $unsigned(((reg636 ? $signed(forvar663) : wire0) ?
                      $signed($signed((8'ha8))) : (reg662 != (wire631 > reg637))));
                  reg641 <= $unsigned(((|$unsigned((8'hb6))) ?
                      ((^~reg664) ?
                          (8'ha3) : ((8'h9c) ?
                              wire632 : reg639)) : wire629[(3'h7):(3'h4)]));
                end
              for (forvar642 = (1'h0); (forvar642 < (1'h0)); forvar642 = (forvar642 + (1'h1)))
                begin
                  if ($unsigned(reg636[(3'h6):(2'h3)]))
                    begin
                      reg643 <= (forvar636 * (^($signed(reg644) ?
                          reg658[(4'h8):(4'h8)] : reg655)));
                    end
                  else
                    begin
                      reg643 <= wire4[(3'h6):(1'h1)];
                    end
                  for (forvar644 = (1'h0); (forvar644 < (2'h2)); forvar644 = (forvar644 + (1'h1)))
                    begin
                      reg645 <= $signed(forvar644[(2'h2):(1'h1)]);
                    end
                  if (reg662)
                    begin
                      reg646 <= $unsigned(($signed(forvar637[(3'h6):(1'h0)]) ?
                          $unsigned($unsigned(reg637)) : reg649[(4'hb):(3'h7)]));
                    end
                  else
                    begin
                      reg646 <= ((~^forvar644) << wire0[(4'hb):(3'h5)]);
                      reg647 <= ((-(~&forvar663)) ?
                          (8'ha7) : $signed(($unsigned(forvar636) ?
                              {forvar643} : reg644[(2'h3):(2'h3)])));
                    end
                  for (forvar648 = (1'h0); (forvar648 < (1'h0)); forvar648 = (forvar648 + (1'h1)))
                    begin
                      reg649 <= reg636;
                      reg650 <= reg648[(3'h6):(2'h2)];
                      reg651 <= $unsigned($signed(reg648));
                    end
                end
              if (((reg658 ?
                  wire631 : $unsigned((!reg651))) >= (reg665 ^~ $signed((~forvar663)))))
                begin
                  for (forvar652 = (1'h0); (forvar652 < (2'h2)); forvar652 = (forvar652 + (1'h1)))
                    begin
                      reg653 <= ($unsigned(((^~reg644) || (^~wire1))) ?
                          $unsigned(($signed(reg643) != (^~wire631))) : (({reg657} - {(8'had)}) ?
                              $unsigned(wire629[(2'h3):(1'h0)]) : ($signed(reg638) ~^ wire0[(4'hb):(4'h9)])));
                      reg654 <= reg644;
                      reg655 <= wire2[(4'h9):(2'h2)];
                      reg656 <= {{$signed((forvar650 & reg658))}};
                    end
                end
              else
                begin
                  if ($signed((((reg649 || forvar644) ^~ reg656[(3'h4):(1'h1)]) >= (~|(reg658 ?
                      reg664 : forvar643)))))
                    begin
                      reg652 <= forvar648;
                      reg653 <= $unsigned(reg662);
                      reg654 <= (-reg647);
                      reg655 <= wire0[(4'h8):(3'h6)];
                    end
                  else
                    begin
                      reg652 <= (~^wire631);
                      reg653 <= (^~wire631);
                    end
                  reg656 <= (($unsigned($unsigned((8'ha6))) ?
                      $unsigned($unsigned(reg650)) : {(forvar651 ^ reg639)}) + $unsigned(reg650));
                end
              if (forvar647[(1'h0):(1'h0)])
                begin
                  if ((($signed(reg653[(1'h0):(1'h0)]) ?
                      {(wire632 << (8'hab))} : reg657[(4'h9):(2'h2)]) < {forvar659}))
                    begin
                      reg657 <= $unsigned((reg660 >= $unsigned($unsigned(reg639))));
                      reg658 <= ($signed((wire631[(3'h6):(1'h1)] == $unsigned(reg637))) ?
                          $signed($unsigned(reg647[(4'h8):(2'h3)])) : ($unsigned(reg641) >> (^reg644)));
                      reg659 <= reg666;
                      reg660 <= $signed($unsigned(reg648[(4'h9):(4'h9)]));
                    end
                  else
                    begin
                      reg657 <= {({$unsigned(reg666)} & $unsigned(wire0[(4'h9):(4'h9)]))};
                      reg658 <= $signed(reg655[(4'h8):(3'h5)]);
                    end
                end
              else
                begin
                  for (forvar657 = (1'h0); (forvar657 < (2'h3)); forvar657 = (forvar657 + (1'h1)))
                    begin
                      reg658 <= (~|reg665[(1'h0):(1'h0)]);
                    end
                  for (forvar659 = (1'h0); (forvar659 < (1'h1)); forvar659 = (forvar659 + (1'h1)))
                    begin
                      reg660 <= reg662[(1'h0):(1'h0)];
                      reg661 <= (~reg639);
                    end
                end
            end
          else
            begin
              for (forvar633 = (1'h0); (forvar633 < (1'h0)); forvar633 = (forvar633 + (1'h1)))
                begin
                  if ($signed($signed($unsigned(wire4))))
                    begin
                      reg634 <= {(~&{(~&reg639)})};
                      reg635 <= forvar642[(3'h5):(3'h4)];
                      reg636 <= reg651[(1'h1):(1'h1)];
                      reg637 <= reg664[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg634 <= ($signed($signed((&(8'haa)))) ?
                          $signed($unsigned((reg659 ?
                              reg651 : reg665))) : (8'ha8));
                      reg635 <= $unsigned((8'ha0));
                    end
                end
              for (forvar638 = (1'h0); (forvar638 < (2'h3)); forvar638 = (forvar638 + (1'h1)))
                begin
                  if ((|((~&(-wire632)) && ((forvar650 >= forvar642) == (~|forvar650)))))
                    begin
                      reg639 <= ((!(^$unsigned(forvar637))) ?
                          reg657[(1'h0):(1'h0)] : forvar648[(4'hb):(4'h8)]);
                      reg640 <= (reg651 >>> ((forvar644 ?
                              $signed(reg658) : reg647[(3'h6):(1'h1)]) ?
                          $unsigned((!reg666)) : (8'ha9)));
                      reg641 <= $signed(($signed((forvar642 ?
                              (8'h9d) : forvar657)) ?
                          reg643 : reg660));
                      reg642 <= $unsigned(({reg661[(3'h4):(3'h4)]} ?
                          ((&wire629) ?
                              (reg635 ?
                                  reg664 : forvar633) : (~forvar643)) : $signed(reg652)));
                    end
                  else
                    begin
                      reg639 <= $signed((~^$unsigned(((8'hba) ?
                          forvar633 : (8'hba)))));
                      reg640 <= $signed($signed(($unsigned(forvar637) ?
                          {forvar633} : $signed(reg649))));
                    end
                  for (forvar643 = (1'h0); (forvar643 < (2'h3)); forvar643 = (forvar643 + (1'h1)))
                    begin
                      reg644 <= (8'hb8);
                      reg645 <= (-($signed((wire1 && (8'had))) | {(forvar633 ?
                              forvar657 : reg662)}));
                      reg646 <= (~|$signed($signed(reg653[(1'h1):(1'h1)])));
                    end
                  reg647 <= forvar651[(1'h0):(1'h0)];
                end
              for (forvar648 = (1'h0); (forvar648 < (1'h1)); forvar648 = (forvar648 + (1'h1)))
                begin
                  if ((^$signed((wire632 ?
                      $unsigned(reg661) : reg641[(2'h2):(1'h1)]))))
                    begin
                      reg649 <= reg646;
                      reg650 <= (&$unsigned((!wire0[(2'h3):(2'h2)])));
                    end
                  else
                    begin
                      reg649 <= $unsigned($unsigned((^$unsigned(forvar643))));
                      reg650 <= $unsigned(forvar652[(2'h2):(1'h0)]);
                    end
                  if (forvar634)
                    begin
                      reg651 <= reg640;
                      reg652 <= ($unsigned($signed($unsigned(forvar637))) << (~^(~|((8'ha1) <= forvar663))));
                    end
                  else
                    begin
                      reg651 <= wire0;
                    end
                  for (forvar653 = (1'h0); (forvar653 < (1'h0)); forvar653 = (forvar653 + (1'h1)))
                    begin
                      reg654 <= (^~forvar650[(2'h2):(2'h2)]);
                      reg655 <= wire629;
                      reg656 <= (reg642 ?
                          (&{$unsigned(wire1)}) : reg635[(3'h7):(2'h2)]);
                    end
                end
              if ($signed($unsigned($signed((reg636 && reg646)))))
                begin
                  reg657 <= ((~^{(forvar648 <<< reg636)}) >= reg651);
                  if (wire632)
                    begin
                      reg658 <= $signed({$unsigned($unsigned(reg664))});
                      reg659 <= {$unsigned($unsigned({reg658}))};
                      reg660 <= forvar659[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg658 <= $signed(forvar659[(1'h1):(1'h0)]);
                      reg659 <= {reg653[(2'h3):(2'h3)]};
                      reg660 <= {$unsigned((~^(reg658 >> reg636)))};
                      reg661 <= {$unsigned(((~forvar633) ?
                              $unsigned(forvar643) : (^forvar638)))};
                    end
                end
              else
                begin
                  if (reg642[(3'h7):(1'h1)])
                    begin
                      reg657 <= {wire2};
                      reg658 <= ({$signed((8'hb0))} ?
                          {({wire2} <<< $unsigned(reg642))} : $signed({(^reg647)}));
                      reg659 <= $unsigned(forvar634);
                      reg660 <= reg665[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg657 <= {wire4};
                      reg658 <= forvar652[(2'h3):(1'h1)];
                      reg659 <= reg658;
                    end
                  for (forvar661 = (1'h0); (forvar661 < (2'h2)); forvar661 = (forvar661 + (1'h1)))
                    begin
                      reg662 <= (reg638[(3'h5):(1'h1)] >= $unsigned(forvar650));
                      reg663 <= $signed(reg659[(3'h5):(2'h2)]);
                    end
                  if ($signed(({reg661[(1'h1):(1'h0)]} ? {(~reg661)} : reg658)))
                    begin
                      reg664 <= (($unsigned(reg650) ?
                          ((reg647 - reg664) ?
                              (reg647 || reg636) : (reg664 >> wire1)) : ((|forvar642) && (!wire2))) <<< (reg646[(1'h0):(1'h0)] ?
                          ((~|reg656) ?
                              $unsigned(wire2) : reg656[(2'h3):(2'h2)]) : {{forvar652}}));
                      reg665 <= $unsigned(reg659[(3'h5):(2'h2)]);
                      reg666 <= reg637;
                      reg667 <= wire1;
                    end
                  else
                    begin
                      reg664 <= {(($unsigned(reg659) ?
                              {forvar663} : (forvar633 ?
                                  forvar634 : (8'hac))) | (~{(8'hac)}))};
                      reg665 <= $signed(forvar647);
                      reg666 <= {forvar647[(4'h8):(3'h4)]};
                      reg667 <= $signed($signed({(forvar643 << reg650)}));
                    end
                  if ((~|(&reg637[(1'h0):(1'h0)])))
                    begin
                      reg668 <= (~&(+$unsigned($unsigned(reg664))));
                      reg669 <= forvar659;
                      reg670 <= $signed((forvar657 + (~&reg645)));
                      reg671 <= $unsigned(reg635[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg668 <= $unsigned($unsigned(((~^forvar659) - (wire631 ~^ forvar659))));
                      reg669 <= ((reg637 >> $signed((~|forvar663))) ?
                          $signed(wire4) : (forvar634 & ($signed(wire0) ?
                              (reg649 && reg657) : {reg656})));
                    end
                end
            end
          for (forvar672 = (1'h0); (forvar672 < (1'h1)); forvar672 = (forvar672 + (1'h1)))
            begin
              for (forvar673 = (1'h0); (forvar673 < (1'h0)); forvar673 = (forvar673 + (1'h1)))
                begin
                  reg674 <= reg666[(4'h9):(3'h5)];
                end
              if (forvar636[(3'h6):(3'h4)])
                begin
                  if (reg651[(3'h6):(3'h5)])
                    begin
                      reg675 <= (~{$signed(((8'hb6) <<< wire631))});
                      reg676 <= $signed($signed(($unsigned(reg657) ?
                          $signed(wire4) : $unsigned(reg666))));
                      reg677 <= ((8'h9c) ?
                          ($signed($unsigned(wire631)) <<< $signed((reg635 ?
                              reg641 : forvar637))) : reg649);
                    end
                  else
                    begin
                      reg675 <= (reg664 ?
                          $unsigned($unsigned(forvar652)) : (($unsigned((8'h9f)) ^ reg641[(4'hf):(3'h5)]) * ($unsigned(reg667) >> reg675[(4'ha):(2'h2)])));
                      reg676 <= wire632[(1'h0):(1'h0)];
                      reg677 <= $signed(forvar650[(1'h1):(1'h0)]);
                      reg678 <= $signed($signed($signed(((8'hb2) ?
                          reg674 : (8'hb6)))));
                    end
                  reg679 <= ($signed((-(reg634 ?
                      reg654 : forvar647))) + ((8'hba) ?
                      $signed({reg640}) : reg645));
                end
              else
                begin
                  if (reg655[(3'h7):(3'h7)])
                    begin
                      reg675 <= {(((wire629 ? reg678 : reg658) ?
                                  reg655 : reg662[(2'h3):(1'h1)]) ?
                              forvar642[(4'h9):(1'h0)] : $unsigned($unsigned(forvar653)))};
                      reg676 <= ({reg662[(3'h4):(3'h4)]} * reg666[(3'h4):(2'h3)]);
                      reg677 <= forvar634[(3'h6):(3'h4)];
                      reg678 <= wire1[(4'ha):(4'ha)];
                    end
                  else
                    begin
                      reg675 <= $signed({reg674[(4'hb):(4'hb)]});
                      reg676 <= {reg674[(4'hd):(3'h7)]};
                    end
                  if ({$unsigned($unsigned((wire629 ? (8'ha0) : (8'hb5))))})
                    begin
                      reg679 <= reg665;
                      reg680 <= $signed($signed(reg637));
                    end
                  else
                    begin
                      reg679 <= (!(wire3[(1'h0):(1'h0)] ~^ $signed(forvar653[(2'h3):(1'h1)])));
                      reg680 <= forvar661[(4'h8):(3'h5)];
                    end
                  if (reg664[(3'h7):(3'h5)])
                    begin
                      reg681 <= reg651[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg681 <= (($signed(reg666[(1'h0):(1'h0)]) | reg667) ?
                          forvar650 : $unsigned(($unsigned(reg676) ?
                              reg644 : ((8'haf) << reg667))));
                    end
                  for (forvar682 = (1'h0); (forvar682 < (1'h0)); forvar682 = (forvar682 + (1'h1)))
                    begin
                      reg683 <= $unsigned(forvar633[(1'h1):(1'h0)]);
                    end
                end
              reg684 <= (8'ha8);
            end
        end
      reg685 <= reg683;
      if ((($signed(reg647[(2'h3):(2'h2)]) ?
          $signed($unsigned(forvar650)) : $unsigned({reg642})) < $unsigned($unsigned(forvar653[(3'h5):(2'h2)]))))
        begin
          if (reg651)
            begin
              for (forvar686 = (1'h0); (forvar686 < (2'h2)); forvar686 = (forvar686 + (1'h1)))
                begin
                  if (((((reg640 | (8'hb6)) ? reg645 : $signed(forvar657)) ?
                          $signed((forvar644 * reg667)) : $unsigned((|reg676))) ?
                      forvar638[(2'h3):(2'h2)] : ($signed((wire632 <<< reg680)) | (reg657[(3'h7):(3'h6)] ?
                          reg640 : {reg685}))))
                    begin
                      reg687 <= ($unsigned((!reg667)) ? (8'ha8) : reg665);
                      reg688 <= (reg656[(2'h3):(1'h0)] >>> $signed((!reg663[(4'ha):(4'h8)])));
                      reg689 <= (($signed((forvar659 ?
                              reg657 : wire2)) + (|(reg653 ?
                              reg645 : reg635))) ?
                          $unsigned((~|reg634)) : $signed((^~forvar650)));
                    end
                  else
                    begin
                      reg687 <= wire632[(4'ha):(1'h0)];
                      reg688 <= (8'haa);
                    end
                  for (forvar690 = (1'h0); (forvar690 < (1'h1)); forvar690 = (forvar690 + (1'h1)))
                    begin
                      reg691 <= (8'hb1);
                    end
                  if ($unsigned(reg662))
                    begin
                      reg692 <= (8'hb2);
                      reg693 <= wire629;
                      reg694 <= $unsigned(($signed((reg648 ? reg645 : reg663)) ?
                          $unsigned((8'ha9)) : ((reg661 && (8'h9d)) ?
                              (+forvar634) : wire631[(3'h6):(1'h0)])));
                      reg695 <= forvar686;
                    end
                  else
                    begin
                      reg692 <= forvar690[(3'h5):(3'h5)];
                      reg693 <= (^~reg675[(4'h8):(3'h4)]);
                    end
                  for (forvar696 = (1'h0); (forvar696 < (2'h3)); forvar696 = (forvar696 + (1'h1)))
                    begin
                      reg697 <= forvar642[(4'hb):(4'h8)];
                      reg698 <= (((8'h9d) ?
                          (^(reg664 ?
                              forvar672 : forvar661)) : forvar690[(1'h1):(1'h0)]) ^ (~&reg652));
                      reg699 <= {(8'ha9)};
                    end
                end
              for (forvar700 = (1'h0); (forvar700 < (1'h1)); forvar700 = (forvar700 + (1'h1)))
                begin
                  for (forvar701 = (1'h0); (forvar701 < (1'h1)); forvar701 = (forvar701 + (1'h1)))
                    begin
                      reg702 <= $unsigned(forvar682[(4'h9):(3'h4)]);
                    end
                  for (forvar703 = (1'h0); (forvar703 < (1'h1)); forvar703 = (forvar703 + (1'h1)))
                    begin
                      reg704 <= reg638;
                      reg705 <= (+$unsigned(((forvar657 ? reg697 : forvar633) ?
                          reg678 : (forvar643 ^~ forvar650))));
                      reg706 <= reg692;
                      reg707 <= (reg698[(2'h2):(1'h1)] * $signed(((forvar633 ?
                          reg658 : forvar653) << $signed(reg642))));
                    end
                end
              reg708 <= (8'h9c);
              for (forvar709 = (1'h0); (forvar709 < (2'h2)); forvar709 = (forvar709 + (1'h1)))
                begin
                  for (forvar710 = (1'h0); (forvar710 < (1'h1)); forvar710 = (forvar710 + (1'h1)))
                    begin
                      reg711 <= ((($signed(reg638) ?
                                  (|reg642) : (reg680 >= reg667)) ?
                              forvar709 : {$unsigned((8'ha5))}) ?
                          $signed(wire629) : (+(+$signed(reg654))));
                      reg712 <= $unsigned($unsigned({(^reg639)}));
                      reg713 <= $signed({reg635[(1'h0):(1'h0)]});
                      reg714 <= forvar700[(4'hc):(4'ha)];
                    end
                  if ((!(reg669 >> $unsigned(reg698[(4'h9):(4'h8)]))))
                    begin
                      reg715 <= $unsigned($signed((wire3 == reg656[(2'h3):(2'h2)])));
                      reg716 <= ($signed(reg635) ?
                          {reg661[(2'h3):(2'h2)]} : (reg702 ?
                              (-forvar633[(1'h0):(1'h0)]) : ($signed(reg634) * (|(8'haa)))));
                      reg717 <= (forvar700[(3'h5):(1'h1)] & ({(reg661 ?
                                  (8'hb9) : forvar650)} ?
                          $unsigned((forvar672 & (8'ha7))) : wire2));
                      reg718 <= (8'hb8);
                    end
                  else
                    begin
                      reg715 <= ((((~^(8'hb2)) ?
                              $signed(reg712) : $unsigned(forvar701)) * wire632) ?
                          {($signed(reg638) ^~ {forvar634})} : ($unsigned($signed(reg666)) ?
                              ($signed(reg692) | $signed(forvar701)) : {$unsigned((8'hb3))}));
                      reg716 <= $signed(({(+reg706)} ^~ (!{reg692})));
                      reg717 <= (~|$signed((~&(8'hb8))));
                      reg718 <= ((~|reg671) ^ reg671);
                    end
                end
            end
          else
            begin
              for (forvar686 = (1'h0); (forvar686 < (1'h0)); forvar686 = (forvar686 + (1'h1)))
                begin
                  for (forvar687 = (1'h0); (forvar687 < (1'h1)); forvar687 = (forvar687 + (1'h1)))
                    begin
                      reg688 <= $unsigned(reg663[(3'h4):(2'h3)]);
                      reg689 <= $unsigned((8'hb7));
                      reg690 <= reg648;
                    end
                end
            end
          for (forvar719 = (1'h0); (forvar719 < (1'h1)); forvar719 = (forvar719 + (1'h1)))
            begin
              reg720 <= $signed(reg677[(2'h2):(1'h0)]);
              reg721 <= (-((((8'ha8) <= reg718) ? (~&reg643) : (&wire0)) ?
                  {(-reg679)} : $signed((reg681 > reg706))));
            end
          for (forvar722 = (1'h0); (forvar722 < (2'h2)); forvar722 = (forvar722 + (1'h1)))
            begin
              for (forvar723 = (1'h0); (forvar723 < (1'h1)); forvar723 = (forvar723 + (1'h1)))
                begin
                  reg724 <= reg644[(2'h2):(2'h2)];
                  for (forvar725 = (1'h0); (forvar725 < (2'h3)); forvar725 = (forvar725 + (1'h1)))
                    begin
                      reg726 <= (~^$signed(reg652[(1'h1):(1'h1)]));
                      reg727 <= ((~|((|reg684) >= {reg702})) ?
                          (8'hb3) : reg684);
                      reg728 <= ({reg691[(1'h1):(1'h1)]} * (!(((8'h9c) ?
                          reg666 : reg647) != $unsigned((8'ha0)))));
                    end
                end
            end
          reg729 <= (~&(8'hb7));
        end
      else
        begin
          if ((reg676 ?
              (reg694 ?
                  (~^(reg683 ? reg692 : forvar701)) : ((~reg718) ?
                      (8'hb9) : wire3[(1'h0):(1'h0)])) : ($signed((reg681 ?
                  reg721 : wire4)) > $unsigned($unsigned((8'hb3))))))
            begin
              for (forvar686 = (1'h0); (forvar686 < (2'h3)); forvar686 = (forvar686 + (1'h1)))
                begin
                  if ((|(8'hb1)))
                    begin
                      reg687 <= reg715;
                      reg688 <= (reg639 ~^ forvar725);
                    end
                  else
                    begin
                      reg687 <= ((+(~(reg684 <<< (8'hba)))) < {({forvar709} & reg690[(1'h0):(1'h0)])});
                      reg688 <= {$unsigned(((8'ha4) ?
                              $unsigned(reg642) : ((8'ha1) << reg712)))};
                      reg689 <= $unsigned((((forvar634 + reg713) ?
                              $unsigned(wire4) : reg708) ?
                          (~|reg720[(1'h1):(1'h0)]) : ((reg648 ?
                                  forvar644 : reg697) ?
                              ((8'hab) ? forvar696 : wire4) : {reg702})));
                      reg690 <= $signed(reg685[(3'h5):(1'h0)]);
                    end
                  if ($signed($unsigned(reg651)))
                    begin
                      reg691 <= (8'ha8);
                      reg692 <= (reg683[(2'h3):(1'h0)] || reg642);
                    end
                  else
                    begin
                      reg691 <= ({forvar636[(4'h9):(3'h7)]} && reg695);
                    end
                  for (forvar693 = (1'h0); (forvar693 < (2'h3)); forvar693 = (forvar693 + (1'h1)))
                    begin
                      reg694 <= $unsigned($signed($signed((reg646 != reg634))));
                    end
                end
              for (forvar695 = (1'h0); (forvar695 < (2'h3)); forvar695 = (forvar695 + (1'h1)))
                begin
                  for (forvar696 = (1'h0); (forvar696 < (2'h3)); forvar696 = (forvar696 + (1'h1)))
                    begin
                      reg697 <= $unsigned(reg713[(1'h1):(1'h1)]);
                      reg698 <= (!(((8'h9f) * $unsigned(reg716)) | {reg634}));
                      reg699 <= forvar719;
                    end
                  for (forvar700 = (1'h0); (forvar700 < (1'h1)); forvar700 = (forvar700 + (1'h1)))
                    begin
                      reg701 <= (((~|$signed(forvar644)) ?
                              {(^~reg637)} : (&(forvar725 ?
                                  forvar703 : forvar695))) ?
                          $signed((&reg640)) : $signed($signed(reg657[(1'h1):(1'h1)])));
                      reg702 <= $unsigned((^reg707));
                      reg703 <= $signed($signed($unsigned(reg676[(2'h3):(1'h0)])));
                    end
                end
              if ($signed(reg651))
                begin
                  for (forvar704 = (1'h0); (forvar704 < (2'h3)); forvar704 = (forvar704 + (1'h1)))
                    begin
                      reg705 <= reg724;
                      reg706 <= ($signed(($signed(wire0) + reg665)) + $unsigned((~|(reg703 ?
                          forvar642 : reg692))));
                      reg707 <= (^$unsigned(reg727[(4'h8):(3'h7)]));
                    end
                  for (forvar708 = (1'h0); (forvar708 < (2'h3)); forvar708 = (forvar708 + (1'h1)))
                    begin
                      reg709 <= (~reg676[(1'h0):(1'h0)]);
                    end
                  for (forvar710 = (1'h0); (forvar710 < (1'h0)); forvar710 = (forvar710 + (1'h1)))
                    begin
                      reg711 <= (reg684 >>> ({wire632[(4'hb):(3'h4)]} > ({forvar672} ?
                          $signed(forvar647) : {reg640})));
                      reg712 <= $unsigned((reg726[(4'h9):(1'h1)] ?
                          ($signed(reg642) ?
                              $signed(wire0) : reg671[(3'h4):(2'h3)]) : (^~(forvar704 + (8'h9d)))));
                      reg713 <= forvar634;
                      reg714 <= ($signed({$signed(forvar701)}) << {reg665[(2'h2):(1'h0)]});
                    end
                  reg715 <= forvar682;
                end
              else
                begin
                  reg704 <= forvar648;
                end
            end
          else
            begin
              for (forvar686 = (1'h0); (forvar686 < (2'h2)); forvar686 = (forvar686 + (1'h1)))
                begin
                  for (forvar687 = (1'h0); (forvar687 < (1'h0)); forvar687 = (forvar687 + (1'h1)))
                    begin
                      reg688 <= $signed(reg641);
                      reg689 <= reg667[(4'hc):(3'h5)];
                    end
                  for (forvar690 = (1'h0); (forvar690 < (1'h0)); forvar690 = (forvar690 + (1'h1)))
                    begin
                      reg691 <= forvar638[(3'h5):(3'h4)];
                    end
                  for (forvar692 = (1'h0); (forvar692 < (2'h3)); forvar692 = (forvar692 + (1'h1)))
                    begin
                      reg693 <= reg654;
                      reg694 <= forvar703[(4'ha):(4'h9)];
                      reg695 <= (8'hb1);
                      reg696 <= (+forvar709);
                    end
                  if (forvar672[(2'h3):(2'h3)])
                    begin
                      reg697 <= reg640;
                      reg698 <= {((~&$signed(wire1)) ?
                              $unsigned(reg666[(1'h1):(1'h0)]) : reg689)};
                    end
                  else
                    begin
                      reg697 <= ((8'hb8) * {reg669});
                      reg698 <= ((8'hb7) ?
                          forvar722 : $unsigned(reg713[(1'h1):(1'h1)]));
                      reg699 <= $unsigned(($unsigned($signed(reg634)) * reg702));
                    end
                end
            end
          if (forvar723[(3'h7):(3'h4)])
            begin
              if (reg659)
                begin
                  for (forvar716 = (1'h0); (forvar716 < (1'h0)); forvar716 = (forvar716 + (1'h1)))
                    begin
                      reg717 <= {(^~$unsigned((reg639 ? reg693 : reg685)))};
                      reg718 <= reg683;
                      reg719 <= $signed(reg675[(3'h4):(1'h1)]);
                      reg720 <= $unsigned({(((8'h9f) || reg684) ?
                              reg698 : (&(8'hb9)))});
                    end
                  if ($unsigned(reg668[(2'h2):(1'h1)]))
                    begin
                      reg721 <= $unsigned(reg646[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg721 <= reg684[(3'h6):(1'h0)];
                      reg722 <= reg702;
                      reg723 <= $unsigned(reg636[(3'h4):(3'h4)]);
                      reg724 <= wire632[(4'he):(4'hc)];
                    end
                  reg725 <= $signed(forvar695);
                  for (forvar726 = (1'h0); (forvar726 < (1'h1)); forvar726 = (forvar726 + (1'h1)))
                    begin
                      reg727 <= reg717[(3'h7):(3'h6)];
                      reg728 <= ((!((!reg678) >= $unsigned(reg707))) ?
                          ($signed(reg679[(4'ha):(1'h0)]) ?
                              forvar636 : ((-forvar633) ?
                                  $unsigned(reg680) : reg645[(1'h1):(1'h0)])) : (^~((~reg648) ?
                              (reg691 ? reg716 : forvar709) : ((8'hba) ?
                                  forvar644 : (8'ha9)))));
                      reg729 <= reg647;
                      reg730 <= (&(8'ha4));
                    end
                end
              else
                begin
                  if (reg659)
                    begin
                      reg716 <= $unsigned(forvar651[(2'h2):(2'h2)]);
                      reg717 <= (^~(($signed(reg662) ?
                          forvar722[(1'h1):(1'h0)] : (reg713 ?
                              reg655 : reg664)) != $signed((~&reg688))));
                      reg718 <= (forvar636[(3'h6):(3'h6)] ^ (~&(reg702[(4'hc):(4'hc)] ?
                          reg730[(2'h3):(1'h0)] : {forvar657})));
                      reg719 <= reg725[(3'h6):(2'h3)];
                    end
                  else
                    begin
                      reg716 <= forvar647[(3'h6):(2'h2)];
                      reg717 <= ($unsigned(((reg721 ? forvar648 : reg718) ?
                          reg727[(4'h8):(4'h8)] : (~|forvar638))) + {(~^(&reg727))});
                      reg718 <= (~((|reg648[(1'h1):(1'h1)]) ?
                          reg698 : ($signed(wire2) ?
                              (reg687 && reg699) : $unsigned(reg643))));
                      reg719 <= (~&(~|$unsigned((reg690 ?
                          forvar719 : reg689))));
                    end
                end
              if (reg647)
                begin
                  if ((~^$signed($signed(reg636[(3'h7):(2'h2)]))))
                    begin
                      reg731 <= (&reg638);
                    end
                  else
                    begin
                      reg731 <= (reg696[(3'h4):(3'h4)] ?
                          (reg707[(1'h0):(1'h0)] ?
                              $signed((reg719 ?
                                  forvar701 : reg697)) : $unsigned(((8'hb9) ^ (8'hba)))) : $signed({reg688}));
                      reg732 <= ($signed(reg716[(5'h10):(4'hd)]) + $signed(((reg654 * forvar682) >> (forvar709 != reg693))));
                      reg733 <= ((((reg690 * forvar703) && (!forvar710)) ?
                              (-reg650) : reg715[(1'h0):(1'h0)]) ?
                          $signed(reg688[(1'h1):(1'h0)]) : ($unsigned(forvar686[(4'hb):(4'ha)]) && {(reg723 && reg647)}));
                    end
                end
              else
                begin
                  if ((8'h9d))
                    begin
                      reg731 <= $unsigned((((reg726 ?
                              reg636 : reg725) <= $signed(forvar703)) ?
                          $unsigned((reg716 == (8'ha0))) : $unsigned({forvar682})));
                      reg732 <= (~^((^~(~^forvar726)) ^ $signed((reg716 ?
                          forvar701 : forvar642))));
                    end
                  else
                    begin
                      reg731 <= wire632[(2'h2):(1'h0)];
                      reg732 <= $unsigned($signed({$signed(reg687)}));
                    end
                  for (forvar733 = (1'h0); (forvar733 < (2'h2)); forvar733 = (forvar733 + (1'h1)))
                    begin
                      reg734 <= reg715;
                    end
                  for (forvar735 = (1'h0); (forvar735 < (2'h3)); forvar735 = (forvar735 + (1'h1)))
                    begin
                      reg736 <= reg659[(3'h5):(3'h4)];
                    end
                  if ((reg639 ? reg666 : $signed((|$signed(forvar735)))))
                    begin
                      reg737 <= $signed(($unsigned((reg715 - reg648)) << ($unsigned((8'haf)) ?
                          reg636 : (reg724 ^ reg648))));
                    end
                  else
                    begin
                      reg737 <= forvar637;
                      reg738 <= reg662;
                    end
                end
            end
          else
            begin
              if ((({(reg697 ?
                          reg721 : forvar704)} - ($signed(reg713) >>> {reg717})) ?
                  {$unsigned((8'ha9))} : (^reg734)))
                begin
                  for (forvar716 = (1'h0); (forvar716 < (2'h2)); forvar716 = (forvar716 + (1'h1)))
                    begin
                      reg717 <= $unsigned(wire3);
                      reg718 <= (reg680 ^ (|(8'hab)));
                    end
                  reg719 <= {(((-(8'ha7)) == $signed(reg638)) | reg651[(3'h5):(2'h3)])};
                  reg720 <= $signed(reg734);
                  for (forvar721 = (1'h0); (forvar721 < (1'h1)); forvar721 = (forvar721 + (1'h1)))
                    begin
                      reg722 <= forvar695;
                      reg723 <= $unsigned(((^~{reg702}) ~^ (+(reg714 ?
                          reg712 : reg709))));
                    end
                end
              else
                begin
                  reg716 <= reg715;
                  if ($unsigned({(reg699[(2'h3):(1'h0)] >> $unsigned(reg730))}))
                    begin
                      reg717 <= $signed($signed(reg677));
                      reg718 <= wire4;
                    end
                  else
                    begin
                      reg717 <= ($signed(reg644[(3'h4):(1'h0)]) ^ $unsigned(forvar695));
                      reg718 <= ({$unsigned({reg652})} ^~ (((reg651 ?
                          forvar633 : wire629) & reg734[(1'h1):(1'h1)]) ^~ reg724));
                    end
                  reg719 <= (($unsigned((wire629 * reg698)) ?
                      reg698[(4'hd):(3'h7)] : (!(8'h9c))) < (^reg715[(4'ha):(1'h1)]));
                  reg720 <= (-forvar642[(3'h6):(3'h4)]);
                end
            end
        end
    end
  module739 #() modinst1087 (wire1086, clk, reg681, reg704, reg716, reg665);
  assign wire1088 = {($unsigned(reg692[(3'h4):(3'h4)]) ?
                            {(~^reg690)} : $signed({reg689}))};
  always
    @(posedge clk) begin
      if (reg707)
        begin
          if (reg717[(3'h6):(1'h0)])
            begin
              reg1089 <= {reg738};
              if ($unsigned(reg730))
                begin
                  reg1090 <= {(^{reg661[(3'h5):(1'h0)]})};
                  for (forvar1091 = (1'h0); (forvar1091 < (1'h1)); forvar1091 = (forvar1091 + (1'h1)))
                    begin
                      reg1092 <= $unsigned(reg668[(1'h0):(1'h0)]);
                      reg1093 <= (!$signed(reg738[(4'hc):(4'h8)]));
                    end
                  for (forvar1094 = (1'h0); (forvar1094 < (2'h3)); forvar1094 = (forvar1094 + (1'h1)))
                    begin
                      reg1095 <= {reg641};
                      reg1096 <= reg738[(4'hb):(2'h3)];
                      reg1097 <= {((wire1086[(3'h5):(3'h4)] ?
                              (reg676 || (8'had)) : (+reg654)) ^~ {(wire2 >> reg665)})};
                      reg1098 <= (8'hb9);
                    end
                  for (forvar1099 = (1'h0); (forvar1099 < (2'h3)); forvar1099 = (forvar1099 + (1'h1)))
                    begin
                      reg1100 <= ($signed(reg724) >>> $signed(reg722));
                    end
                end
              else
                begin
                  if (reg736[(1'h1):(1'h0)])
                    begin
                      reg1090 <= $unsigned($signed(($signed(reg729) ^ $signed(forvar1091))));
                      reg1091 <= $signed($signed($signed((8'hae))));
                      reg1092 <= ($signed((reg685[(2'h3):(1'h0)] << $signed(reg728))) >>> $signed(reg729));
                    end
                  else
                    begin
                      reg1090 <= reg683[(1'h1):(1'h0)];
                    end
                end
            end
          else
            begin
              if (((($unsigned(reg726) ? (reg694 + reg726) : (-(8'hb2))) ?
                  reg655 : ((reg690 ?
                      reg723 : (8'ha6)) <= {reg667})) > ({$signed(reg736)} ^ (reg655[(3'h7):(3'h4)] <<< reg726[(3'h4):(2'h3)]))))
                begin
                  if ($unsigned(($signed((&(8'h9c))) ?
                      reg699[(4'hf):(1'h0)] : (|forvar1091[(1'h0):(1'h0)]))))
                    begin
                      reg1089 <= {((reg726[(3'h6):(2'h2)] >> (reg716 < reg652)) || ({reg725} >> $unsigned(reg667)))};
                      reg1090 <= reg650[(3'h4):(3'h4)];
                      reg1091 <= ({(((8'ha8) ? reg730 : reg706) ?
                              wire4[(3'h6):(3'h6)] : $signed(reg698))} + ((~|(!reg693)) && ((-(8'had)) << (&reg704))));
                    end
                  else
                    begin
                      reg1089 <= reg690;
                      reg1090 <= (~^(reg644 >= reg726));
                    end
                  if ((8'hb2))
                    begin
                      reg1092 <= {(reg702 != ({reg734} ?
                              (reg718 ?
                                  (8'h9c) : (8'h9c)) : (reg1093 && reg638)))};
                      reg1093 <= reg646;
                      reg1094 <= $signed(($signed(reg723) ?
                          (~^(+(8'hb7))) : (reg669 == reg701)));
                    end
                  else
                    begin
                      reg1092 <= reg653[(3'h4):(2'h3)];
                      reg1093 <= ($unsigned({reg724}) ?
                          ((~{reg1093}) ?
                              (reg687 > reg641) : $unsigned(reg679)) : (wire1[(3'h5):(2'h2)] ^ (|$unsigned(reg663))));
                      reg1094 <= reg699[(4'hf):(3'h7)];
                      reg1095 <= $unsigned($signed($unsigned((&reg687))));
                    end
                  if ((!reg649))
                    begin
                      reg1096 <= (reg736[(2'h2):(1'h1)] ?
                          $signed((~|reg728)) : ((|reg725) ?
                              reg655 : (wire0[(4'hd):(1'h0)] ~^ {reg647})));
                      reg1097 <= $unsigned(reg702);
                      reg1098 <= reg647;
                      reg1099 <= reg636[(3'h6):(1'h0)];
                    end
                  else
                    begin
                      reg1096 <= (8'haf);
                      reg1097 <= (+$signed((~(8'hb3))));
                      reg1098 <= $unsigned(reg638[(3'h6):(1'h1)]);
                    end
                end
              else
                begin
                  reg1089 <= (8'hb5);
                  for (forvar1090 = (1'h0); (forvar1090 < (1'h1)); forvar1090 = (forvar1090 + (1'h1)))
                    begin
                      reg1091 <= ((wire3[(3'h4):(3'h4)] * (-reg685[(4'h8):(3'h7)])) ?
                          (((reg702 && reg731) ^ reg703) ?
                              ($unsigned(reg724) ?
                                  (reg645 ?
                                      reg694 : reg689) : {reg1097}) : wire629) : $signed(reg707));
                      reg1092 <= (8'hb6);
                      reg1093 <= {($unsigned(((8'ha7) < reg685)) ?
                              reg654[(2'h3):(1'h0)] : ((wire629 >> reg685) ?
                                  $unsigned((8'ha3)) : {reg684}))};
                    end
                end
            end
          reg1101 <= ((reg643[(3'h7):(3'h5)] != (-$signed(reg639))) << (&reg713));
          if (reg683[(1'h0):(1'h0)])
            begin
              if (forvar1099)
                begin
                  if (reg683[(1'h0):(1'h0)])
                    begin
                      reg1102 <= {(|(+((8'ha8) ? reg717 : reg723)))};
                      reg1103 <= reg671[(4'h8):(2'h3)];
                    end
                  else
                    begin
                      reg1102 <= $unsigned(((+$signed(reg641)) | ($signed(reg699) * $unsigned((8'ha3)))));
                      reg1103 <= $signed({{$signed(reg707)}});
                      reg1104 <= ($signed($unsigned($unsigned(reg667))) ?
                          $unsigned(reg674[(3'h6):(3'h4)]) : $unsigned($signed(reg659[(3'h5):(3'h4)])));
                      reg1105 <= wire629;
                    end
                end
              else
                begin
                  reg1102 <= ($unsigned(($signed(reg1098) ?
                          (reg718 ? reg1089 : reg704) : {reg733})) ?
                      ($unsigned((reg662 ^ reg724)) ^~ wire1088[(2'h2):(1'h0)]) : (8'hb2));
                  reg1103 <= (reg723[(2'h2):(1'h1)] << $signed((8'hb6)));
                  reg1104 <= $signed($signed((^(-reg634))));
                  if ({$unsigned((reg717 ? (reg1097 & reg727) : {reg711}))})
                    begin
                      reg1105 <= reg714[(3'h4):(2'h3)];
                      reg1106 <= reg1092;
                      reg1107 <= ((($unsigned(reg644) ?
                              (reg719 ? reg667 : reg668) : (reg694 ?
                                  reg659 : reg657)) - reg676[(1'h0):(1'h0)]) ?
                          reg737 : ((~reg675) + $unsigned((reg676 ?
                              (8'hb4) : reg667))));
                      reg1108 <= {$signed(((reg1096 ?
                              reg635 : reg1094) & reg731))};
                    end
                  else
                    begin
                      reg1105 <= {(^~(^reg1089))};
                      reg1106 <= (~(forvar1094[(2'h3):(2'h2)] ?
                          reg731[(2'h2):(2'h2)] : (-$unsigned((8'ha3)))));
                      reg1107 <= (8'ha2);
                    end
                end
            end
          else
            begin
              for (forvar1102 = (1'h0); (forvar1102 < (1'h1)); forvar1102 = (forvar1102 + (1'h1)))
                begin
                  for (forvar1103 = (1'h0); (forvar1103 < (1'h1)); forvar1103 = (forvar1103 + (1'h1)))
                    begin
                      reg1104 <= (($unsigned((-reg657)) * $signed($unsigned(reg1093))) * (^~({reg681} ?
                          $unsigned(reg696) : (^~reg653))));
                      reg1105 <= (reg698 * $unsigned(reg645));
                      reg1106 <= (~^(~|($signed(reg668) ^ (reg1096 && forvar1094))));
                    end
                end
              for (forvar1107 = (1'h0); (forvar1107 < (2'h3)); forvar1107 = (forvar1107 + (1'h1)))
                begin
                  for (forvar1108 = (1'h0); (forvar1108 < (2'h3)); forvar1108 = (forvar1108 + (1'h1)))
                    begin
                      reg1109 <= ((((reg713 && reg1108) || (reg680 ?
                          reg676 : reg690)) & ((~|reg702) ?
                          $signed(reg657) : (|reg738))) >>> reg662);
                    end
                  if ((reg1093 ?
                      reg653 : (reg690[(1'h0):(1'h0)] ?
                          $signed({reg1093}) : ($signed(forvar1103) ?
                              $unsigned(reg1097) : (reg709 ?
                                  wire1086 : reg666)))))
                    begin
                      reg1110 <= reg1104;
                      reg1111 <= ((^$unsigned($signed(reg717))) - ({reg650} ?
                          reg1092 : (reg696 & reg687[(3'h4):(2'h2)])));
                      reg1112 <= (~|forvar1091[(1'h1):(1'h0)]);
                      reg1113 <= $unsigned($unsigned(reg636));
                    end
                  else
                    begin
                      reg1110 <= (8'h9e);
                      reg1111 <= reg723[(2'h2):(1'h1)];
                      reg1112 <= ($unsigned((reg727 >> {reg1105})) >>> (&$unsigned(((8'ha9) ?
                          reg706 : reg657))));
                      reg1113 <= reg730[(2'h3):(2'h2)];
                    end
                end
              reg1114 <= wire631[(3'h6):(3'h4)];
              if (reg684[(3'h6):(2'h2)])
                begin
                  for (forvar1115 = (1'h0); (forvar1115 < (2'h3)); forvar1115 = (forvar1115 + (1'h1)))
                    begin
                      reg1116 <= (reg662 <= $unsigned((!$signed(reg659))));
                      reg1117 <= reg687[(3'h4):(1'h1)];
                      reg1118 <= ($unsigned(reg1113) ^ $unsigned((reg638[(1'h0):(1'h0)] ?
                          (forvar1115 ? wire1 : reg709) : {reg732})));
                    end
                  reg1119 <= reg689;
                  for (forvar1120 = (1'h0); (forvar1120 < (2'h2)); forvar1120 = (forvar1120 + (1'h1)))
                    begin
                      reg1121 <= ({(((8'ha2) ? wire1 : reg654) >> {reg716})} ?
                          ($signed(reg654) ?
                              {{reg653}} : (reg647 ?
                                  forvar1099 : (reg659 ?
                                      wire0 : (8'hb9)))) : $signed($signed({reg653})));
                      reg1122 <= ($signed($signed(reg634)) ?
                          $unsigned(reg1107[(3'h4):(1'h1)]) : (+($signed(forvar1107) >>> reg1114)));
                    end
                  if (wire2[(4'he):(1'h0)])
                    begin
                      reg1123 <= forvar1094[(1'h0):(1'h0)];
                      reg1124 <= $unsigned((~(~^reg1093)));
                      reg1125 <= (($signed($signed(reg1111)) ?
                              $unsigned(reg696) : $signed($signed(wire1))) ?
                          (reg702[(3'h6):(2'h2)] ?
                              reg637[(3'h5):(2'h2)] : {$signed((8'hb1))}) : (((reg654 + reg722) == {reg663}) << ((reg669 ?
                                  reg637 : reg1089) ?
                              ((8'ha2) > reg1093) : reg640)));
                      reg1126 <= reg1093;
                    end
                  else
                    begin
                      reg1123 <= (~(((reg634 + reg656) && (reg729 ?
                              reg688 : (8'ha5))) ?
                          (~&$signed(forvar1108)) : (reg731[(1'h1):(1'h1)] >>> reg653[(3'h5):(2'h2)])));
                    end
                end
              else
                begin
                  for (forvar1115 = (1'h0); (forvar1115 < (1'h1)); forvar1115 = (forvar1115 + (1'h1)))
                    begin
                      reg1116 <= ((($signed(reg691) + (~&(8'ha6))) << $signed((~&wire1))) ^ $signed((-{reg713})));
                      reg1117 <= {{(|((8'ha3) << reg664))}};
                    end
                  if ({{reg650}})
                    begin
                      reg1118 <= $signed((!$signed($unsigned(reg1123))));
                      reg1119 <= ({$unsigned(reg684)} << $unsigned(reg714[(3'h5):(2'h3)]));
                      reg1120 <= reg696;
                      reg1121 <= ((^~$unsigned({reg689})) ?
                          reg708[(4'h9):(2'h3)] : reg1118[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1118 <= reg692;
                      reg1119 <= $unsigned((|reg732[(1'h0):(1'h0)]));
                    end
                  for (forvar1122 = (1'h0); (forvar1122 < (2'h3)); forvar1122 = (forvar1122 + (1'h1)))
                    begin
                      reg1123 <= (wire4[(3'h4):(2'h3)] ?
                          ((^((8'hb1) == wire4)) ?
                              (~|$signed(reg651)) : $unsigned($unsigned(reg641))) : $unsigned(reg724[(2'h3):(1'h1)]));
                      reg1124 <= $unsigned(((^~((8'had) ? reg704 : wire632)) ?
                          reg708[(3'h4):(3'h4)] : ($unsigned(reg715) & $signed(reg1092))));
                      reg1125 <= ($unsigned((~|$unsigned(wire631))) ?
                          $unsigned($signed((~|reg1092))) : $signed(wire631));
                    end
                end
            end
          reg1127 <= (+reg696[(5'h10):(4'hf)]);
        end
      else
        begin
          for (forvar1089 = (1'h0); (forvar1089 < (1'h1)); forvar1089 = (forvar1089 + (1'h1)))
            begin
              for (forvar1090 = (1'h0); (forvar1090 < (2'h2)); forvar1090 = (forvar1090 + (1'h1)))
                begin
                  if ($signed($unsigned((reg697 || (!reg1109)))))
                    begin
                      reg1091 <= (reg711[(2'h3):(1'h1)] != reg730[(3'h4):(2'h3)]);
                      reg1092 <= ($signed((^reg1101[(4'hb):(4'hb)])) ?
                          wire2 : forvar1094[(4'hc):(1'h0)]);
                      reg1093 <= ((+reg722[(2'h3):(2'h2)]) * wire3);
                    end
                  else
                    begin
                      reg1091 <= $signed(reg687[(3'h4):(1'h1)]);
                      reg1092 <= reg696;
                      reg1093 <= (($signed(reg636) > ($unsigned(reg687) ?
                          (^reg1106) : $unsigned(reg684))) <<< (((~&reg727) ?
                          $signed((8'hb5)) : $signed(forvar1089)) | ($signed((8'haa)) >>> (^reg1105))));
                    end
                end
              for (forvar1094 = (1'h0); (forvar1094 < (1'h1)); forvar1094 = (forvar1094 + (1'h1)))
                begin
                  if (((~|reg1123[(4'hb):(4'hb)]) ?
                      ({reg1120[(3'h5):(1'h1)]} ?
                          ({(8'ha5)} ?
                              $signed(forvar1115) : $unsigned(reg646)) : ((!reg676) * $signed(reg1105))) : (({reg1113} << (reg657 < (8'hb7))) ?
                          {reg661} : $signed((~^reg659)))))
                    begin
                      reg1095 <= reg707[(2'h2):(2'h2)];
                      reg1096 <= {$signed((reg678 + reg707))};
                      reg1097 <= $signed(reg638[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1095 <= (^~reg668[(1'h0):(1'h0)]);
                      reg1096 <= {{{(reg699 ^ reg727)}}};
                      reg1097 <= ($signed((8'ha5)) >= $unsigned($unsigned($signed(reg1120))));
                    end
                  if (forvar1099[(1'h1):(1'h0)])
                    begin
                      reg1098 <= $signed(({reg645[(1'h1):(1'h0)]} - {$unsigned((8'ha8))}));
                    end
                  else
                    begin
                      reg1098 <= ((({reg736} + {forvar1103}) ?
                          reg685[(1'h1):(1'h0)] : ((reg734 ?
                              reg1106 : reg727) >> $unsigned(reg683))) == $unsigned(((reg692 >>> reg707) ?
                          (reg671 <<< reg637) : ((8'ha7) ?
                              forvar1089 : reg1095))));
                    end
                  if ((8'ha7))
                    begin
                      reg1099 <= (reg715 ?
                          $unsigned($unsigned((8'ha7))) : $unsigned($unsigned($unsigned((8'hb7)))));
                      reg1100 <= $unsigned($signed(forvar1108[(2'h2):(1'h0)]));
                      reg1101 <= {reg725[(4'h9):(2'h3)]};
                      reg1102 <= ($unsigned({(8'haf)}) ?
                          ($signed(reg1111) && $signed(reg664)) : $signed($unsigned({reg1089})));
                    end
                  else
                    begin
                      reg1099 <= reg638[(3'h6):(1'h1)];
                      reg1100 <= (-$unsigned(($signed(reg1094) ?
                          (reg723 ? reg667 : reg681) : $unsigned(reg1099))));
                    end
                  if (reg670[(2'h3):(2'h2)])
                    begin
                      reg1103 <= $unsigned((&(~(reg1098 ? reg705 : reg655))));
                      reg1104 <= (reg640[(2'h2):(1'h1)] ?
                          reg1127[(4'h8):(3'h6)] : {((wire1086 ?
                                      reg683 : (8'hb5)) ?
                                  wire1[(4'h8):(1'h1)] : (reg698 >>> (8'haa)))});
                    end
                  else
                    begin
                      reg1103 <= ((^~((reg647 ?
                              reg1110 : reg1091) ~^ $signed(reg1093))) ?
                          (+(reg720 <<< (reg736 ?
                              reg1120 : (8'ha3)))) : reg698[(4'he):(3'h4)]);
                      reg1104 <= reg1107;
                      reg1105 <= $unsigned((^~($signed((8'hab)) | reg1097)));
                      reg1106 <= ({(^$signed(reg685))} ?
                          {(~(reg651 ? (8'haf) : reg703))} : (((reg634 ?
                              (8'had) : reg635) & wire1086) <<< $signed((wire631 ?
                              (8'h9f) : reg694))));
                    end
                end
              for (forvar1107 = (1'h0); (forvar1107 < (2'h2)); forvar1107 = (forvar1107 + (1'h1)))
                begin
                  if (((&reg701[(1'h0):(1'h0)]) ?
                      reg645[(1'h1):(1'h0)] : {($unsigned((8'hab)) <= ((8'hac) ?
                              reg1102 : reg1098))}))
                    begin
                      reg1108 <= (~(reg653 ?
                          (forvar1094 ? (8'hab) : reg727) : reg643));
                    end
                  else
                    begin
                      reg1108 <= $signed((reg1109 ?
                          ((forvar1102 ^ reg689) & (reg637 ?
                              reg701 : (8'ha1))) : (|((8'ha4) ?
                              reg1104 : reg702))));
                      reg1109 <= ({($signed(reg1119) - $signed(reg730))} < reg657[(3'h7):(3'h4)]);
                    end
                  for (forvar1110 = (1'h0); (forvar1110 < (1'h1)); forvar1110 = (forvar1110 + (1'h1)))
                    begin
                      reg1111 <= $unsigned($unsigned($unsigned((reg1117 ?
                          reg709 : reg1105))));
                    end
                  for (forvar1112 = (1'h0); (forvar1112 < (2'h3)); forvar1112 = (forvar1112 + (1'h1)))
                    begin
                      reg1113 <= $signed((reg1126[(1'h1):(1'h1)] ?
                          reg728[(1'h1):(1'h0)] : (^~(reg1113 ?
                              (8'ha5) : (8'hb4)))));
                      reg1114 <= {reg652[(4'h8):(4'h8)]};
                    end
                  if ({{reg733[(4'ha):(4'h9)]}})
                    begin
                      reg1115 <= reg1104[(1'h1):(1'h0)];
                      reg1116 <= $unsigned(($signed($unsigned(reg669)) ^~ ($unsigned(reg712) ?
                          reg738[(3'h7):(1'h1)] : ((8'hb8) || (8'ha6)))));
                      reg1117 <= {reg1116};
                      reg1118 <= $signed({$signed(reg1092)});
                    end
                  else
                    begin
                      reg1115 <= $signed(reg676);
                      reg1116 <= $signed((8'ha0));
                    end
                end
            end
          reg1119 <= $unsigned((|(forvar1110 ?
              (reg646 ? wire1086 : (8'ha4)) : (reg1102 & reg1113))));
          for (forvar1120 = (1'h0); (forvar1120 < (2'h2)); forvar1120 = (forvar1120 + (1'h1)))
            begin
              if ({({reg654[(2'h2):(1'h0)]} ?
                      $signed((reg643 ?
                          (8'ha0) : reg707)) : $signed($unsigned((8'ha9))))})
                begin
                  for (forvar1121 = (1'h0); (forvar1121 < (1'h0)); forvar1121 = (forvar1121 + (1'h1)))
                    begin
                      reg1122 <= $unsigned(reg712[(4'he):(3'h4)]);
                    end
                  if ($unsigned($signed((((8'hb3) - reg1121) * (|reg722)))))
                    begin
                      reg1123 <= (~|wire3);
                      reg1124 <= (wire2[(1'h1):(1'h0)] <<< reg664[(3'h4):(2'h3)]);
                      reg1125 <= ($signed(((~^reg1110) ^~ $signed(reg1127))) & (reg1091[(1'h0):(1'h0)] ?
                          ((+reg738) | (reg697 >>> reg695)) : $unsigned((~^(8'hb6)))));
                    end
                  else
                    begin
                      reg1123 <= $unsigned(($unsigned(reg657[(1'h0):(1'h0)]) << ((reg1109 ?
                              reg715 : (8'hb8)) ?
                          {wire1088} : ((8'ha5) ? reg1089 : reg1115))));
                    end
                  for (forvar1126 = (1'h0); (forvar1126 < (2'h2)); forvar1126 = (forvar1126 + (1'h1)))
                    begin
                      reg1127 <= $unsigned(((~^$signed((8'ha7))) ?
                          reg654 : ((reg640 ? reg725 : reg725) || (reg698 ?
                              reg637 : reg658))));
                    end
                end
              else
                begin
                  for (forvar1121 = (1'h0); (forvar1121 < (1'h0)); forvar1121 = (forvar1121 + (1'h1)))
                    begin
                      reg1122 <= forvar1091;
                      reg1123 <= ($signed(forvar1090) <<< {(wire1086 > {reg649})});
                      reg1124 <= $unsigned(($unsigned($signed((8'haa))) ?
                          (-reg658) : {(+reg659)}));
                    end
                end
              reg1128 <= $signed((~|((reg1117 ? reg654 : (8'hb6)) ?
                  reg649 : (reg678 ? reg1115 : reg675))));
              for (forvar1129 = (1'h0); (forvar1129 < (2'h2)); forvar1129 = (forvar1129 + (1'h1)))
                begin
                  if ((forvar1115[(3'h7):(1'h1)] < (^~$unsigned($signed(reg1121)))))
                    begin
                      reg1130 <= $signed(reg714);
                    end
                  else
                    begin
                      reg1130 <= (&($unsigned((^~reg707)) | $unsigned((&(8'hae)))));
                      reg1131 <= ($signed((reg1091[(4'he):(4'hb)] ?
                              (reg719 & reg732) : reg722[(1'h0):(1'h0)])) ?
                          {$unsigned({(8'ha2)})} : wire1086);
                      reg1132 <= (+$signed(reg677[(1'h1):(1'h0)]));
                    end
                  for (forvar1133 = (1'h0); (forvar1133 < (2'h2)); forvar1133 = (forvar1133 + (1'h1)))
                    begin
                      reg1134 <= $unsigned((reg668 ?
                          (((8'hb9) & reg643) ?
                              {reg655} : $unsigned((8'hb8))) : ((wire0 == (8'h9e)) <= reg640[(4'h9):(1'h1)])));
                      reg1135 <= (((8'hac) ?
                          reg653 : $unsigned(reg1091[(4'h8):(2'h2)])) > ($signed({(8'ha4)}) ?
                          reg657[(3'h4):(1'h0)] : $signed(reg711[(1'h0):(1'h0)])));
                      reg1136 <= (8'hb4);
                    end
                end
            end
        end
      for (forvar1137 = (1'h0); (forvar1137 < (2'h3)); forvar1137 = (forvar1137 + (1'h1)))
        begin
          for (forvar1138 = (1'h0); (forvar1138 < (1'h1)); forvar1138 = (forvar1138 + (1'h1)))
            begin
              for (forvar1139 = (1'h0); (forvar1139 < (2'h2)); forvar1139 = (forvar1139 + (1'h1)))
                begin
                  reg1140 <= reg646;
                  for (forvar1141 = (1'h0); (forvar1141 < (2'h2)); forvar1141 = (forvar1141 + (1'h1)))
                    begin
                      reg1142 <= $signed(((~&reg675) >> ((reg720 * reg641) <<< {reg662})));
                      reg1143 <= {$signed(reg641)};
                      reg1144 <= $signed(((^reg704) ?
                          ($unsigned(reg690) ?
                              (reg683 || reg737) : (^~(8'hb2))) : reg1143));
                    end
                end
              if ({$signed(reg1132)})
                begin
                  for (forvar1145 = (1'h0); (forvar1145 < (1'h0)); forvar1145 = (forvar1145 + (1'h1)))
                    begin
                      reg1146 <= $signed({(8'had)});
                      reg1147 <= ({$unsigned((-reg1110))} - reg1121[(2'h3):(1'h1)]);
                      reg1148 <= $signed($signed($unsigned({reg675})));
                      reg1149 <= $signed(((~|(reg655 ? reg1132 : reg1101)) ?
                          $unsigned($unsigned(forvar1091)) : wire632[(3'h6):(2'h2)]));
                    end
                  for (forvar1150 = (1'h0); (forvar1150 < (1'h1)); forvar1150 = (forvar1150 + (1'h1)))
                    begin
                      reg1151 <= reg712[(4'he):(2'h3)];
                      reg1152 <= ((reg699 || ({forvar1107} ?
                              ((8'ha8) & forvar1091) : reg719)) ?
                          $unsigned((~|(reg1134 > reg1115))) : $unsigned(reg658[(4'h8):(3'h7)]));
                      reg1153 <= (8'haa);
                      reg1154 <= reg721;
                    end
                end
              else
                begin
                  for (forvar1145 = (1'h0); (forvar1145 < (1'h1)); forvar1145 = (forvar1145 + (1'h1)))
                    begin
                      reg1146 <= $unsigned(reg1127[(1'h1):(1'h1)]);
                      reg1147 <= ({{reg738}} ?
                          $signed(((reg676 ? (8'ha3) : wire1088) ?
                              reg1095 : (~reg702))) : (!$unsigned({(8'ha7)})));
                      reg1148 <= $signed($unsigned((^reg707[(1'h0):(1'h0)])));
                      reg1149 <= ((({reg738} < reg639[(3'h5):(2'h2)]) ?
                              reg1143 : (|(forvar1145 << reg671))) ?
                          $unsigned((+reg675[(4'h8):(3'h6)])) : ($unsigned(reg642) ?
                              $unsigned(reg683) : reg693[(3'h7):(3'h5)]));
                    end
                end
            end
          for (forvar1155 = (1'h0); (forvar1155 < (1'h0)); forvar1155 = (forvar1155 + (1'h1)))
            begin
              for (forvar1156 = (1'h0); (forvar1156 < (1'h0)); forvar1156 = (forvar1156 + (1'h1)))
                begin
                  for (forvar1157 = (1'h0); (forvar1157 < (1'h0)); forvar1157 = (forvar1157 + (1'h1)))
                    begin
                      reg1158 <= (reg1134 ?
                          $unsigned($signed({reg662})) : reg1126[(1'h1):(1'h0)]);
                      reg1159 <= $unsigned(reg1125);
                      reg1160 <= reg669;
                      reg1161 <= $signed($signed($unsigned({(8'hae)})));
                    end
                end
            end
        end
      for (forvar1162 = (1'h0); (forvar1162 < (1'h0)); forvar1162 = (forvar1162 + (1'h1)))
        begin
          for (forvar1163 = (1'h0); (forvar1163 < (2'h3)); forvar1163 = (forvar1163 + (1'h1)))
            begin
              for (forvar1164 = (1'h0); (forvar1164 < (2'h3)); forvar1164 = (forvar1164 + (1'h1)))
                begin
                  if ($unsigned((+reg638)))
                    begin
                      reg1165 <= {reg679[(2'h3):(2'h2)]};
                      reg1166 <= (($unsigned((~&reg726)) ?
                              ((reg737 ?
                                  forvar1099 : reg711) == (forvar1121 << reg676)) : {$unsigned(forvar1102)}) ?
                          ((^(wire1086 ?
                              reg1152 : reg736)) & $unsigned((~&wire1086))) : (forvar1122 ?
                              (~^(~(8'hb8))) : wire4));
                      reg1167 <= $signed(reg1144);
                      reg1168 <= reg703;
                    end
                  else
                    begin
                      reg1165 <= ($unsigned($signed((&reg1120))) | (reg1108 ^ ($unsigned(reg656) == (8'h9d))));
                    end
                  for (forvar1169 = (1'h0); (forvar1169 < (1'h1)); forvar1169 = (forvar1169 + (1'h1)))
                    begin
                      reg1170 <= ($signed($signed(reg1099)) ?
                          ((reg722[(1'h0):(1'h0)] >> $signed(forvar1150)) ?
                              {{(8'hac)}} : (~|(reg1158 ?
                                  reg722 : forvar1133))) : $unsigned(reg637));
                    end
                end
            end
        end
    end
  module1171 #() modinst1754 (wire1753, clk, reg659, reg1110, reg1151, reg664, reg647);
  always
    @(posedge clk) begin
      for (forvar1755 = (1'h0); (forvar1755 < (2'h2)); forvar1755 = (forvar1755 + (1'h1)))
        begin
          if (((~($signed((8'ha0)) ?
              (8'hb0) : (reg634 || reg1167))) >= ({(reg675 - (8'ha4))} > $unsigned({reg1170}))))
            begin
              for (forvar1756 = (1'h0); (forvar1756 < (1'h0)); forvar1756 = (forvar1756 + (1'h1)))
                begin
                  reg1757 <= $unsigned(reg680);
                  reg1758 <= forvar1756;
                  for (forvar1759 = (1'h0); (forvar1759 < (1'h1)); forvar1759 = (forvar1759 + (1'h1)))
                    begin
                      reg1760 <= $signed((~$unsigned(reg691[(2'h2):(1'h1)])));
                    end
                  reg1761 <= ($unsigned({$signed((8'haf))}) ?
                      (($signed(reg646) ?
                          {(8'hba)} : reg1131) != $signed((+reg736))) : $signed(reg696));
                end
              if ($signed((~&((reg1107 ~^ reg1108) & (reg1118 ?
                  reg715 : (8'haa))))))
                begin
                  for (forvar1762 = (1'h0); (forvar1762 < (1'h1)); forvar1762 = (forvar1762 + (1'h1)))
                    begin
                      reg1763 <= ((($unsigned(reg722) ?
                          $signed(reg641) : (8'ha7)) + (8'hb6)) | (~|(~|$unsigned((8'h9c)))));
                      reg1764 <= (reg1109[(2'h3):(2'h2)] != reg1109[(1'h1):(1'h1)]);
                      reg1765 <= $unsigned((~$unsigned($signed(reg668))));
                      reg1766 <= $unsigned(reg1098);
                    end
                  if (((($unsigned(reg1143) ? (~^reg733) : $signed((8'hb4))) ?
                          $signed((8'hb3)) : ($unsigned(reg662) ?
                              reg1128 : $unsigned(reg1100))) ?
                      $signed((((8'hb0) ? reg1160 : (8'ha7)) ?
                          reg1100[(4'ha):(4'h8)] : (~^reg1121))) : reg1159))
                    begin
                      reg1767 <= wire2;
                    end
                  else
                    begin
                      reg1767 <= reg730[(1'h1):(1'h0)];
                    end
                  for (forvar1768 = (1'h0); (forvar1768 < (1'h1)); forvar1768 = (forvar1768 + (1'h1)))
                    begin
                      reg1769 <= reg651;
                      reg1770 <= {((reg1097[(1'h0):(1'h0)] < reg671) ?
                              reg1098 : $signed($unsigned(reg1091)))};
                    end
                end
              else
                begin
                  if ((reg708[(3'h5):(2'h2)] || reg712))
                    begin
                      reg1762 <= $unsigned(reg663);
                      reg1763 <= $signed($unsigned(((reg680 | wire1753) ?
                          {reg1125} : (8'hb1))));
                      reg1764 <= (~^reg651);
                      reg1765 <= (($signed((+(8'hae))) == (~&(~&(8'ha8)))) ?
                          (~^(~|(8'h9f))) : ($unsigned(((8'hac) <<< reg664)) ?
                              (8'had) : ($unsigned(reg697) < (reg1092 >>> reg662))));
                    end
                  else
                    begin
                      reg1762 <= $unsigned((~^(reg656 ?
                          $unsigned(reg1769) : {reg734})));
                      reg1763 <= (|($signed($unsigned(reg694)) ?
                          $unsigned({reg1117}) : reg661[(3'h5):(3'h5)]));
                    end
                end
              if ((wire629[(3'h5):(1'h1)] ?
                  (+reg1764) : $unsigned($unsigned((reg695 ?
                      reg1765 : (8'ha3))))))
                begin
                  if ($signed(($unsigned((reg1166 | reg693)) ?
                      $unsigned((8'hb2)) : (~^$signed(reg730)))))
                    begin
                      reg1771 <= $unsigned($signed(((reg1167 <<< reg716) ?
                          (^reg1106) : $unsigned(wire4))));
                      reg1772 <= (reg1153 <<< ($signed((|reg1100)) ?
                          reg724 : {$signed(reg687)}));
                      reg1773 <= reg728;
                    end
                  else
                    begin
                      reg1771 <= $unsigned($signed($unsigned(reg1091)));
                    end
                  reg1774 <= $signed((~(+reg1160)));
                end
              else
                begin
                  reg1771 <= ((~^$signed(reg734)) ?
                      (reg1140 * ($signed(reg1168) <= $signed(wire1086))) : ((^~$signed(wire3)) ?
                          reg1763 : reg664[(2'h2):(1'h0)]));
                end
              reg1775 <= (reg703 ?
                  (reg737[(4'ha):(3'h6)] ?
                      (|(reg644 ?
                          reg1771 : reg1771)) : $signed(reg699[(3'h7):(3'h7)])) : ($signed((wire632 ?
                      reg694 : reg1116)) << ({reg1136} ?
                      $unsigned(reg1120) : ((8'haa) ? reg1766 : reg1132))));
            end
          else
            begin
              for (forvar1756 = (1'h0); (forvar1756 < (2'h2)); forvar1756 = (forvar1756 + (1'h1)))
                begin
                  for (forvar1757 = (1'h0); (forvar1757 < (2'h2)); forvar1757 = (forvar1757 + (1'h1)))
                    begin
                      reg1758 <= $unsigned({reg1127});
                      reg1759 <= ({(reg1140[(4'hf):(4'he)] - reg1154[(1'h0):(1'h0)])} ?
                          (~|$unsigned({reg1115})) : (+$signed($signed(reg1758))));
                      reg1760 <= (^~{$signed($unsigned(reg674))});
                      reg1761 <= ({(~reg1757)} ?
                          (wire631 ?
                              reg1120[(2'h2):(1'h0)] : reg722) : forvar1756[(4'h9):(2'h2)]);
                    end
                  for (forvar1762 = (1'h0); (forvar1762 < (2'h2)); forvar1762 = (forvar1762 + (1'h1)))
                    begin
                      reg1763 <= $signed(reg1108);
                      reg1764 <= (reg639[(3'h4):(1'h0)] >>> $signed((&reg1765[(2'h3):(1'h0)])));
                    end
                  for (forvar1765 = (1'h0); (forvar1765 < (2'h3)); forvar1765 = (forvar1765 + (1'h1)))
                    begin
                      reg1766 <= ((reg647 >= $unsigned($signed(reg1146))) ?
                          reg712 : ((-reg1135[(4'hd):(4'hb)]) << (-$unsigned((8'h9c)))));
                      reg1767 <= ((-{$unsigned(reg1089)}) ?
                          reg1093[(3'h4):(2'h3)] : (8'ha9));
                      reg1768 <= $unsigned($unsigned(((|reg697) ^~ (~&reg729))));
                      reg1769 <= reg1113[(2'h2):(1'h1)];
                    end
                  for (forvar1770 = (1'h0); (forvar1770 < (2'h3)); forvar1770 = (forvar1770 + (1'h1)))
                    begin
                      reg1771 <= $unsigned({$unsigned({(8'hb7)})});
                      reg1772 <= reg643;
                      reg1773 <= (-(8'hae));
                    end
                end
              if (({((reg1758 < wire1086) ?
                      (|reg665) : (reg663 && reg698))} || (reg643 ?
                  reg1118 : reg1126)))
                begin
                  if (($unsigned(($signed(reg1159) * $signed(reg640))) && (reg1149[(3'h6):(3'h5)] - (~^$unsigned(reg689)))))
                    begin
                      reg1774 <= (^~(({reg1127} ?
                              $signed(reg1775) : (^(8'hb0))) ?
                          (reg1142[(2'h2):(2'h2)] < reg703) : ($signed((8'hac)) ?
                              reg1760[(3'h6):(1'h1)] : ((8'h9e) >>> reg1130))));
                    end
                  else
                    begin
                      reg1774 <= reg734;
                      reg1775 <= $unsigned(((reg727 * $unsigned((8'haa))) ?
                          $unsigned($signed(reg723)) : $unsigned((~(8'h9d)))));
                    end
                  if ({reg654[(2'h2):(1'h1)]})
                    begin
                      reg1776 <= $signed((!$signed($unsigned(reg1106))));
                      reg1777 <= reg1095[(4'h8):(4'h8)];
                      reg1778 <= ($unsigned((~(|wire632))) >= ({(reg651 ?
                              reg711 : reg721)} ^~ {$unsigned(reg1104)}));
                    end
                  else
                    begin
                      reg1776 <= reg1147[(1'h1):(1'h0)];
                      reg1777 <= reg647[(4'he):(3'h4)];
                      reg1778 <= reg664[(3'h6):(2'h3)];
                      reg1779 <= $signed(reg1757[(2'h2):(1'h1)]);
                    end
                  if ((&reg1170))
                    begin
                      reg1780 <= ($unsigned({(reg638 ?
                              reg661 : (8'ha6))}) + reg1122[(1'h1):(1'h0)]);
                      reg1781 <= (+{reg1109[(1'h1):(1'h1)]});
                    end
                  else
                    begin
                      reg1780 <= reg1769[(3'h4):(2'h2)];
                      reg1781 <= ($unsigned({reg648[(4'h9):(4'h9)]}) ?
                          $unsigned(forvar1768[(3'h4):(2'h3)]) : (({reg649} ?
                                  (8'h9e) : {reg734}) ?
                              $signed($unsigned(wire632)) : $unsigned((reg1115 ^ (8'hb7)))));
                    end
                end
              else
                begin
                  if ($signed((~|{$unsigned(reg644)})))
                    begin
                      reg1774 <= wire1086[(1'h1):(1'h1)];
                      reg1775 <= reg654;
                      reg1776 <= $signed(($unsigned(reg1134) ?
                          $unsigned($unsigned((8'h9c))) : $unsigned((reg1165 ?
                              (8'hac) : wire3))));
                    end
                  else
                    begin
                      reg1774 <= $signed($signed(($signed(reg1101) ?
                          reg1124[(1'h0):(1'h0)] : {(8'haf)})));
                      reg1775 <= $signed($unsigned((reg1120[(3'h5):(3'h4)] >> (~&reg646))));
                      reg1776 <= reg1093;
                      reg1777 <= $signed(reg660);
                    end
                  for (forvar1778 = (1'h0); (forvar1778 < (2'h3)); forvar1778 = (forvar1778 + (1'h1)))
                    begin
                      reg1779 <= $unsigned($signed($unsigned((~&reg1099))));
                      reg1780 <= (&$unsigned($signed($unsigned(reg679))));
                      reg1781 <= ((^{{reg667}}) ?
                          $unsigned($unsigned($signed(reg1124))) : $signed(reg1131));
                    end
                  if ($signed(((reg646 ?
                          (reg641 ? reg707 : reg683) : ((8'had) ?
                              reg652 : reg727)) ?
                      $unsigned(reg1124[(2'h2):(2'h2)]) : $unsigned((reg656 >>> reg1765)))))
                    begin
                      reg1782 <= reg1092;
                      reg1783 <= reg653[(3'h5):(3'h5)];
                      reg1784 <= (({$signed((8'had))} ?
                              $unsigned((reg736 != reg656)) : reg678[(3'h4):(2'h3)]) ?
                          (~&((!reg681) * (reg1122 >= wire1086))) : $unsigned((reg652 && reg1111)));
                      reg1785 <= (^~reg1090[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg1782 <= reg1762;
                      reg1783 <= (^$signed(wire1086));
                      reg1784 <= (-{reg1768});
                    end
                  for (forvar1786 = (1'h0); (forvar1786 < (1'h1)); forvar1786 = (forvar1786 + (1'h1)))
                    begin
                      reg1787 <= $unsigned($signed(($signed((8'ha3)) <= $signed(reg1114))));
                    end
                end
              reg1788 <= ($signed(((reg1096 ~^ (8'hb6)) ?
                      $signed((8'ha1)) : reg1109[(1'h0):(1'h0)])) ?
                  $signed(($signed(forvar1755) ?
                      {reg683} : $unsigned(reg647))) : ((8'h9c) | (~|(reg1779 ?
                      reg718 : wire629))));
            end
          reg1789 <= (($unsigned(reg729[(4'ha):(3'h4)]) == $unsigned((reg1131 ?
              reg728 : reg1765))) - (8'ha8));
          for (forvar1790 = (1'h0); (forvar1790 < (2'h2)); forvar1790 = (forvar1790 + (1'h1)))
            begin
              if ($unsigned(reg657))
                begin
                  if (($unsigned($signed({(8'hb0)})) ?
                      (!(reg1775 & (reg1116 >>> reg659))) : (-$signed((&reg1166)))))
                    begin
                      reg1791 <= reg1773;
                    end
                  else
                    begin
                      reg1791 <= wire4;
                      reg1792 <= {(((!(8'hb1)) > $unsigned(reg666)) ?
                              {(|reg1784)} : ($signed(reg650) ^~ (~|wire629)))};
                      reg1793 <= reg1772[(3'h6):(2'h3)];
                    end
                  if (forvar1768[(3'h5):(2'h3)])
                    begin
                      reg1794 <= (8'hba);
                      reg1795 <= (8'haf);
                      reg1796 <= (((8'hb7) ?
                              $unsigned((reg666 ?
                                  forvar1790 : reg1773)) : {(-forvar1759)}) ?
                          (~(+(reg1119 ^ reg697))) : $signed($unsigned($unsigned(reg1091))));
                    end
                  else
                    begin
                      reg1794 <= $signed(reg635[(3'h5):(3'h5)]);
                      reg1795 <= ({reg693[(4'hb):(4'hb)]} << {$signed($unsigned(reg1112))});
                      reg1796 <= (8'hb1);
                    end
                  for (forvar1797 = (1'h0); (forvar1797 < (1'h1)); forvar1797 = (forvar1797 + (1'h1)))
                    begin
                      reg1798 <= reg664[(3'h6):(2'h3)];
                      reg1799 <= forvar1790[(3'h5):(3'h4)];
                    end
                  for (forvar1800 = (1'h0); (forvar1800 < (2'h3)); forvar1800 = (forvar1800 + (1'h1)))
                    begin
                      reg1801 <= reg1775;
                    end
                end
              else
                begin
                  if (reg1114)
                    begin
                      reg1791 <= $unsigned(((((8'hb4) >= reg663) || (+reg695)) * reg1143[(2'h3):(2'h2)]));
                      reg1792 <= $signed($signed((-(+reg691))));
                    end
                  else
                    begin
                      reg1791 <= reg689[(4'hd):(1'h0)];
                      reg1792 <= {(wire2 && reg1104)};
                      reg1793 <= ($signed({(reg1114 >> (8'ha0))}) <<< (reg703 ?
                          reg677 : (~&reg1781[(3'h6):(2'h3)])));
                    end
                end
              for (forvar1802 = (1'h0); (forvar1802 < (2'h2)); forvar1802 = (forvar1802 + (1'h1)))
                begin
                  if ((-reg1789[(3'h4):(2'h2)]))
                    begin
                      reg1803 <= (8'hb4);
                      reg1804 <= (8'haf);
                      reg1805 <= $signed($signed((!{(8'ha2)})));
                    end
                  else
                    begin
                      reg1803 <= $unsigned(reg713);
                      reg1804 <= wire1[(4'h9):(3'h5)];
                      reg1805 <= {(reg1144 < reg680[(2'h2):(1'h1)])};
                    end
                  if (((((8'ha0) ? (~^reg658) : reg704) ?
                          reg640[(4'hb):(3'h5)] : wire3) ?
                      (^$signed((reg1792 ?
                          reg1154 : reg1804))) : (~|(reg1115[(3'h7):(3'h7)] ^~ $unsigned(reg1111)))))
                    begin
                      reg1806 <= $unsigned(reg675);
                      reg1807 <= (|$unsigned($unsigned((-forvar1802))));
                    end
                  else
                    begin
                      reg1806 <= reg688;
                      reg1807 <= $unsigned({(((8'hb6) - reg1123) ?
                              (reg638 < reg697) : $unsigned(reg719))});
                      reg1808 <= (~^$signed((((8'hb4) ? reg1784 : (8'haf)) ?
                          reg647[(3'h7):(1'h1)] : {reg658})));
                    end
                  reg1809 <= (~&$signed(($unsigned(reg647) > $unsigned(reg1783))));
                  for (forvar1810 = (1'h0); (forvar1810 < (1'h1)); forvar1810 = (forvar1810 + (1'h1)))
                    begin
                      reg1811 <= reg1130[(1'h1):(1'h0)];
                    end
                end
            end
          for (forvar1812 = (1'h0); (forvar1812 < (1'h0)); forvar1812 = (forvar1812 + (1'h1)))
            begin
              if ($signed(((&reg1089[(3'h7):(3'h7)]) ?
                  {$signed(reg683)} : ($unsigned(reg1098) <= (reg635 >> reg679)))))
                begin
                  for (forvar1813 = (1'h0); (forvar1813 < (1'h0)); forvar1813 = (forvar1813 + (1'h1)))
                    begin
                      reg1814 <= (&(($unsigned(reg1787) < {reg1760}) < reg1761));
                    end
                  reg1815 <= $signed(((reg665[(3'h4):(3'h4)] + reg1104[(1'h1):(1'h1)]) ?
                      (8'ha0) : (reg692 * $unsigned(reg722))));
                  reg1816 <= reg1093[(1'h0):(1'h0)];
                end
              else
                begin
                  for (forvar1813 = (1'h0); (forvar1813 < (2'h2)); forvar1813 = (forvar1813 + (1'h1)))
                    begin
                      reg1814 <= (reg1773 >> (reg1125[(4'hd):(4'hb)] << {(8'h9c)}));
                      reg1815 <= $unsigned((^~$signed($signed(reg1123))));
                    end
                  reg1816 <= ((reg1128 - (+(^~reg1806))) ?
                      (reg715 ? reg707 : {reg1109[(1'h0):(1'h0)]}) : reg1135);
                  for (forvar1817 = (1'h0); (forvar1817 < (2'h2)); forvar1817 = (forvar1817 + (1'h1)))
                    begin
                      reg1818 <= $unsigned($unsigned($unsigned($signed(reg654))));
                      reg1819 <= $unsigned(reg1096[(1'h0):(1'h0)]);
                    end
                end
              reg1820 <= (reg1795 ?
                  {$unsigned(reg1109[(2'h3):(1'h0)])} : (|(~&$unsigned(reg1092))));
            end
        end
    end
  assign wire1821 = $unsigned(($unsigned((wire1086 ? reg1779 : reg648)) ?
                        reg676 : reg1135));
  assign wire1822 = reg1777[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      if (wire3[(3'h6):(3'h6)])
        begin
          if (reg1816[(3'h5):(3'h4)])
            begin
              for (forvar1823 = (1'h0); (forvar1823 < (2'h2)); forvar1823 = (forvar1823 + (1'h1)))
                begin
                  if ((((&(reg733 ? (8'ha9) : reg702)) ?
                      reg1098[(2'h2):(1'h0)] : (^~(reg1166 ?
                          reg1773 : wire631))) <= reg1168[(1'h0):(1'h0)]))
                    begin
                      reg1824 <= (reg1095 ?
                          (reg655 ?
                              ($unsigned(reg1089) && reg685[(1'h0):(1'h0)]) : reg1094[(4'ha):(3'h4)]) : (-(~&(8'h9d))));
                      reg1825 <= ((+(~$signed(reg692))) | reg1768);
                      reg1826 <= reg664;
                      reg1827 <= reg659;
                    end
                  else
                    begin
                      reg1824 <= ($signed({(reg715 ?
                              reg660 : reg641)}) - $unsigned(reg656));
                      reg1825 <= (reg1798 - $signed($unsigned(reg707)));
                    end
                  for (forvar1828 = (1'h0); (forvar1828 < (1'h0)); forvar1828 = (forvar1828 + (1'h1)))
                    begin
                      reg1829 <= $unsigned(reg693);
                      reg1830 <= {$signed((reg1153[(3'h6):(3'h6)] ?
                              $signed(reg693) : (reg692 ? reg650 : reg1774)))};
                      reg1831 <= $unsigned(((8'hb7) ?
                          $unsigned((reg1096 * reg713)) : (|$signed(reg1103))));
                      reg1832 <= (^~reg636[(4'ha):(4'h8)]);
                    end
                  for (forvar1833 = (1'h0); (forvar1833 < (2'h3)); forvar1833 = (forvar1833 + (1'h1)))
                    begin
                      reg1834 <= ($unsigned(forvar1823) == {(~(reg1128 >>> reg1787))});
                      reg1835 <= reg696;
                      reg1836 <= reg663[(3'h4):(3'h4)];
                    end
                  if ($unsigned($signed(reg1113[(2'h2):(2'h2)])))
                    begin
                      reg1837 <= reg693;
                    end
                  else
                    begin
                      reg1837 <= reg1127;
                      reg1838 <= (reg737 ?
                          {($signed(reg1114) ^~ $unsigned(reg638))} : $unsigned(reg1152));
                    end
                end
            end
          else
            begin
              for (forvar1823 = (1'h0); (forvar1823 < (2'h2)); forvar1823 = (forvar1823 + (1'h1)))
                begin
                  reg1824 <= reg662[(1'h1):(1'h0)];
                  if (reg1107[(4'hc):(1'h1)])
                    begin
                      reg1825 <= ($unsigned(reg1160) <= {($unsigned(wire0) ?
                              (8'ha8) : $signed(wire1086))});
                      reg1826 <= $unsigned(((~&reg714[(1'h1):(1'h0)]) ?
                          $signed({reg1111}) : reg1775));
                    end
                  else
                    begin
                      reg1825 <= ((^~$unsigned(reg1780)) ?
                          (reg642[(3'h7):(1'h0)] ?
                              (!(reg1094 ?
                                  (8'ha4) : reg1130)) : ($unsigned(reg1123) >= reg1151[(1'h0):(1'h0)])) : (~($signed(reg721) ^~ (reg1818 ?
                              reg1805 : reg1136))));
                    end
                end
              for (forvar1827 = (1'h0); (forvar1827 < (2'h3)); forvar1827 = (forvar1827 + (1'h1)))
                begin
                  if ({(&$signed($signed(reg1836)))})
                    begin
                      reg1828 <= wire3[(3'h7):(3'h7)];
                    end
                  else
                    begin
                      reg1828 <= $signed((($signed(reg667) + $signed((8'hab))) >>> $signed($signed((8'ha2)))));
                      reg1829 <= $signed(reg1834);
                      reg1830 <= reg647[(3'h5):(1'h0)];
                      reg1831 <= $signed((8'ha7));
                    end
                  reg1832 <= ((-$signed($signed(reg1759))) != $unsigned((reg711[(3'h4):(2'h2)] > $unsigned(reg1149))));
                  for (forvar1833 = (1'h0); (forvar1833 < (1'h1)); forvar1833 = (forvar1833 + (1'h1)))
                    begin
                      reg1834 <= reg1757;
                    end
                  for (forvar1835 = (1'h0); (forvar1835 < (2'h2)); forvar1835 = (forvar1835 + (1'h1)))
                    begin
                      reg1836 <= ((reg1775 ?
                          ($signed((8'ha5)) && $unsigned(forvar1828)) : ((reg722 >> reg1151) >> (reg1788 ?
                              reg662 : reg1837))) ~^ {$unsigned($unsigned(reg1095))});
                      reg1837 <= ((^($unsigned((8'ha2)) == reg657)) ?
                          (&((wire631 <= reg706) ?
                              (~^reg731) : reg1808[(2'h2):(1'h0)])) : ((~|reg1832[(3'h4):(3'h4)]) ?
                              (8'hb9) : reg1128));
                    end
                end
            end
          for (forvar1839 = (1'h0); (forvar1839 < (1'h1)); forvar1839 = (forvar1839 + (1'h1)))
            begin
              if ($unsigned(reg723[(2'h2):(1'h0)]))
                begin
                  if ((-$unsigned(reg679[(3'h5):(2'h2)])))
                    begin
                      reg1840 <= (reg1776 ?
                          (((reg1781 < (8'had)) ?
                              wire1822[(3'h4):(1'h1)] : reg1110[(3'h5):(2'h2)]) | (+$signed(reg638))) : reg644);
                      reg1841 <= reg1135[(4'he):(3'h4)];
                    end
                  else
                    begin
                      reg1840 <= ($signed($signed($signed(reg1828))) ?
                          reg1096 : reg1161[(3'h5):(1'h1)]);
                      reg1841 <= (8'ha1);
                      reg1842 <= (((+$signed(reg685)) != $unsigned(reg1125[(2'h2):(1'h1)])) ?
                          reg1149 : reg1147[(1'h0):(1'h0)]);
                    end
                  for (forvar1843 = (1'h0); (forvar1843 < (1'h1)); forvar1843 = (forvar1843 + (1'h1)))
                    begin
                      reg1844 <= $signed({($unsigned(reg1170) && {reg719})});
                      reg1845 <= $signed(reg683);
                      reg1846 <= (~&(((reg1771 && wire1) ?
                              (~&reg1794) : $signed(reg1094)) ?
                          wire1[(3'h5):(3'h5)] : (8'had)));
                    end
                  for (forvar1847 = (1'h0); (forvar1847 < (2'h3)); forvar1847 = (forvar1847 + (1'h1)))
                    begin
                      reg1848 <= {(reg695 >>> wire4)};
                      reg1849 <= {($signed(reg642[(2'h3):(1'h0)]) * $signed(reg1167[(3'h6):(3'h5)]))};
                    end
                end
              else
                begin
                  reg1840 <= reg1158[(3'h6):(3'h6)];
                end
              if ($signed($unsigned($unsigned((reg663 <<< reg1144)))))
                begin
                  for (forvar1850 = (1'h0); (forvar1850 < (2'h2)); forvar1850 = (forvar1850 + (1'h1)))
                    begin
                      reg1851 <= ({((reg728 ? reg1824 : reg678) ?
                                  $signed(reg1828) : reg1768)} ?
                          $unsigned($unsigned(reg1117[(1'h0):(1'h0)])) : {reg698});
                      reg1852 <= ($unsigned(reg1127[(4'hb):(1'h1)]) ?
                          {reg1765} : $unsigned((~^{forvar1847})));
                      reg1853 <= (-(|$signed(reg668)));
                    end
                  reg1854 <= reg1770[(4'hb):(4'hb)];
                  for (forvar1855 = (1'h0); (forvar1855 < (1'h1)); forvar1855 = (forvar1855 + (1'h1)))
                    begin
                      reg1856 <= (-(~^$signed($signed(reg1146))));
                    end
                end
              else
                begin
                  for (forvar1850 = (1'h0); (forvar1850 < (1'h0)); forvar1850 = (forvar1850 + (1'h1)))
                    begin
                      reg1851 <= {$unsigned(($signed((8'hb8)) ?
                              ((8'had) ?
                                  reg1835 : reg1781) : $signed(reg728)))};
                    end
                  for (forvar1852 = (1'h0); (forvar1852 < (2'h3)); forvar1852 = (forvar1852 + (1'h1)))
                    begin
                      reg1853 <= $signed((reg699[(2'h3):(1'h0)] ~^ (reg1795[(1'h1):(1'h0)] <<< (reg684 ?
                          reg638 : reg718))));
                      reg1854 <= reg727[(4'hd):(4'hc)];
                      reg1855 <= $signed((reg738 + $signed((8'ha2))));
                      reg1856 <= ($unsigned({reg1777}) ?
                          (((-reg1807) | (8'hb2)) ?
                              reg1793[(4'hf):(4'hd)] : ($signed(reg679) ^ $unsigned(reg726))) : (((|reg1100) ?
                                  reg715[(3'h4):(1'h0)] : reg688[(1'h1):(1'h1)]) ?
                              {((8'haf) ?
                                      reg694 : (8'hb0))} : forvar1823[(1'h0):(1'h0)]));
                    end
                  if (reg706)
                    begin
                      reg1857 <= (~|(reg666 ?
                          reg1807[(1'h1):(1'h1)] : $unsigned(((8'hb8) ?
                              reg726 : reg1830))));
                    end
                  else
                    begin
                      reg1857 <= $unsigned($unsigned($signed(reg1804[(4'h8):(3'h4)])));
                      reg1858 <= (|$unsigned(((~&reg1779) + ((8'h9e) ?
                          reg1110 : reg663))));
                      reg1859 <= $signed((reg1103[(2'h2):(1'h1)] ?
                          (~&((8'hb8) >>> reg1820)) : (+forvar1835[(1'h1):(1'h0)])));
                    end
                  if (reg731[(1'h1):(1'h1)])
                    begin
                      reg1860 <= reg677;
                    end
                  else
                    begin
                      reg1860 <= ((reg661 ?
                          (reg696[(4'ha):(2'h2)] & reg1762[(2'h2):(2'h2)]) : {(reg729 == reg714)}) ~^ $unsigned({((8'ha9) + reg693)}));
                      reg1861 <= ((((8'ha7) ?
                              (reg643 ?
                                  reg1806 : reg1796) : {(8'h9d)}) << (((8'ha9) ?
                              reg1757 : reg730) ^ {reg1846})) ?
                          {($unsigned(reg709) ?
                                  $unsigned(reg674) : $unsigned(reg1799))} : $unsigned($unsigned(reg1805[(2'h3):(1'h0)])));
                      reg1862 <= (reg1861 ~^ ($unsigned($signed(reg1788)) - ({reg687} ?
                          (reg1819 <= reg716) : (reg1143 >>> reg720))));
                      reg1863 <= $signed(reg1844);
                    end
                end
              for (forvar1864 = (1'h0); (forvar1864 < (1'h1)); forvar1864 = (forvar1864 + (1'h1)))
                begin
                  if (reg1127[(3'h4):(2'h3)])
                    begin
                      reg1865 <= $unsigned(reg1758);
                      reg1866 <= $unsigned(($signed({reg1089}) ?
                          reg715 : $signed(reg654[(3'h5):(1'h0)])));
                      reg1867 <= ((((-reg1134) ?
                              reg727[(4'h8):(3'h6)] : $unsigned((8'hb2))) < $unsigned(reg651)) ?
                          $signed(({reg1780} & $signed(reg1826))) : reg1096);
                    end
                  else
                    begin
                      reg1865 <= forvar1864;
                      reg1866 <= $unsigned((wire631 ?
                          $signed((reg638 ?
                              reg1793 : reg1867)) : $signed({(8'hb1)})));
                      reg1867 <= ($unsigned((reg1857 ?
                              (wire632 ? (8'h9d) : reg1816) : reg659)) ?
                          (!($unsigned(reg1126) + $unsigned(reg1865))) : (($unsigned(reg661) ?
                                  ((8'ha9) ?
                                      (8'hb9) : reg1136) : $unsigned(reg1831)) ?
                              {$signed((8'ha3))} : reg1153));
                      reg1868 <= {reg1168[(1'h1):(1'h0)]};
                    end
                  reg1869 <= reg690;
                  for (forvar1870 = (1'h0); (forvar1870 < (1'h1)); forvar1870 = (forvar1870 + (1'h1)))
                    begin
                      reg1871 <= reg1805[(1'h1):(1'h0)];
                      reg1872 <= ({$unsigned((~&reg1109))} ~^ ({$unsigned(forvar1833)} * reg1820[(4'hb):(4'hb)]));
                      reg1873 <= (~&(+$unsigned(((8'h9f) ? reg1785 : reg698))));
                      reg1874 <= (~&(reg1110[(1'h0):(1'h0)] * $unsigned(reg1151[(3'h7):(2'h2)])));
                    end
                  if ($unsigned((~|$signed($unsigned((8'hb2))))))
                    begin
                      reg1875 <= $unsigned($unsigned(reg1841[(3'h5):(2'h2)]));
                      reg1876 <= $unsigned({{(-reg1819)}});
                      reg1877 <= reg719[(2'h3):(2'h3)];
                      reg1878 <= (^$signed($unsigned((~^reg701))));
                    end
                  else
                    begin
                      reg1875 <= (reg1110 ?
                          $signed(reg734) : ((~^$unsigned(reg1829)) >= reg636));
                    end
                end
              reg1879 <= (^reg705[(2'h2):(1'h0)]);
            end
        end
      else
        begin
          reg1823 <= {($signed($unsigned((8'hb1))) ?
                  reg1841 : ((reg1149 ? (8'ha0) : reg733) ?
                      reg1798 : reg1115))};
          for (forvar1824 = (1'h0); (forvar1824 < (2'h3)); forvar1824 = (forvar1824 + (1'h1)))
            begin
              reg1825 <= $unsigned((reg1766[(3'h5):(1'h0)] ?
                  (-reg1793[(3'h5):(3'h5)]) : reg1858[(3'h5):(2'h2)]));
            end
        end
      for (forvar1880 = (1'h0); (forvar1880 < (2'h2)); forvar1880 = (forvar1880 + (1'h1)))
        begin
          for (forvar1881 = (1'h0); (forvar1881 < (1'h0)); forvar1881 = (forvar1881 + (1'h1)))
            begin
              for (forvar1882 = (1'h0); (forvar1882 < (1'h0)); forvar1882 = (forvar1882 + (1'h1)))
                begin
                  for (forvar1883 = (1'h0); (forvar1883 < (2'h2)); forvar1883 = (forvar1883 + (1'h1)))
                    begin
                      reg1884 <= $unsigned(($unsigned((reg694 | reg1131)) ^~ $signed((reg649 ?
                          reg726 : reg738))));
                    end
                  if (reg1760)
                    begin
                      reg1885 <= (reg674[(2'h3):(1'h0)] ?
                          reg1100[(4'h9):(2'h3)] : reg701[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg1885 <= {$unsigned(reg695)};
                      reg1886 <= reg1115[(4'hd):(1'h1)];
                    end
                end
              reg1887 <= {$unsigned(($signed(reg659) <<< $signed(wire1)))};
              for (forvar1888 = (1'h0); (forvar1888 < (1'h1)); forvar1888 = (forvar1888 + (1'h1)))
                begin
                  reg1889 <= (~&{($signed((8'hb8)) + {reg685})});
                  for (forvar1890 = (1'h0); (forvar1890 < (2'h3)); forvar1890 = (forvar1890 + (1'h1)))
                    begin
                      reg1891 <= (~&$unsigned($signed((reg1762 ?
                          reg1838 : reg656))));
                    end
                  for (forvar1892 = (1'h0); (forvar1892 < (2'h3)); forvar1892 = (forvar1892 + (1'h1)))
                    begin
                      reg1893 <= $signed(reg1089);
                    end
                end
            end
          for (forvar1894 = (1'h0); (forvar1894 < (1'h1)); forvar1894 = (forvar1894 + (1'h1)))
            begin
              if ((^reg1865))
                begin
                  if ((($unsigned((reg1119 && reg639)) - reg1108) ?
                      (~&$unsigned($unsigned(reg714))) : (reg1859 ?
                          reg731 : wire1086[(3'h5):(1'h0)])))
                    begin
                      reg1895 <= $signed($signed(reg1886[(3'h6):(2'h3)]));
                      reg1896 <= ({((8'h9e) > forvar1827[(1'h1):(1'h1)])} > reg1134[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg1895 <= (~$unsigned($signed((reg1808 ?
                          reg1830 : reg725))));
                      reg1896 <= ((|wire1822) > (($signed(reg1836) ?
                          (reg709 ^ reg1854) : (reg702 ?
                              reg696 : reg1877)) && reg1104));
                      reg1897 <= $unsigned((^~($unsigned(reg1808) ?
                          (~(8'h9d)) : reg679[(2'h2):(2'h2)])));
                    end
                  reg1898 <= $unsigned(reg1166[(3'h5):(1'h1)]);
                  reg1899 <= reg690[(3'h7):(3'h6)];
                end
              else
                begin
                  if (reg1127[(4'h8):(3'h6)])
                    begin
                      reg1895 <= $signed($unsigned((+forvar1843[(2'h2):(1'h1)])));
                    end
                  else
                    begin
                      reg1895 <= ((forvar1880[(1'h0):(1'h0)] ?
                              {(~|reg1867)} : reg1778[(1'h1):(1'h0)]) ?
                          ((reg1787[(1'h1):(1'h0)] ?
                                  (reg1119 < reg1120) : reg732[(3'h6):(2'h3)]) ?
                              {(!reg684)} : ((reg1838 ?
                                  reg1849 : wire631) < (reg1132 ?
                                  reg1889 : (8'hae)))) : (^~({wire1821} <<< (~(8'ha0)))));
                      reg1896 <= (({$unsigned(wire1)} >= reg1823[(3'h4):(1'h0)]) ?
                          (!$signed((!reg1818))) : reg1132);
                      reg1897 <= ((reg1784 - ((reg1124 ? (8'ha9) : reg1789) ?
                              reg1842 : {(8'hb8)})) ?
                          {(|(~^forvar1864))} : (8'ha6));
                    end
                end
            end
          reg1900 <= $unsigned(reg1873[(1'h0):(1'h0)]);
          reg1901 <= (|reg1101[(3'h4):(2'h2)]);
        end
    end
  assign wire1902 = reg1124;
  assign wire1903 = (~(~^(-(reg1760 ? reg1774 : reg1115))));
  assign wire1904 = ((-reg689) ?
                        $unsigned(reg1153) : {((reg677 << (8'hb0)) ^~ $signed(wire631))});
  assign wire1905 = ((reg1846[(4'h9):(3'h5)] ?
                        (|((8'h9c) | reg1799)) : {reg1122[(1'h0):(1'h0)]}) ^~ $signed(reg1846));
  assign wire1906 = reg737[(1'h0):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1171
#(parameter param1752 = {((-((8'ha9) >>> (8'hb0))) ? (!(~&(8'hb4))) : (((8'h9d) | (8'hac)) < ((8'ha0) | (8'ha5))))})
(y, clk, wire1176, wire1175, wire1174, wire1173, wire1172);
  output wire [(32'h896):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire1176;
  input wire signed [(4'h8):(1'h0)] wire1175;
  input wire [(2'h3):(1'h0)] wire1174;
  input wire signed [(4'hb):(1'h0)] wire1173;
  input wire signed [(4'hf):(1'h0)] wire1172;
  wire [(4'he):(1'h0)] wire1751;
  wire [(4'h8):(1'h0)] wire1683;
  wire [(4'hb):(1'h0)] wire1682;
  wire signed [(4'hf):(1'h0)] wire1681;
  wire signed [(2'h2):(1'h0)] wire1531;
  wire [(4'h9):(1'h0)] wire1178;
  wire signed [(4'hc):(1'h0)] wire1177;
  reg [(4'ha):(1'h0)] reg1750 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1749 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1748 = (1'h0);
  reg [(4'hd):(1'h0)] reg1747 = (1'h0);
  reg [(3'h5):(1'h0)] reg1746 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1745 = (1'h0);
  reg [(2'h3):(1'h0)] reg1744 = (1'h0);
  reg [(4'h8):(1'h0)] reg1743 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1742 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1741 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1739 = (1'h0);
  reg [(4'h8):(1'h0)] reg1734 = (1'h0);
  reg [(3'h4):(1'h0)] reg1738 = (1'h0);
  reg [(3'h6):(1'h0)] reg1737 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1736 = (1'h0);
  reg [(4'hc):(1'h0)] reg1735 = (1'h0);
  reg [(4'hc):(1'h0)] reg1733 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1730 = (1'h0);
  reg [(4'he):(1'h0)] reg1729 = (1'h0);
  reg [(4'ha):(1'h0)] reg1727 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1726 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1725 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1723 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1718 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1712 = (1'h0);
  reg [(4'he):(1'h0)] reg1710 = (1'h0);
  reg [(3'h4):(1'h0)] reg1707 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1699 = (1'h0);
  reg [(3'h4):(1'h0)] reg1698 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1689 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1722 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1721 = (1'h0);
  reg [(3'h7):(1'h0)] reg1720 = (1'h0);
  reg [(2'h2):(1'h0)] reg1719 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1717 = (1'h0);
  reg [(4'h9):(1'h0)] reg1716 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1715 = (1'h0);
  reg [(3'h4):(1'h0)] reg1714 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1713 = (1'h0);
  reg [(4'h8):(1'h0)] reg1711 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1709 = (1'h0);
  reg [(3'h4):(1'h0)] reg1708 = (1'h0);
  reg [(3'h5):(1'h0)] reg1706 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1705 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1704 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1703 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1702 = (1'h0);
  reg [(4'hf):(1'h0)] reg1701 = (1'h0);
  reg [(4'ha):(1'h0)] reg1700 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1697 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1696 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1695 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1694 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1693 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1692 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1691 = (1'h0);
  reg [(5'h10):(1'h0)] reg1690 = (1'h0);
  reg [(4'hf):(1'h0)] reg1688 = (1'h0);
  reg [(4'he):(1'h0)] reg1686 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1684 = (1'h0);
  reg [(4'ha):(1'h0)] reg1673 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1680 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1679 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1678 = (1'h0);
  reg [(2'h3):(1'h0)] reg1677 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1676 = (1'h0);
  reg [(3'h5):(1'h0)] reg1675 = (1'h0);
  reg [(2'h2):(1'h0)] reg1674 = (1'h0);
  reg [(3'h4):(1'h0)] reg1672 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1671 = (1'h0);
  reg [(4'hc):(1'h0)] reg1670 = (1'h0);
  reg [(4'hb):(1'h0)] reg1669 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1668 = (1'h0);
  reg [(4'h9):(1'h0)] reg1667 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1666 = (1'h0);
  reg [(4'ha):(1'h0)] reg1665 = (1'h0);
  reg [(2'h3):(1'h0)] reg1664 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1662 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1661 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1660 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1657 = (1'h0);
  reg [(2'h2):(1'h0)] reg1656 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1652 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1651 = (1'h0);
  reg [(4'h9):(1'h0)] reg1639 = (1'h0);
  reg [(3'h6):(1'h0)] reg1636 = (1'h0);
  reg [(4'hd):(1'h0)] reg1635 = (1'h0);
  reg [(4'h8):(1'h0)] reg1650 = (1'h0);
  reg [(2'h3):(1'h0)] reg1649 = (1'h0);
  reg [(4'h8):(1'h0)] reg1648 = (1'h0);
  reg [(4'he):(1'h0)] reg1647 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1646 = (1'h0);
  reg [(3'h6):(1'h0)] reg1644 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1643 = (1'h0);
  reg [(3'h5):(1'h0)] reg1642 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1641 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1640 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1637 = (1'h0);
  reg [(4'h9):(1'h0)] reg1626 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1634 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1633 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1632 = (1'h0);
  reg [(3'h4):(1'h0)] reg1631 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1630 = (1'h0);
  reg [(4'hd):(1'h0)] reg1629 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1628 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1627 = (1'h0);
  reg [(5'h10):(1'h0)] reg1625 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1623 = (1'h0);
  reg [(4'h8):(1'h0)] reg1622 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1621 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1620 = (1'h0);
  reg [(4'ha):(1'h0)] reg1618 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1617 = (1'h0);
  reg [(3'h5):(1'h0)] reg1615 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1614 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1613 = (1'h0);
  reg [(4'h8):(1'h0)] reg1612 = (1'h0);
  reg [(3'h7):(1'h0)] reg1611 = (1'h0);
  reg [(2'h3):(1'h0)] reg1598 = (1'h0);
  reg [(3'h7):(1'h0)] reg1609 = (1'h0);
  reg [(4'h9):(1'h0)] reg1608 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1607 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1606 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1605 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1603 = (1'h0);
  reg [(3'h4):(1'h0)] reg1602 = (1'h0);
  reg [(4'h9):(1'h0)] reg1601 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1600 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1599 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1597 = (1'h0);
  reg [(4'hd):(1'h0)] reg1596 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1594 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1593 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1592 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1591 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1590 = (1'h0);
  reg [(4'he):(1'h0)] reg1589 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1587 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1584 = (1'h0);
  reg [(4'hf):(1'h0)] reg1583 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1582 = (1'h0);
  reg [(2'h3):(1'h0)] reg1581 = (1'h0);
  reg [(3'h5):(1'h0)] reg1579 = (1'h0);
  reg [(4'he):(1'h0)] reg1578 = (1'h0);
  reg [(5'h10):(1'h0)] reg1577 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1576 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1573 = (1'h0);
  reg [(4'h8):(1'h0)] reg1570 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1569 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1568 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1567 = (1'h0);
  reg [(3'h4):(1'h0)] reg1566 = (1'h0);
  reg [(2'h3):(1'h0)] reg1565 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1564 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1563 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1562 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1561 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1559 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1558 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1557 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1555 = (1'h0);
  reg [(3'h4):(1'h0)] reg1554 = (1'h0);
  reg [(3'h6):(1'h0)] reg1553 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1552 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1549 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1546 = (1'h0);
  reg [(4'ha):(1'h0)] reg1542 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1548 = (1'h0);
  reg [(4'hb):(1'h0)] reg1547 = (1'h0);
  reg [(3'h4):(1'h0)] reg1545 = (1'h0);
  reg [(4'he):(1'h0)] reg1544 = (1'h0);
  reg [(4'ha):(1'h0)] reg1543 = (1'h0);
  reg [(4'ha):(1'h0)] reg1541 = (1'h0);
  reg [(4'hb):(1'h0)] reg1540 = (1'h0);
  reg [(4'h8):(1'h0)] reg1539 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1538 = (1'h0);
  reg [(3'h5):(1'h0)] reg1537 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1740 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1734 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1732 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1731 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1728 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1724 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1721 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1709 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1708 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1702 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1696 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1695 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1694 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1688 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1714 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1718 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1712 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1710 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1707 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1699 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1698 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1689 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1687 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1685 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1673 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1663 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1659 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1658 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1655 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1654 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1653 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1650 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1642 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1631 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1647 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1645 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1639 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1638 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1636 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1635 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1625 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1626 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1624 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1619 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1616 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1610 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1604 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1598 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1595 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1588 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1586 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1585 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1580 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1575 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1574 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1572 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1571 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1560 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1556 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1551 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1550 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1546 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1542 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1536 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1535 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1534 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1533 = (1'h0);
  assign y = {wire1751,
                 wire1683,
                 wire1682,
                 wire1681,
                 wire1531,
                 wire1178,
                 wire1177,
                 reg1750,
                 reg1749,
                 reg1748,
                 reg1747,
                 reg1746,
                 reg1745,
                 reg1744,
                 reg1743,
                 reg1742,
                 reg1741,
                 reg1739,
                 reg1734,
                 reg1738,
                 reg1737,
                 reg1736,
                 reg1735,
                 reg1733,
                 reg1730,
                 reg1729,
                 reg1727,
                 reg1726,
                 reg1725,
                 reg1723,
                 reg1718,
                 reg1712,
                 reg1710,
                 reg1707,
                 reg1699,
                 reg1698,
                 reg1689,
                 reg1722,
                 reg1721,
                 reg1720,
                 reg1719,
                 reg1717,
                 reg1716,
                 reg1715,
                 reg1714,
                 reg1713,
                 reg1711,
                 reg1709,
                 reg1708,
                 reg1706,
                 reg1705,
                 reg1704,
                 reg1703,
                 reg1702,
                 reg1701,
                 reg1700,
                 reg1697,
                 reg1696,
                 reg1695,
                 reg1694,
                 reg1693,
                 reg1692,
                 reg1691,
                 reg1690,
                 reg1688,
                 reg1686,
                 reg1684,
                 reg1673,
                 reg1680,
                 reg1679,
                 reg1678,
                 reg1677,
                 reg1676,
                 reg1675,
                 reg1674,
                 reg1672,
                 reg1671,
                 reg1670,
                 reg1669,
                 reg1668,
                 reg1667,
                 reg1666,
                 reg1665,
                 reg1664,
                 reg1662,
                 reg1661,
                 reg1660,
                 reg1657,
                 reg1656,
                 reg1652,
                 reg1651,
                 reg1639,
                 reg1636,
                 reg1635,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1647,
                 reg1646,
                 reg1644,
                 reg1643,
                 reg1642,
                 reg1641,
                 reg1640,
                 reg1637,
                 reg1626,
                 reg1634,
                 reg1633,
                 reg1632,
                 reg1631,
                 reg1630,
                 reg1629,
                 reg1628,
                 reg1627,
                 reg1625,
                 reg1623,
                 reg1622,
                 reg1621,
                 reg1620,
                 reg1618,
                 reg1617,
                 reg1615,
                 reg1614,
                 reg1613,
                 reg1612,
                 reg1611,
                 reg1598,
                 reg1609,
                 reg1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1603,
                 reg1602,
                 reg1601,
                 reg1600,
                 reg1599,
                 reg1597,
                 reg1596,
                 reg1594,
                 reg1593,
                 reg1592,
                 reg1591,
                 reg1590,
                 reg1589,
                 reg1587,
                 reg1584,
                 reg1583,
                 reg1582,
                 reg1581,
                 reg1579,
                 reg1578,
                 reg1577,
                 reg1576,
                 reg1573,
                 reg1570,
                 reg1569,
                 reg1568,
                 reg1567,
                 reg1566,
                 reg1565,
                 reg1564,
                 reg1563,
                 reg1562,
                 reg1561,
                 reg1559,
                 reg1558,
                 reg1557,
                 reg1555,
                 reg1554,
                 reg1553,
                 reg1552,
                 reg1549,
                 reg1546,
                 reg1542,
                 reg1548,
                 reg1547,
                 reg1545,
                 reg1544,
                 reg1543,
                 reg1541,
                 reg1540,
                 reg1539,
                 reg1538,
                 reg1537,
                 forvar1740,
                 forvar1734,
                 forvar1732,
                 forvar1731,
                 forvar1728,
                 forvar1724,
                 forvar1721,
                 forvar1709,
                 forvar1708,
                 forvar1702,
                 forvar1696,
                 forvar1695,
                 forvar1694,
                 forvar1688,
                 forvar1714,
                 forvar1718,
                 forvar1712,
                 forvar1710,
                 forvar1707,
                 forvar1699,
                 forvar1698,
                 forvar1689,
                 forvar1687,
                 forvar1685,
                 forvar1673,
                 forvar1663,
                 forvar1659,
                 forvar1658,
                 forvar1655,
                 forvar1654,
                 forvar1653,
                 forvar1650,
                 forvar1642,
                 forvar1631,
                 forvar1647,
                 forvar1645,
                 forvar1639,
                 forvar1638,
                 forvar1636,
                 forvar1635,
                 forvar1625,
                 forvar1626,
                 forvar1624,
                 forvar1619,
                 forvar1616,
                 forvar1610,
                 forvar1604,
                 forvar1598,
                 forvar1595,
                 forvar1588,
                 forvar1586,
                 forvar1585,
                 forvar1580,
                 forvar1575,
                 forvar1574,
                 forvar1572,
                 forvar1571,
                 forvar1560,
                 forvar1556,
                 forvar1551,
                 forvar1550,
                 forvar1546,
                 forvar1542,
                 forvar1536,
                 forvar1535,
                 forvar1534,
                 forvar1533,
                 (1'h0)};
  assign wire1177 = (^~wire1176[(3'h6):(3'h5)]);
  assign wire1178 = wire1177;
  module1179 #() modinst1532 (.wire1182(wire1177), .wire1181(wire1173), .y(wire1531), .wire1180(wire1175), .clk(clk), .wire1183(wire1172));
  always
    @(posedge clk) begin
      for (forvar1533 = (1'h0); (forvar1533 < (1'h1)); forvar1533 = (forvar1533 + (1'h1)))
        begin
          for (forvar1534 = (1'h0); (forvar1534 < (1'h1)); forvar1534 = (forvar1534 + (1'h1)))
            begin
              for (forvar1535 = (1'h0); (forvar1535 < (1'h1)); forvar1535 = (forvar1535 + (1'h1)))
                begin
                  for (forvar1536 = (1'h0); (forvar1536 < (2'h3)); forvar1536 = (forvar1536 + (1'h1)))
                    begin
                      reg1537 <= ((^~$signed(forvar1534[(4'h9):(3'h6)])) * ($signed(wire1531) ?
                          ($unsigned(forvar1534) ^ $unsigned((8'ha5))) : wire1178[(1'h1):(1'h0)]));
                      reg1538 <= (((&(&reg1537)) ?
                          (wire1176 <= (forvar1533 ^ wire1173)) : ((forvar1534 ~^ forvar1534) ?
                              (!wire1178) : $unsigned(wire1177))) < $unsigned(($unsigned((8'ha8)) ?
                          wire1178 : $unsigned(wire1174))));
                      reg1539 <= forvar1535;
                      reg1540 <= $unsigned($signed((forvar1533[(3'h6):(1'h1)] * reg1538[(1'h1):(1'h1)])));
                    end
                end
              reg1541 <= reg1539;
              if (((!$unsigned((~&wire1175))) > wire1177[(3'h4):(1'h0)]))
                begin
                  for (forvar1542 = (1'h0); (forvar1542 < (1'h1)); forvar1542 = (forvar1542 + (1'h1)))
                    begin
                      reg1543 <= wire1176;
                      reg1544 <= wire1531;
                      reg1545 <= $unsigned($unsigned((|forvar1534[(4'hc):(4'ha)])));
                    end
                  for (forvar1546 = (1'h0); (forvar1546 < (2'h2)); forvar1546 = (forvar1546 + (1'h1)))
                    begin
                      reg1547 <= (((reg1538[(3'h4):(1'h1)] ?
                          reg1539[(3'h4):(1'h1)] : ((8'ha8) < wire1176)) & $unsigned($unsigned(reg1540))) >> $signed((^(forvar1534 ?
                          wire1177 : reg1540))));
                      reg1548 <= ($unsigned(reg1547[(3'h5):(1'h1)]) != $unsigned(wire1173));
                    end
                end
              else
                begin
                  reg1542 <= forvar1535[(3'h5):(2'h2)];
                  reg1543 <= $unsigned({{reg1543}});
                  if (($signed((8'had)) - reg1540))
                    begin
                      reg1544 <= $signed(wire1174[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1544 <= forvar1535;
                      reg1545 <= (((&(+wire1172)) >> $unsigned(((8'hb9) <= reg1540))) ?
                          $unsigned((8'had)) : (((reg1547 * (8'hb6)) || (forvar1533 ?
                                  (8'hb4) : wire1175)) ?
                              (&$unsigned(wire1173)) : {(wire1531 ?
                                      (8'ha8) : reg1545)}));
                      reg1546 <= (~&reg1540[(3'h7):(3'h5)]);
                    end
                end
            end
          if ($unsigned((8'ha7)))
            begin
              reg1549 <= (~^$signed(reg1542[(2'h2):(1'h0)]));
              for (forvar1550 = (1'h0); (forvar1550 < (2'h2)); forvar1550 = (forvar1550 + (1'h1)))
                begin
                  for (forvar1551 = (1'h0); (forvar1551 < (1'h1)); forvar1551 = (forvar1551 + (1'h1)))
                    begin
                      reg1552 <= (|forvar1551);
                      reg1553 <= ((((forvar1542 >> forvar1535) | (^~(8'h9d))) >> forvar1551[(4'hd):(3'h4)]) > $signed(($signed(reg1552) + (&(8'h9c)))));
                      reg1554 <= forvar1551[(4'hd):(1'h0)];
                    end
                  reg1555 <= (reg1553 * wire1178[(2'h2):(2'h2)]);
                  for (forvar1556 = (1'h0); (forvar1556 < (1'h1)); forvar1556 = (forvar1556 + (1'h1)))
                    begin
                      reg1557 <= $signed((~&{$signed(reg1554)}));
                      reg1558 <= wire1174[(2'h3):(1'h0)];
                      reg1559 <= $signed((~reg1547));
                    end
                end
            end
          else
            begin
              reg1549 <= ($unsigned((forvar1536 ?
                      reg1559[(3'h4):(1'h1)] : (reg1554 > wire1173))) ?
                  (+reg1549) : reg1540);
            end
          for (forvar1560 = (1'h0); (forvar1560 < (2'h3)); forvar1560 = (forvar1560 + (1'h1)))
            begin
              if ({(((&(8'hb5)) | $unsigned(forvar1534)) ?
                      ((wire1176 | reg1552) ?
                          reg1541[(2'h2):(2'h2)] : (-reg1555)) : reg1552[(3'h5):(1'h1)])})
                begin
                  if ($unsigned(({$unsigned((8'hab))} <<< {{reg1558}})))
                    begin
                      reg1561 <= wire1175[(4'h8):(4'h8)];
                    end
                  else
                    begin
                      reg1561 <= $unsigned((($signed((8'hb1)) + reg1554[(2'h3):(1'h1)]) ?
                          $unsigned((forvar1551 ?
                              forvar1546 : reg1553)) : ($signed(reg1549) ?
                              $unsigned(reg1541) : (~(8'ha9)))));
                      reg1562 <= (-(^~wire1173));
                      reg1563 <= ((($signed(forvar1536) ?
                              (!(8'hb6)) : (reg1537 ? reg1538 : reg1541)) ?
                          reg1559 : reg1559) == ((reg1562 > $signed(reg1537)) == reg1547));
                    end
                  if ($unsigned(reg1538[(3'h5):(1'h0)]))
                    begin
                      reg1564 <= {(8'h9f)};
                      reg1565 <= reg1543[(3'h5):(1'h1)];
                      reg1566 <= $unsigned({{reg1544[(4'h8):(2'h3)]}});
                    end
                  else
                    begin
                      reg1564 <= $signed({forvar1533[(4'hd):(3'h4)]});
                    end
                  if ({$signed(($unsigned(wire1176) & (reg1546 == reg1539)))})
                    begin
                      reg1567 <= (~$unsigned($unsigned({reg1554})));
                      reg1568 <= $signed($signed(reg1546));
                      reg1569 <= $signed((((reg1563 ? reg1541 : (8'ha9)) ?
                          $unsigned(reg1568) : (8'ha6)) - ($unsigned((8'hb8)) >> $signed(reg1553))));
                      reg1570 <= ($unsigned($unsigned((wire1172 + forvar1556))) ?
                          {reg1543} : {wire1173[(4'h9):(3'h5)]});
                    end
                  else
                    begin
                      reg1567 <= ($unsigned((^~(reg1570 == forvar1546))) >> reg1539[(4'h8):(2'h2)]);
                      reg1568 <= ((8'hb5) | ((reg1570 == $signed(forvar1533)) + {$unsigned((8'hba))}));
                    end
                end
              else
                begin
                  if ({forvar1542[(2'h2):(1'h1)]})
                    begin
                      reg1561 <= ((~^$signed($unsigned(reg1552))) << $unsigned((!$unsigned(wire1177))));
                    end
                  else
                    begin
                      reg1561 <= (^~{(~^(reg1537 ? reg1555 : wire1172))});
                      reg1562 <= (^~((forvar1551 ?
                          $signed(forvar1536) : $signed(reg1537)) * forvar1536[(2'h3):(2'h3)]));
                    end
                end
              for (forvar1571 = (1'h0); (forvar1571 < (1'h0)); forvar1571 = (forvar1571 + (1'h1)))
                begin
                  for (forvar1572 = (1'h0); (forvar1572 < (1'h1)); forvar1572 = (forvar1572 + (1'h1)))
                    begin
                      reg1573 <= $unsigned($unsigned(($unsigned((8'hba)) ^ reg1546)));
                    end
                end
              for (forvar1574 = (1'h0); (forvar1574 < (1'h0)); forvar1574 = (forvar1574 + (1'h1)))
                begin
                  for (forvar1575 = (1'h0); (forvar1575 < (2'h2)); forvar1575 = (forvar1575 + (1'h1)))
                    begin
                      reg1576 <= reg1542;
                    end
                  if (reg1539[(3'h7):(2'h2)])
                    begin
                      reg1577 <= reg1555[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg1577 <= (|wire1178[(1'h0):(1'h0)]);
                      reg1578 <= (wire1174 < (~^(~|$unsigned(forvar1536))));
                      reg1579 <= $unsigned((reg1568[(1'h1):(1'h1)] || ($signed(reg1562) <= wire1531)));
                    end
                  for (forvar1580 = (1'h0); (forvar1580 < (2'h2)); forvar1580 = (forvar1580 + (1'h1)))
                    begin
                      reg1581 <= (^~$unsigned($unsigned(forvar1533[(3'h4):(2'h3)])));
                      reg1582 <= $unsigned(((-forvar1534[(3'h7):(3'h6)]) ?
                          ($signed((8'h9d)) >>> (forvar1551 ?
                              reg1561 : (8'ha0))) : $signed((reg1542 ?
                              reg1547 : reg1569))));
                      reg1583 <= (($signed($signed(wire1173)) < ($signed(reg1582) ?
                              (^forvar1580) : $signed(forvar1580))) ?
                          (forvar1533 >= reg1566[(1'h0):(1'h0)]) : ($signed((~&reg1559)) ?
                              {forvar1571} : (~wire1175[(3'h5):(1'h0)])));
                      reg1584 <= (($unsigned($unsigned(forvar1535)) > (+$unsigned(forvar1556))) ?
                          ($unsigned((reg1539 ?
                              (8'ha4) : (8'ha8))) >> $signed($signed((8'ha6)))) : forvar1550[(1'h0):(1'h0)]);
                    end
                end
              for (forvar1585 = (1'h0); (forvar1585 < (1'h1)); forvar1585 = (forvar1585 + (1'h1)))
                begin
                  for (forvar1586 = (1'h0); (forvar1586 < (2'h3)); forvar1586 = (forvar1586 + (1'h1)))
                    begin
                      reg1587 <= (^((reg1577[(4'hd):(2'h2)] ?
                          $signed(wire1531) : ((8'ha2) ?
                              forvar1580 : reg1538)) | reg1543[(2'h2):(2'h2)]));
                    end
                  for (forvar1588 = (1'h0); (forvar1588 < (2'h3)); forvar1588 = (forvar1588 + (1'h1)))
                    begin
                      reg1589 <= (~&forvar1551[(2'h2):(1'h0)]);
                    end
                  reg1590 <= (!(($unsigned(forvar1550) ^ $signed((8'h9d))) ?
                      ((~reg1547) ?
                          (reg1554 ?
                              (8'ha5) : reg1563) : reg1559) : ((forvar1586 <= forvar1560) ?
                          (+wire1174) : $unsigned((8'hb1)))));
                  if ($signed($signed($signed((~forvar1551)))))
                    begin
                      reg1591 <= forvar1550;
                      reg1592 <= (~|(&(|reg1545[(3'h4):(1'h0)])));
                      reg1593 <= (8'had);
                      reg1594 <= (((~|reg1569) && $signed(forvar1585[(2'h2):(1'h1)])) ?
                          (8'h9f) : (reg1563[(3'h6):(3'h5)] - reg1576));
                    end
                  else
                    begin
                      reg1591 <= {$signed(((&forvar1556) ?
                              (~|wire1172) : forvar1574))};
                      reg1592 <= ($signed((+{reg1559})) ?
                          ({$signed((8'hb2))} >>> $unsigned($signed(wire1173))) : $signed($signed(reg1543[(2'h2):(1'h0)])));
                      reg1593 <= (reg1564[(3'h7):(3'h4)] ?
                          $signed(forvar1560) : (+($unsigned(reg1592) == (reg1589 ?
                              forvar1572 : forvar1560))));
                    end
                end
            end
          for (forvar1595 = (1'h0); (forvar1595 < (1'h0)); forvar1595 = (forvar1595 + (1'h1)))
            begin
              reg1596 <= reg1558[(2'h2):(2'h2)];
              reg1597 <= reg1568;
              if ((~^((~&$unsigned(forvar1542)) & reg1579[(2'h2):(1'h0)])))
                begin
                  for (forvar1598 = (1'h0); (forvar1598 < (1'h1)); forvar1598 = (forvar1598 + (1'h1)))
                    begin
                      reg1599 <= (~$signed(reg1577[(3'h7):(3'h6)]));
                      reg1600 <= {($unsigned((~&reg1566)) ?
                              (~|$signed(reg1568)) : forvar1546)};
                      reg1601 <= $signed((forvar1535 >>> ((reg1582 ?
                              reg1596 : reg1576) ?
                          reg1599[(2'h2):(1'h0)] : (!reg1564))));
                      reg1602 <= $signed(reg1579[(1'h1):(1'h1)]);
                    end
                  reg1603 <= (({(forvar1585 ? forvar1551 : reg1554)} ?
                          ((reg1601 ? reg1597 : forvar1588) ~^ (forvar1585 ?
                              forvar1534 : forvar1572)) : ((wire1174 * reg1545) * (forvar1535 ?
                              (8'ha6) : reg1584))) ?
                      $signed({reg1564}) : reg1537[(3'h5):(2'h3)]);
                  for (forvar1604 = (1'h0); (forvar1604 < (1'h1)); forvar1604 = (forvar1604 + (1'h1)))
                    begin
                      reg1605 <= (({(8'hb7)} | (&$signed(reg1578))) || {reg1552[(2'h3):(2'h3)]});
                      reg1606 <= $signed(reg1542[(4'ha):(2'h3)]);
                      reg1607 <= reg1558[(2'h2):(2'h2)];
                      reg1608 <= reg1584;
                    end
                  reg1609 <= reg1567;
                end
              else
                begin
                  reg1598 <= ($signed((reg1579[(3'h4):(2'h2)] + wire1176)) >> {((~reg1542) ?
                          $signed(reg1566) : $signed((8'ha8)))});
                end
              for (forvar1610 = (1'h0); (forvar1610 < (1'h0)); forvar1610 = (forvar1610 + (1'h1)))
                begin
                  if ($signed($unsigned($signed(forvar1571[(1'h0):(1'h0)]))))
                    begin
                      reg1611 <= $signed({(8'hb9)});
                      reg1612 <= reg1603;
                      reg1613 <= $unsigned($unsigned(reg1557[(1'h1):(1'h0)]));
                      reg1614 <= reg1598[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg1611 <= (~&(reg1591 != $signed(reg1568)));
                      reg1612 <= (!(((reg1601 >> (8'haa)) * (reg1582 >> reg1541)) ?
                          $signed(forvar1534) : $unsigned((~^wire1175))));
                      reg1613 <= (((~|reg1591[(4'h8):(1'h0)]) ?
                          reg1549 : {(reg1590 != reg1547)}) ~^ (((reg1579 ?
                              reg1548 : reg1565) ?
                          reg1583 : $unsigned(reg1554)) + reg1577[(4'hd):(4'h9)]));
                      reg1614 <= $signed({(|reg1547[(4'h8):(3'h5)])});
                    end
                  reg1615 <= {(~&$unsigned(reg1592[(1'h0):(1'h0)]))};
                  for (forvar1616 = (1'h0); (forvar1616 < (1'h1)); forvar1616 = (forvar1616 + (1'h1)))
                    begin
                      reg1617 <= forvar1551;
                      reg1618 <= ((reg1577 | {$unsigned(reg1606)}) <= $unsigned($signed($unsigned((8'hb5)))));
                    end
                  for (forvar1619 = (1'h0); (forvar1619 < (2'h2)); forvar1619 = (forvar1619 + (1'h1)))
                    begin
                      reg1620 <= (forvar1616[(3'h7):(2'h2)] >> (reg1568[(1'h1):(1'h1)] ?
                          $unsigned($signed(forvar1572)) : (reg1576 ?
                              (~&(8'hb6)) : reg1596[(4'hb):(3'h6)])));
                      reg1621 <= reg1596;
                      reg1622 <= forvar1535;
                      reg1623 <= (+((reg1582 ?
                          $signed((8'hae)) : (~^(8'hb9))) << reg1622[(3'h4):(3'h4)]));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ({(($signed(reg1564) ? $signed(reg1622) : (^~reg1599)) ?
              ((~^(8'ha4)) ?
                  (reg1602 ? reg1558 : reg1605) : reg1542) : $signed((8'hb1)))})
        begin
          for (forvar1624 = (1'h0); (forvar1624 < (2'h2)); forvar1624 = (forvar1624 + (1'h1)))
            begin
              if ({reg1552[(4'hc):(2'h3)]})
                begin
                  reg1625 <= (($unsigned(reg1590) ?
                      ((reg1592 > (8'h9e)) ~^ (reg1564 ?
                          reg1577 : (8'ha1))) : (~|$signed(reg1583))) * (reg1578[(1'h1):(1'h0)] ?
                      reg1612 : $unsigned({reg1539})));
                  for (forvar1626 = (1'h0); (forvar1626 < (2'h2)); forvar1626 = (forvar1626 + (1'h1)))
                    begin
                      reg1627 <= (^~(^((reg1564 ?
                          forvar1626 : (8'hab)) ~^ (reg1559 ?
                          reg1620 : (8'h9d)))));
                      reg1628 <= reg1594[(3'h4):(1'h0)];
                      reg1629 <= (($unsigned((^~(8'hb1))) ?
                              (|(reg1591 ?
                                  reg1547 : reg1592)) : $unsigned((reg1567 == reg1546))) ?
                          ($signed((wire1531 > wire1172)) < (-$unsigned(reg1579))) : $signed($signed($unsigned(reg1622))));
                      reg1630 <= ($signed((^$unsigned((8'ha6)))) || (reg1602[(1'h0):(1'h0)] ?
                          $unsigned((reg1566 == reg1565)) : $unsigned($signed(reg1583))));
                    end
                  if ($signed(forvar1626))
                    begin
                      reg1631 <= wire1174[(1'h0):(1'h0)];
                      reg1632 <= $signed($signed(((~reg1597) <= $unsigned(reg1579))));
                      reg1633 <= (((^~(^~(8'hb8))) <<< $signed((reg1566 ?
                          reg1559 : (8'hba)))) && $signed({((8'hb1) == reg1541)}));
                    end
                  else
                    begin
                      reg1631 <= {((~$unsigned(reg1623)) ?
                              ((reg1632 < reg1620) + $signed(reg1587)) : (((8'h9e) ?
                                  reg1573 : reg1563) <<< (wire1177 ?
                                  reg1594 : reg1573)))};
                      reg1632 <= ((!{reg1553[(1'h0):(1'h0)]}) ?
                          reg1570 : (((reg1592 << reg1538) ?
                              wire1177[(4'hc):(4'hb)] : {reg1632}) | (reg1559 << (reg1615 * wire1177))));
                      reg1633 <= ((((reg1582 ? reg1557 : reg1537) ?
                          $signed((8'ha2)) : (&reg1600)) + (reg1622[(3'h5):(1'h1)] <= $signed(reg1564))) && reg1609[(3'h4):(1'h0)]);
                    end
                  reg1634 <= (($unsigned((~|forvar1626)) ?
                      $signed((reg1618 ?
                          (8'hb2) : reg1590)) : $unsigned({reg1627})) ~^ $unsigned($signed(reg1594)));
                end
              else
                begin
                  for (forvar1625 = (1'h0); (forvar1625 < (1'h1)); forvar1625 = (forvar1625 + (1'h1)))
                    begin
                      reg1626 <= {reg1544};
                      reg1627 <= ((wire1176 ?
                              ($unsigned(reg1621) && $signed(reg1570)) : $unsigned(reg1541)) ?
                          reg1540 : $signed($signed(reg1568)));
                      reg1628 <= $unsigned((|reg1593));
                      reg1629 <= ((wire1172 ?
                          wire1176 : reg1564) >>> (reg1630 * reg1593));
                    end
                end
            end
          for (forvar1635 = (1'h0); (forvar1635 < (2'h3)); forvar1635 = (forvar1635 + (1'h1)))
            begin
              for (forvar1636 = (1'h0); (forvar1636 < (1'h0)); forvar1636 = (forvar1636 + (1'h1)))
                begin
                  reg1637 <= (8'haa);
                end
              for (forvar1638 = (1'h0); (forvar1638 < (1'h1)); forvar1638 = (forvar1638 + (1'h1)))
                begin
                  for (forvar1639 = (1'h0); (forvar1639 < (2'h2)); forvar1639 = (forvar1639 + (1'h1)))
                    begin
                      reg1640 <= {((!$signed(reg1546)) ?
                              $unsigned($unsigned(reg1543)) : $signed(reg1631[(2'h2):(1'h0)]))};
                      reg1641 <= reg1612[(2'h2):(1'h0)];
                      reg1642 <= $signed(((~&(reg1542 ?
                          (8'ha9) : (8'hb4))) <<< $unsigned((~reg1561))));
                      reg1643 <= $signed((((reg1590 ?
                              reg1539 : reg1600) >> (wire1178 & wire1173)) ?
                          ((reg1630 ? reg1590 : reg1633) ?
                              $signed((8'had)) : {reg1577}) : reg1558));
                    end
                end
              if ($unsigned($unsigned(((reg1611 & forvar1638) != reg1558[(2'h3):(1'h1)]))))
                begin
                  reg1644 <= $unsigned(reg1600[(1'h1):(1'h1)]);
                  for (forvar1645 = (1'h0); (forvar1645 < (2'h2)); forvar1645 = (forvar1645 + (1'h1)))
                    begin
                      reg1646 <= reg1537;
                      reg1647 <= ((reg1538[(1'h0):(1'h0)] ?
                              $unsigned(reg1553[(3'h4):(1'h0)]) : reg1613[(4'hd):(4'hc)]) ?
                          reg1599 : ($signed($signed(reg1570)) > reg1559[(3'h5):(1'h1)]));
                      reg1648 <= ($unsigned(($unsigned(wire1531) + reg1642[(3'h4):(1'h0)])) ?
                          $unsigned(reg1623[(1'h0):(1'h0)]) : (^$unsigned($unsigned(reg1617))));
                      reg1649 <= $unsigned(((~^reg1641[(3'h7):(3'h5)]) ^~ ($unsigned(forvar1635) && wire1175)));
                    end
                end
              else
                begin
                  reg1644 <= {$unsigned(reg1563)};
                  for (forvar1645 = (1'h0); (forvar1645 < (1'h1)); forvar1645 = (forvar1645 + (1'h1)))
                    begin
                      reg1646 <= $signed(reg1631);
                    end
                  for (forvar1647 = (1'h0); (forvar1647 < (1'h1)); forvar1647 = (forvar1647 + (1'h1)))
                    begin
                      reg1648 <= $unsigned(((~|(reg1557 ?
                          reg1547 : (8'h9d))) > {(forvar1636 != forvar1636)}));
                      reg1649 <= {$unsigned($unsigned(reg1569))};
                      reg1650 <= reg1549;
                    end
                end
            end
        end
      else
        begin
          for (forvar1624 = (1'h0); (forvar1624 < (1'h1)); forvar1624 = (forvar1624 + (1'h1)))
            begin
              for (forvar1625 = (1'h0); (forvar1625 < (2'h3)); forvar1625 = (forvar1625 + (1'h1)))
                begin
                  for (forvar1626 = (1'h0); (forvar1626 < (1'h0)); forvar1626 = (forvar1626 + (1'h1)))
                    begin
                      reg1627 <= reg1555[(1'h1):(1'h0)];
                      reg1628 <= $unsigned(((reg1554[(3'h4):(2'h2)] ?
                          (reg1622 ?
                              (8'ha3) : forvar1625) : $unsigned((8'ha6))) != forvar1638[(2'h2):(1'h0)]));
                      reg1629 <= reg1630[(2'h2):(2'h2)];
                    end
                  reg1630 <= ((~{(reg1612 ? reg1642 : reg1582)}) ?
                      reg1644 : (8'hb3));
                  for (forvar1631 = (1'h0); (forvar1631 < (1'h0)); forvar1631 = (forvar1631 + (1'h1)))
                    begin
                      reg1632 <= wire1177[(1'h0):(1'h0)];
                      reg1633 <= (8'ha9);
                      reg1634 <= {$signed({(reg1547 ~^ reg1562)})};
                      reg1635 <= (^(8'had));
                    end
                  if ($signed($unsigned(reg1578[(4'hb):(4'hb)])))
                    begin
                      reg1636 <= $unsigned((+reg1577[(4'hd):(4'h9)]));
                    end
                  else
                    begin
                      reg1636 <= {$unsigned((~(reg1630 ? reg1593 : (8'haf))))};
                      reg1637 <= (~^reg1540);
                    end
                end
            end
          for (forvar1638 = (1'h0); (forvar1638 < (2'h2)); forvar1638 = (forvar1638 + (1'h1)))
            begin
              if ((!({(reg1636 ? reg1581 : (8'hb6))} || ((8'ha0) ?
                  {forvar1647} : $signed(forvar1639)))))
                begin
                  for (forvar1639 = (1'h0); (forvar1639 < (2'h2)); forvar1639 = (forvar1639 + (1'h1)))
                    begin
                      reg1640 <= (^$signed(reg1632));
                      reg1641 <= reg1543;
                    end
                end
              else
                begin
                  if (((-reg1567[(1'h1):(1'h1)]) == (($unsigned(reg1602) | {forvar1636}) ~^ $signed((reg1566 + (8'hb8))))))
                    begin
                      reg1639 <= $unsigned((((reg1540 && reg1596) >> (reg1590 ?
                          reg1549 : forvar1639)) & reg1545[(2'h3):(2'h2)]));
                      reg1640 <= (($unsigned(reg1576[(1'h1):(1'h1)]) ?
                              ($signed(reg1631) <<< (reg1609 ?
                                  reg1565 : (8'ha4))) : {$unsigned(reg1555)}) ?
                          $unsigned(((reg1603 >> reg1631) ?
                              reg1573[(4'h8):(3'h6)] : (wire1176 ?
                                  (8'hb6) : wire1176))) : $unsigned({(reg1633 ?
                                  reg1554 : reg1593)}));
                      reg1641 <= (8'ha0);
                    end
                  else
                    begin
                      reg1639 <= ((reg1639 ? $signed(reg1622) : reg1540) ?
                          (reg1557[(2'h2):(2'h2)] ?
                              reg1648 : ($signed(reg1596) ?
                                  $unsigned(reg1568) : $signed(reg1543))) : $signed(($signed(wire1173) != (~|wire1178))));
                      reg1640 <= ({$signed($signed((8'hb1)))} ?
                          reg1614[(4'h8):(3'h4)] : reg1579);
                    end
                  for (forvar1642 = (1'h0); (forvar1642 < (2'h2)); forvar1642 = (forvar1642 + (1'h1)))
                    begin
                      reg1643 <= ((reg1642 * ($unsigned(reg1578) ?
                          reg1634 : $unsigned(reg1546))) * reg1539);
                      reg1644 <= reg1629;
                    end
                  for (forvar1645 = (1'h0); (forvar1645 < (1'h1)); forvar1645 = (forvar1645 + (1'h1)))
                    begin
                      reg1646 <= $signed({$signed((^reg1573))});
                      reg1647 <= (8'hb9);
                      reg1648 <= (!$unsigned($unsigned({reg1537})));
                      reg1649 <= reg1635[(4'h8):(1'h1)];
                    end
                  for (forvar1650 = (1'h0); (forvar1650 < (1'h0)); forvar1650 = (forvar1650 + (1'h1)))
                    begin
                      reg1651 <= $signed((wire1177[(2'h3):(1'h1)] ?
                          $signed($signed(reg1576)) : (~$signed(reg1553))));
                      reg1652 <= $unsigned((|$signed((reg1611 ?
                          reg1564 : reg1573))));
                    end
                end
            end
          for (forvar1653 = (1'h0); (forvar1653 < (1'h0)); forvar1653 = (forvar1653 + (1'h1)))
            begin
              for (forvar1654 = (1'h0); (forvar1654 < (2'h2)); forvar1654 = (forvar1654 + (1'h1)))
                begin
                  for (forvar1655 = (1'h0); (forvar1655 < (1'h0)); forvar1655 = (forvar1655 + (1'h1)))
                    begin
                      reg1656 <= ($signed((reg1603[(3'h4):(1'h1)] ?
                          (reg1552 | reg1649) : $unsigned((8'h9c)))) > (reg1617[(3'h4):(2'h3)] >>> $signed($unsigned(forvar1639))));
                      reg1657 <= {$unsigned({$signed(forvar1650)})};
                    end
                end
              for (forvar1658 = (1'h0); (forvar1658 < (2'h3)); forvar1658 = (forvar1658 + (1'h1)))
                begin
                  for (forvar1659 = (1'h0); (forvar1659 < (1'h1)); forvar1659 = (forvar1659 + (1'h1)))
                    begin
                      reg1660 <= reg1632;
                      reg1661 <= $unsigned(($signed($signed(forvar1625)) ~^ $signed((|reg1597))));
                      reg1662 <= $signed((-($signed(reg1601) ?
                          {reg1632} : forvar1635)));
                    end
                  for (forvar1663 = (1'h0); (forvar1663 < (2'h2)); forvar1663 = (forvar1663 + (1'h1)))
                    begin
                      reg1664 <= {reg1644[(3'h4):(1'h0)]};
                      reg1665 <= reg1558[(2'h2):(2'h2)];
                    end
                  if ($unsigned((~$unsigned(reg1540[(1'h1):(1'h1)]))))
                    begin
                      reg1666 <= {$unsigned(reg1632[(1'h1):(1'h1)])};
                      reg1667 <= (8'had);
                    end
                  else
                    begin
                      reg1666 <= reg1598;
                      reg1667 <= (~^(+(^~forvar1647[(3'h6):(3'h6)])));
                      reg1668 <= (&$signed({reg1568[(2'h3):(1'h1)]}));
                    end
                  if ({reg1646[(3'h6):(2'h3)]})
                    begin
                      reg1669 <= $unsigned(((((8'ha0) ?
                          reg1623 : reg1613) < reg1629) == reg1564));
                      reg1670 <= (wire1531[(1'h1):(1'h0)] ?
                          $signed((^~$unsigned((8'ha5)))) : reg1643);
                    end
                  else
                    begin
                      reg1669 <= ((reg1568[(2'h3):(2'h2)] ?
                              ((&wire1173) > $signed(reg1649)) : reg1593) ?
                          reg1568[(3'h4):(2'h3)] : $unsigned(wire1174));
                      reg1670 <= reg1569[(3'h7):(1'h1)];
                      reg1671 <= (~$signed((reg1561 >>> (!reg1559))));
                    end
                end
              if (reg1577)
                begin
                  reg1672 <= $signed(forvar1655);
                  for (forvar1673 = (1'h0); (forvar1673 < (1'h1)); forvar1673 = (forvar1673 + (1'h1)))
                    begin
                      reg1674 <= {$signed($unsigned((reg1553 ?
                              reg1665 : forvar1639)))};
                    end
                  if (reg1614[(3'h6):(1'h1)])
                    begin
                      reg1675 <= ({$signed(reg1545[(3'h4):(2'h3)])} * (~&(|reg1621[(3'h6):(1'h0)])));
                      reg1676 <= reg1594;
                      reg1677 <= (~^({$unsigned((8'hb7))} ?
                          ($unsigned((8'hb5)) ^ (~^reg1676)) : reg1584));
                      reg1678 <= reg1607[(4'h8):(4'h8)];
                    end
                  else
                    begin
                      reg1675 <= ((reg1557[(1'h0):(1'h0)] + ((reg1593 < forvar1658) ?
                              (forvar1635 ?
                                  reg1581 : forvar1624) : (reg1598 < reg1627))) ?
                          {(~&reg1657)} : $signed((|{reg1646})));
                      reg1676 <= $signed($signed($unsigned($signed((8'hb7)))));
                      reg1677 <= (8'hae);
                      reg1678 <= ((+wire1177[(4'hc):(4'hc)]) ?
                          reg1603[(4'h8):(3'h7)] : $unsigned(wire1176[(1'h0):(1'h0)]));
                    end
                  if ($unsigned(($unsigned($unsigned(reg1656)) && wire1176)))
                    begin
                      reg1679 <= ((~&{(reg1576 ? reg1555 : reg1627)}) ?
                          $signed(((!reg1660) ?
                              {reg1579} : ((8'hb0) == reg1617))) : reg1546[(1'h1):(1'h0)]);
                      reg1680 <= ((reg1613 ?
                              {$unsigned(reg1593)} : (reg1541 ?
                                  (~|reg1626) : $signed(reg1562))) ?
                          reg1636 : (~&(8'hb2)));
                    end
                  else
                    begin
                      reg1679 <= (({(reg1680 || (8'ha6))} << reg1593[(2'h3):(1'h0)]) && (!$signed({reg1674})));
                      reg1680 <= (^{$signed(reg1643)});
                    end
                end
              else
                begin
                  if ($signed(reg1635[(4'h9):(4'h8)]))
                    begin
                      reg1672 <= reg1540;
                    end
                  else
                    begin
                      reg1672 <= ($unsigned((~|forvar1673[(1'h1):(1'h0)])) - {reg1557[(3'h4):(3'h4)]});
                      reg1673 <= (({reg1671[(1'h0):(1'h0)]} >> $signed($signed(reg1552))) << $signed((+(reg1591 ?
                          reg1633 : reg1596))));
                      reg1674 <= reg1545[(1'h0):(1'h0)];
                    end
                  if (((~&($unsigned(reg1668) ~^ ((8'ha1) ^~ (8'hb8)))) ?
                      (~&(8'hac)) : (-reg1621[(3'h6):(1'h1)])))
                    begin
                      reg1675 <= reg1633;
                      reg1676 <= (({{reg1634}} == $signed($unsigned((8'hb6)))) ?
                          (~^reg1542) : reg1615);
                      reg1677 <= {($signed((+reg1620)) ? reg1544 : (8'hb2))};
                    end
                  else
                    begin
                      reg1675 <= forvar1635[(2'h2):(1'h0)];
                      reg1676 <= {(~(((8'ha0) ? reg1680 : reg1593) ?
                              $unsigned(reg1618) : (|wire1173)))};
                      reg1677 <= wire1176;
                      reg1678 <= reg1637;
                    end
                  if (reg1602)
                    begin
                      reg1679 <= reg1680[(4'hb):(2'h2)];
                      reg1680 <= (((forvar1635[(1'h1):(1'h0)] <= {wire1176}) & $signed((reg1630 ?
                              reg1565 : reg1561))) ?
                          $signed(forvar1653[(3'h4):(1'h1)]) : (reg1597[(3'h6):(3'h4)] ^ $unsigned($signed((8'ha6)))));
                    end
                  else
                    begin
                      reg1679 <= (+{forvar1663[(1'h0):(1'h0)]});
                      reg1680 <= $unsigned($unsigned(reg1563[(3'h4):(1'h1)]));
                    end
                end
            end
        end
    end
  assign wire1681 = reg1647[(4'h8):(2'h3)];
  assign wire1682 = reg1567;
  assign wire1683 = reg1608;
  always
    @(posedge clk) begin
      reg1684 <= reg1650[(3'h4):(3'h4)];
      for (forvar1685 = (1'h0); (forvar1685 < (2'h3)); forvar1685 = (forvar1685 + (1'h1)))
        begin
          reg1686 <= $signed((($unsigned(reg1622) ?
              (reg1639 >>> reg1576) : (reg1541 ?
                  reg1548 : reg1581)) - reg1656));
        end
      if ((-reg1601))
        begin
          for (forvar1687 = (1'h0); (forvar1687 < (2'h2)); forvar1687 = (forvar1687 + (1'h1)))
            begin
              reg1688 <= $unsigned($unsigned({(reg1598 ? reg1564 : reg1642)}));
              for (forvar1689 = (1'h0); (forvar1689 < (2'h3)); forvar1689 = (forvar1689 + (1'h1)))
                begin
                  if ((|((~^(reg1662 >> reg1669)) ?
                      ((reg1582 ? (8'hba) : reg1664) ?
                          reg1569 : (^(8'hb9))) : $signed((reg1600 ^~ reg1579)))))
                    begin
                      reg1690 <= (+$signed((8'hb0)));
                      reg1691 <= reg1591;
                    end
                  else
                    begin
                      reg1690 <= $signed($unsigned($unsigned(reg1578[(4'ha):(2'h3)])));
                      reg1691 <= $signed(reg1589);
                      reg1692 <= ((~^reg1598[(1'h0):(1'h0)]) ?
                          ((^{reg1558}) >>> ((reg1630 ^~ reg1669) <= (8'h9c))) : reg1657);
                    end
                  reg1693 <= (reg1639 ?
                      reg1639 : (((reg1603 || reg1665) ?
                          (reg1576 ?
                              reg1639 : wire1682) : reg1552[(3'h6):(2'h3)]) >= ((~(8'ha7)) ?
                          (-reg1564) : (reg1554 ? (8'hb1) : reg1546))));
                  if (((|$signed(reg1540[(3'h4):(2'h2)])) >>> reg1646))
                    begin
                      reg1694 <= $unsigned((-{(reg1646 ?
                              reg1605 : forvar1685)}));
                      reg1695 <= reg1546[(2'h3):(2'h3)];
                      reg1696 <= (~reg1549[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg1694 <= (^$signed(reg1549[(3'h4):(2'h2)]));
                      reg1695 <= $signed($signed(reg1643));
                      reg1696 <= (($signed($unsigned(reg1545)) ?
                          reg1555 : $unsigned({(8'hb8)})) <<< forvar1685[(4'hb):(3'h6)]);
                      reg1697 <= $unsigned($unsigned((8'hb5)));
                    end
                end
              for (forvar1698 = (1'h0); (forvar1698 < (2'h3)); forvar1698 = (forvar1698 + (1'h1)))
                begin
                  for (forvar1699 = (1'h0); (forvar1699 < (2'h3)); forvar1699 = (forvar1699 + (1'h1)))
                    begin
                      reg1700 <= reg1630;
                      reg1701 <= reg1542;
                      reg1702 <= {reg1690};
                    end
                  if (((wire1682 && reg1669) ?
                      (({reg1648} ? $unsigned((8'hae)) : reg1656) ?
                          (reg1613[(4'hc):(1'h0)] <<< reg1583[(4'h8):(3'h7)]) : ($unsigned(reg1606) & (reg1608 != reg1677))) : ((!$unsigned((8'ha4))) & reg1650[(3'h4):(2'h3)])))
                    begin
                      reg1703 <= ($unsigned((!(reg1565 ? reg1584 : reg1568))) ?
                          reg1587 : reg1601);
                      reg1704 <= (-{$unsigned($signed(reg1589))});
                      reg1705 <= $signed($unsigned((reg1670[(4'h8):(3'h7)] ?
                          (^reg1582) : reg1549[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg1703 <= (+{($signed(reg1546) ?
                              (reg1667 != wire1173) : $signed(reg1666))});
                      reg1704 <= $unsigned(($unsigned(reg1591[(4'hf):(4'hb)]) ?
                          reg1690[(2'h3):(2'h2)] : $signed($unsigned(reg1620))));
                    end
                end
              reg1706 <= reg1602[(2'h2):(1'h0)];
            end
          for (forvar1707 = (1'h0); (forvar1707 < (2'h2)); forvar1707 = (forvar1707 + (1'h1)))
            begin
              reg1708 <= ((-({(8'ha6)} ?
                  reg1547 : (reg1548 ?
                      reg1706 : (8'hb7)))) << $unsigned(reg1555[(1'h0):(1'h0)]));
              reg1709 <= (reg1543 >> ((reg1637[(4'h9):(1'h0)] > $signed(reg1612)) ?
                  (^~$signed(reg1598)) : (8'hb0)));
              for (forvar1710 = (1'h0); (forvar1710 < (1'h0)); forvar1710 = (forvar1710 + (1'h1)))
                begin
                  reg1711 <= $signed($unsigned((-(reg1549 ^~ reg1644))));
                end
            end
          for (forvar1712 = (1'h0); (forvar1712 < (2'h2)); forvar1712 = (forvar1712 + (1'h1)))
            begin
              reg1713 <= $unsigned($signed(reg1675));
              if (reg1688)
                begin
                  reg1714 <= reg1678[(1'h1):(1'h0)];
                  if ($unsigned(wire1174[(1'h0):(1'h0)]))
                    begin
                      reg1715 <= reg1617[(1'h0):(1'h0)];
                      reg1716 <= $unsigned(reg1640);
                      reg1717 <= reg1680;
                    end
                  else
                    begin
                      reg1715 <= (8'hab);
                      reg1716 <= $signed((~reg1696[(1'h0):(1'h0)]));
                    end
                  for (forvar1718 = (1'h0); (forvar1718 < (2'h3)); forvar1718 = (forvar1718 + (1'h1)))
                    begin
                      reg1719 <= ((reg1639 ?
                          (reg1636 <<< reg1714[(3'h4):(2'h3)]) : {(^~reg1548)}) ~^ (((~&reg1598) << (reg1640 ?
                              reg1693 : (8'hb5))) ?
                          reg1608[(1'h1):(1'h1)] : reg1700));
                      reg1720 <= reg1649;
                      reg1721 <= $signed($unsigned(reg1567[(3'h5):(3'h4)]));
                      reg1722 <= (((+forvar1718) ?
                          reg1702 : $unsigned($unsigned(reg1672))) >>> (|($unsigned(reg1558) ?
                          $signed(reg1690) : {reg1641})));
                    end
                end
              else
                begin
                  for (forvar1714 = (1'h0); (forvar1714 < (2'h2)); forvar1714 = (forvar1714 + (1'h1)))
                    begin
                      reg1715 <= ((~&reg1561) ?
                          $signed(($signed(reg1649) ~^ (reg1587 != reg1715))) : (reg1714[(1'h0):(1'h0)] >>> (8'hb5)));
                      reg1716 <= reg1557[(2'h2):(1'h1)];
                      reg1717 <= reg1660[(1'h1):(1'h0)];
                    end
                  for (forvar1718 = (1'h0); (forvar1718 < (2'h3)); forvar1718 = (forvar1718 + (1'h1)))
                    begin
                      reg1719 <= reg1555[(2'h2):(1'h1)];
                    end
                end
            end
        end
      else
        begin
          if ((~reg1720[(1'h0):(1'h0)]))
            begin
              for (forvar1687 = (1'h0); (forvar1687 < (1'h1)); forvar1687 = (forvar1687 + (1'h1)))
                begin
                  for (forvar1688 = (1'h0); (forvar1688 < (2'h2)); forvar1688 = (forvar1688 + (1'h1)))
                    begin
                      reg1689 <= (wire1175 ?
                          ((^$signed(reg1715)) << {wire1174}) : (^~$unsigned($signed(reg1564))));
                      reg1690 <= ((($signed(reg1679) ~^ (reg1686 != reg1716)) ?
                          reg1689 : (!$signed(reg1640))) - (($unsigned(reg1648) & (reg1672 && reg1577)) ?
                          reg1719[(1'h1):(1'h1)] : $unsigned((~^(8'hb3)))));
                      reg1691 <= (~|reg1686[(2'h3):(2'h2)]);
                    end
                  reg1692 <= ((&(~^(reg1662 * reg1570))) >= (~(^(reg1606 != reg1596))));
                  reg1693 <= reg1714[(3'h4):(1'h0)];
                end
              for (forvar1694 = (1'h0); (forvar1694 < (2'h3)); forvar1694 = (forvar1694 + (1'h1)))
                begin
                  for (forvar1695 = (1'h0); (forvar1695 < (2'h2)); forvar1695 = (forvar1695 + (1'h1)))
                    begin
                      reg1696 <= ((-($unsigned(reg1661) != (reg1599 ?
                          reg1554 : reg1617))) == ((reg1587[(2'h3):(2'h2)] ?
                          reg1637[(1'h1):(1'h0)] : (8'ha4)) << ($signed(reg1543) >>> reg1700[(2'h2):(1'h1)])));
                    end
                end
            end
          else
            begin
              for (forvar1687 = (1'h0); (forvar1687 < (2'h2)); forvar1687 = (forvar1687 + (1'h1)))
                begin
                  reg1688 <= $unsigned($unsigned((reg1600[(3'h6):(2'h3)] ?
                      (+reg1650) : ((8'ha1) <= reg1688))));
                  for (forvar1689 = (1'h0); (forvar1689 < (2'h2)); forvar1689 = (forvar1689 + (1'h1)))
                    begin
                      reg1690 <= reg1665[(3'h5):(3'h4)];
                      reg1691 <= $unsigned(reg1635[(3'h7):(3'h6)]);
                      reg1692 <= (8'hb8);
                      reg1693 <= $unsigned($unsigned(reg1579));
                    end
                  for (forvar1694 = (1'h0); (forvar1694 < (1'h1)); forvar1694 = (forvar1694 + (1'h1)))
                    begin
                      reg1695 <= ($unsigned(($unsigned((8'hb9)) ?
                          reg1552[(4'he):(4'h8)] : (reg1608 && reg1558))) * $unsigned((wire1172[(1'h0):(1'h0)] ?
                          $signed((8'hb6)) : (reg1622 ? reg1599 : (8'haf)))));
                    end
                end
              for (forvar1696 = (1'h0); (forvar1696 < (2'h3)); forvar1696 = (forvar1696 + (1'h1)))
                begin
                  if ((reg1555[(1'h0):(1'h0)] >> ((8'ha5) >> {$unsigned((8'hb5))})))
                    begin
                      reg1697 <= reg1717[(3'h7):(2'h3)];
                      reg1698 <= forvar1710;
                      reg1699 <= ((^{$signed(reg1568)}) < reg1623[(1'h1):(1'h1)]);
                      reg1700 <= reg1705[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg1697 <= reg1688;
                      reg1698 <= $signed($unsigned(((reg1628 ?
                              (8'hb5) : reg1704) ?
                          {reg1676} : $signed(forvar1695))));
                      reg1699 <= (8'h9d);
                    end
                  reg1701 <= reg1631[(3'h4):(1'h1)];
                  for (forvar1702 = (1'h0); (forvar1702 < (1'h1)); forvar1702 = (forvar1702 + (1'h1)))
                    begin
                      reg1703 <= (reg1713[(3'h6):(3'h4)] ?
                          $signed(reg1634) : ((^(reg1589 ?
                              reg1679 : reg1546)) < {$unsigned((8'ha5))}));
                      reg1704 <= ({reg1639[(4'h9):(2'h3)]} != reg1711[(4'h8):(2'h3)]);
                      reg1705 <= reg1640;
                      reg1706 <= reg1695;
                    end
                end
            end
          reg1707 <= reg1689[(1'h1):(1'h0)];
          for (forvar1708 = (1'h0); (forvar1708 < (2'h3)); forvar1708 = (forvar1708 + (1'h1)))
            begin
              if ($signed((($unsigned((8'h9d)) >>> (reg1719 ?
                  reg1713 : reg1692)) || reg1609[(1'h0):(1'h0)])))
                begin
                  for (forvar1709 = (1'h0); (forvar1709 < (2'h3)); forvar1709 = (forvar1709 + (1'h1)))
                    begin
                      reg1710 <= wire1174[(2'h3):(2'h2)];
                      reg1711 <= (((reg1641[(2'h3):(1'h0)] ~^ (8'ha7)) != reg1702) ?
                          reg1615 : (+reg1593));
                      reg1712 <= (8'ha7);
                    end
                  if (($signed(((reg1545 == reg1612) ?
                      $signed(reg1669) : $unsigned(reg1676))) * reg1644[(3'h4):(2'h3)]))
                    begin
                      reg1713 <= $unsigned(reg1642);
                      reg1714 <= (&(^(reg1553 ?
                          $signed(reg1721) : (~&reg1635))));
                    end
                  else
                    begin
                      reg1713 <= (8'had);
                      reg1714 <= reg1702[(4'ha):(2'h3)];
                      reg1715 <= (8'ha0);
                    end
                  reg1716 <= reg1577;
                  if (wire1178)
                    begin
                      reg1717 <= $unsigned((|(~reg1680[(1'h0):(1'h0)])));
                      reg1718 <= (~^{$unsigned($unsigned(reg1543))});
                      reg1719 <= $unsigned(reg1704[(4'hc):(4'h8)]);
                      reg1720 <= $signed($signed($signed((reg1555 ^~ reg1706))));
                    end
                  else
                    begin
                      reg1717 <= (&reg1652[(1'h0):(1'h0)]);
                      reg1718 <= $signed((reg1623[(2'h3):(2'h2)] * (&$signed(reg1559))));
                      reg1719 <= reg1667;
                    end
                end
              else
                begin
                  reg1709 <= reg1597;
                  for (forvar1710 = (1'h0); (forvar1710 < (1'h0)); forvar1710 = (forvar1710 + (1'h1)))
                    begin
                      reg1711 <= {forvar1695[(4'he):(4'hb)]};
                      reg1712 <= $unsigned((reg1710[(4'hc):(4'hc)] & $unsigned((+reg1554))));
                      reg1713 <= reg1718[(4'he):(2'h3)];
                      reg1714 <= reg1706;
                    end
                  reg1715 <= ($unsigned(reg1684[(1'h1):(1'h1)]) ?
                      reg1696[(1'h0):(1'h0)] : reg1714);
                end
              for (forvar1721 = (1'h0); (forvar1721 < (1'h0)); forvar1721 = (forvar1721 + (1'h1)))
                begin
                  if (($unsigned(reg1647[(4'hc):(4'hb)]) || (~&$signed((!reg1617)))))
                    begin
                      reg1722 <= ($signed((~(reg1584 ?
                          reg1599 : reg1581))) & $signed(((reg1599 ?
                              reg1720 : reg1591) ?
                          (reg1568 ?
                              reg1613 : reg1579) : (reg1674 == reg1692))));
                    end
                  else
                    begin
                      reg1722 <= {$signed(reg1597[(1'h0):(1'h0)])};
                      reg1723 <= (reg1709[(2'h3):(2'h2)] ?
                          $signed(((forvar1709 >>> reg1549) >> reg1555[(1'h0):(1'h0)])) : $unsigned($unsigned((-reg1677))));
                    end
                  for (forvar1724 = (1'h0); (forvar1724 < (1'h0)); forvar1724 = (forvar1724 + (1'h1)))
                    begin
                      reg1725 <= $unsigned(((8'hb0) | ((^~wire1683) ?
                          reg1712 : (reg1614 ? reg1718 : reg1539))));
                      reg1726 <= (reg1709 ?
                          ($signed($signed((8'hb9))) ~^ reg1567) : reg1539);
                      reg1727 <= reg1623;
                    end
                  for (forvar1728 = (1'h0); (forvar1728 < (1'h0)); forvar1728 = (forvar1728 + (1'h1)))
                    begin
                      reg1729 <= $unsigned($signed(reg1557[(1'h0):(1'h0)]));
                      reg1730 <= (((reg1559[(4'h9):(3'h4)] << reg1644[(3'h6):(3'h4)]) ?
                              reg1637 : reg1539) ?
                          (((|reg1632) < $unsigned(reg1696)) ?
                              ((reg1635 ? reg1557 : wire1174) ?
                                  (reg1557 ^~ reg1607) : (reg1618 ?
                                      (8'ha0) : reg1711)) : ($unsigned(reg1600) ?
                                  $signed(reg1567) : $signed(reg1569))) : reg1678);
                    end
                end
            end
        end
      for (forvar1731 = (1'h0); (forvar1731 < (2'h3)); forvar1731 = (forvar1731 + (1'h1)))
        begin
          for (forvar1732 = (1'h0); (forvar1732 < (2'h2)); forvar1732 = (forvar1732 + (1'h1)))
            begin
              if (((forvar1689[(2'h2):(2'h2)] ?
                      reg1559 : (((8'hb0) <= reg1542) ?
                          reg1547 : (reg1692 > (8'had)))) ?
                  forvar1718[(2'h3):(2'h2)] : $unsigned(((wire1174 ?
                          reg1628 : reg1684) ?
                      $unsigned(forvar1710) : (reg1538 >= reg1699)))))
                begin
                  reg1733 <= wire1174[(2'h2):(1'h1)];
                  for (forvar1734 = (1'h0); (forvar1734 < (1'h0)); forvar1734 = (forvar1734 + (1'h1)))
                    begin
                      reg1735 <= ((~$signed((reg1573 ?
                          reg1592 : reg1712))) && reg1543);
                      reg1736 <= {(reg1688[(2'h3):(2'h3)] ?
                              (~&(~&reg1591)) : {(reg1710 >= forvar1734)})};
                      reg1737 <= $unsigned(($signed(forvar1698) << $signed((forvar1699 ?
                          reg1710 : reg1684))));
                      reg1738 <= {(^~(+$signed(reg1695)))};
                    end
                end
              else
                begin
                  reg1733 <= ((reg1555[(1'h1):(1'h1)] ?
                      (8'ha8) : $signed((~&(8'hb3)))) <= $signed(((|reg1601) ?
                      $unsigned(forvar1732) : reg1546)));
                  if (((-$unsigned((reg1648 ? reg1727 : reg1733))) == reg1635))
                    begin
                      reg1734 <= $signed(reg1678[(2'h2):(1'h1)]);
                      reg1735 <= (reg1579[(2'h3):(2'h2)] ?
                          (!{(reg1694 ?
                                  reg1709 : reg1578)}) : {$unsigned($signed((8'hac)))});
                      reg1736 <= ((~|reg1628) > ((reg1559[(4'h8):(4'h8)] ?
                          $unsigned(reg1709) : reg1720[(1'h1):(1'h0)]) || $signed(forvar1710)));
                    end
                  else
                    begin
                      reg1734 <= (wire1177[(3'h6):(3'h4)] < $signed(((reg1656 && reg1670) * $signed(reg1722))));
                    end
                  reg1737 <= $signed(reg1633);
                  if ((!((+(^~reg1590)) ?
                      reg1719[(2'h2):(2'h2)] : ((reg1643 ^ reg1666) > reg1573))))
                    begin
                      reg1738 <= (~&reg1630[(4'h8):(2'h2)]);
                    end
                  else
                    begin
                      reg1738 <= (|reg1631);
                      reg1739 <= (reg1661 ?
                          reg1627[(2'h3):(1'h0)] : $signed(((^forvar1721) ?
                              {reg1606} : forvar1708[(4'h8):(3'h4)])));
                    end
                end
              if (reg1641[(2'h2):(1'h1)])
                begin
                  for (forvar1740 = (1'h0); (forvar1740 < (1'h0)); forvar1740 = (forvar1740 + (1'h1)))
                    begin
                      reg1741 <= $signed($unsigned(wire1172[(2'h3):(2'h2)]));
                      reg1742 <= forvar1708;
                      reg1743 <= $signed(reg1674);
                      reg1744 <= {(~&reg1730[(3'h7):(1'h1)])};
                    end
                end
              else
                begin
                  for (forvar1740 = (1'h0); (forvar1740 < (2'h3)); forvar1740 = (forvar1740 + (1'h1)))
                    begin
                      reg1741 <= ((^~(~^(forvar1688 >= (8'hb7)))) <= $signed(((|reg1641) ?
                          (forvar1694 << reg1661) : (forvar1731 ?
                              reg1547 : reg1581))));
                      reg1742 <= $unsigned({({reg1670} ?
                              (~|(8'hba)) : reg1691)});
                      reg1743 <= {$unsigned((~^(reg1605 >> reg1670)))};
                      reg1744 <= ((&((forvar1721 ~^ reg1722) ?
                              $unsigned((8'hb8)) : (reg1689 ^~ reg1613))) ?
                          reg1725[(2'h2):(2'h2)] : $unsigned(({(8'h9d)} ?
                              (wire1177 ? reg1675 : reg1539) : (reg1667 ?
                                  reg1628 : reg1590))));
                    end
                  reg1745 <= (|(($signed(reg1677) & reg1552) ?
                      (-$signed(reg1590)) : {(reg1628 ? reg1608 : reg1662)}));
                  reg1746 <= (reg1657 <= {$signed((^~reg1692))});
                  if (reg1717[(3'h4):(1'h1)])
                    begin
                      reg1747 <= reg1611[(3'h7):(3'h7)];
                      reg1748 <= reg1615[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg1747 <= reg1697;
                      reg1748 <= reg1581[(2'h2):(1'h0)];
                      reg1749 <= {(-reg1727)};
                      reg1750 <= $signed(((reg1719 ?
                              (reg1623 == forvar1694) : ((8'hb9) ?
                                  reg1555 : forvar1732)) ?
                          $signed(reg1680) : ({wire1172} ?
                              $unsigned(reg1546) : $unsigned(reg1718))));
                    end
                end
            end
        end
    end
  assign wire1751 = $signed(($unsigned((reg1673 ?
                        (8'ha0) : reg1557)) + reg1667[(1'h0):(1'h0)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module739
#(parameter param1085 = (({((8'h9d) ? (8'ha2) : (8'hba))} + ({(8'hab)} < ((8'haa) ^ (8'ha1)))) * (((^~(8'had)) == (^(8'h9f))) ? (!((8'h9d) ? (8'hb4) : (8'ha0))) : (-(8'hb6)))))
(y, clk, wire743, wire742, wire741, wire740);
  output wire [(32'hdbe):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire743;
  input wire signed [(4'ha):(1'h0)] wire742;
  input wire signed [(4'hb):(1'h0)] wire741;
  input wire [(4'hd):(1'h0)] wire740;
  wire [(2'h3):(1'h0)] wire838;
  wire signed [(4'h9):(1'h0)] wire745;
  wire [(4'hc):(1'h0)] wire744;
  reg signed [(4'h8):(1'h0)] reg1084 = (1'h0);
  reg [(3'h5):(1'h0)] reg1083 = (1'h0);
  reg [(3'h6):(1'h0)] reg1082 = (1'h0);
  reg [(4'hd):(1'h0)] reg1081 = (1'h0);
  reg [(3'h5):(1'h0)] reg1079 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1057 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1069 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1077 = (1'h0);
  reg [(3'h7):(1'h0)] reg1076 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1075 = (1'h0);
  reg [(4'he):(1'h0)] reg1074 = (1'h0);
  reg [(3'h7):(1'h0)] reg1072 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1071 = (1'h0);
  reg [(4'h9):(1'h0)] reg1070 = (1'h0);
  reg [(3'h4):(1'h0)] reg1068 = (1'h0);
  reg [(4'hf):(1'h0)] reg1067 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1066 = (1'h0);
  reg [(4'h8):(1'h0)] reg1065 = (1'h0);
  reg [(5'h10):(1'h0)] reg1063 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1062 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1061 = (1'h0);
  reg [(4'hd):(1'h0)] reg1060 = (1'h0);
  reg [(4'he):(1'h0)] reg1059 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1058 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1056 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1055 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1054 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1053 = (1'h0);
  reg [(4'h8):(1'h0)] reg1051 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1046 = (1'h0);
  reg [(4'hd):(1'h0)] reg1044 = (1'h0);
  reg [(4'hf):(1'h0)] reg1042 = (1'h0);
  reg [(4'he):(1'h0)] reg1050 = (1'h0);
  reg [(4'he):(1'h0)] reg1049 = (1'h0);
  reg [(3'h4):(1'h0)] reg1048 = (1'h0);
  reg [(4'he):(1'h0)] reg1047 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1045 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1043 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1041 = (1'h0);
  reg [(4'he):(1'h0)] reg1040 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1038 = (1'h0);
  reg [(4'hc):(1'h0)] reg1037 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1035 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1034 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1032 = (1'h0);
  reg [(4'hd):(1'h0)] reg1031 = (1'h0);
  reg [(2'h2):(1'h0)] reg1030 = (1'h0);
  reg [(3'h7):(1'h0)] reg1029 = (1'h0);
  reg [(4'h9):(1'h0)] reg1026 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1025 = (1'h0);
  reg [(5'h10):(1'h0)] reg1024 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1023 = (1'h0);
  reg [(4'hc):(1'h0)] reg1011 = (1'h0);
  reg [(4'hc):(1'h0)] reg1006 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1019 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1018 = (1'h0);
  reg [(4'h8):(1'h0)] reg1017 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1016 = (1'h0);
  reg [(4'ha):(1'h0)] reg1014 = (1'h0);
  reg [(4'he):(1'h0)] reg1013 = (1'h0);
  reg [(5'h10):(1'h0)] reg1012 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1003 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1010 = (1'h0);
  reg [(4'ha):(1'h0)] reg1009 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1008 = (1'h0);
  reg [(4'ha):(1'h0)] reg1007 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1005 = (1'h0);
  reg [(2'h3):(1'h0)] reg1004 = (1'h0);
  reg [(4'hc):(1'h0)] reg1002 = (1'h0);
  reg [(4'he):(1'h0)] reg1001 = (1'h0);
  reg [(4'hd):(1'h0)] reg1000 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg999 = (1'h0);
  reg [(4'hd):(1'h0)] reg998 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg996 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg995 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg994 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg993 = (1'h0);
  reg [(2'h3):(1'h0)] reg992 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg990 = (1'h0);
  reg [(4'h8):(1'h0)] reg989 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg988 = (1'h0);
  reg [(3'h7):(1'h0)] reg987 = (1'h0);
  reg [(3'h5):(1'h0)] reg985 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg986 = (1'h0);
  reg [(3'h4):(1'h0)] reg984 = (1'h0);
  reg [(4'h8):(1'h0)] reg983 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg982 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg981 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg978 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg977 = (1'h0);
  reg [(2'h2):(1'h0)] reg976 = (1'h0);
  reg [(4'he):(1'h0)] reg975 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg974 = (1'h0);
  reg [(3'h7):(1'h0)] reg973 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg970 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg972 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg971 = (1'h0);
  reg [(3'h7):(1'h0)] reg969 = (1'h0);
  reg [(4'hb):(1'h0)] reg968 = (1'h0);
  reg [(3'h4):(1'h0)] reg966 = (1'h0);
  reg [(4'hc):(1'h0)] reg965 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg964 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg963 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg962 = (1'h0);
  reg [(3'h4):(1'h0)] reg955 = (1'h0);
  reg [(4'hf):(1'h0)] reg954 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg952 = (1'h0);
  reg [(2'h2):(1'h0)] reg942 = (1'h0);
  reg signed [(4'he):(1'h0)] reg945 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg943 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg960 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg959 = (1'h0);
  reg [(4'hd):(1'h0)] reg958 = (1'h0);
  reg [(5'h10):(1'h0)] reg957 = (1'h0);
  reg [(2'h3):(1'h0)] reg956 = (1'h0);
  reg [(2'h3):(1'h0)] reg953 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg951 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg950 = (1'h0);
  reg [(4'ha):(1'h0)] reg949 = (1'h0);
  reg [(5'h10):(1'h0)] reg948 = (1'h0);
  reg [(4'h9):(1'h0)] reg947 = (1'h0);
  reg [(3'h4):(1'h0)] reg946 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg944 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg940 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg939 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg938 = (1'h0);
  reg [(3'h7):(1'h0)] reg937 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg936 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg935 = (1'h0);
  reg [(3'h7):(1'h0)] reg934 = (1'h0);
  reg [(4'hd):(1'h0)] reg932 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg931 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg930 = (1'h0);
  reg [(3'h4):(1'h0)] reg929 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg928 = (1'h0);
  reg [(3'h5):(1'h0)] reg927 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg926 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg925 = (1'h0);
  reg signed [(4'he):(1'h0)] reg923 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg922 = (1'h0);
  reg [(3'h5):(1'h0)] reg921 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg919 = (1'h0);
  reg [(4'hf):(1'h0)] reg918 = (1'h0);
  reg [(4'h9):(1'h0)] reg917 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg916 = (1'h0);
  reg signed [(4'he):(1'h0)] reg915 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg914 = (1'h0);
  reg [(4'ha):(1'h0)] reg913 = (1'h0);
  reg [(4'ha):(1'h0)] reg910 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg907 = (1'h0);
  reg [(4'hc):(1'h0)] reg912 = (1'h0);
  reg [(4'he):(1'h0)] reg911 = (1'h0);
  reg [(3'h4):(1'h0)] reg909 = (1'h0);
  reg [(4'he):(1'h0)] reg908 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg906 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg905 = (1'h0);
  reg signed [(4'he):(1'h0)] reg904 = (1'h0);
  reg signed [(4'he):(1'h0)] reg888 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg901 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg900 = (1'h0);
  reg [(3'h4):(1'h0)] reg898 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg897 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg896 = (1'h0);
  reg [(3'h5):(1'h0)] reg895 = (1'h0);
  reg [(2'h3):(1'h0)] reg894 = (1'h0);
  reg [(2'h3):(1'h0)] reg893 = (1'h0);
  reg [(4'h8):(1'h0)] reg892 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg891 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg890 = (1'h0);
  reg [(3'h6):(1'h0)] reg889 = (1'h0);
  reg [(4'h9):(1'h0)] reg886 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg885 = (1'h0);
  reg [(4'ha):(1'h0)] reg884 = (1'h0);
  reg [(4'hb):(1'h0)] reg883 = (1'h0);
  reg [(4'hb):(1'h0)] reg882 = (1'h0);
  reg [(3'h4):(1'h0)] reg881 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg880 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg875 = (1'h0);
  reg [(5'h10):(1'h0)] reg872 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg862 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg878 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg877 = (1'h0);
  reg [(5'h10):(1'h0)] reg876 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg874 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg873 = (1'h0);
  reg [(3'h4):(1'h0)] reg865 = (1'h0);
  reg [(2'h2):(1'h0)] reg871 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg870 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg869 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg868 = (1'h0);
  reg [(3'h5):(1'h0)] reg867 = (1'h0);
  reg [(3'h4):(1'h0)] reg866 = (1'h0);
  reg [(3'h4):(1'h0)] reg864 = (1'h0);
  reg [(4'hc):(1'h0)] reg863 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg861 = (1'h0);
  reg signed [(4'he):(1'h0)] reg860 = (1'h0);
  reg [(3'h4):(1'h0)] reg859 = (1'h0);
  reg [(3'h7):(1'h0)] reg858 = (1'h0);
  reg [(4'hc):(1'h0)] reg857 = (1'h0);
  reg [(3'h7):(1'h0)] reg855 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg854 = (1'h0);
  reg [(4'h8):(1'h0)] reg850 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg845 = (1'h0);
  reg [(4'ha):(1'h0)] reg853 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg852 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg851 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg849 = (1'h0);
  reg [(4'hb):(1'h0)] reg848 = (1'h0);
  reg [(4'h9):(1'h0)] reg847 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg846 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg844 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg840 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg837 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg836 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg835 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg833 = (1'h0);
  reg [(4'hf):(1'h0)] reg832 = (1'h0);
  reg signed [(4'he):(1'h0)] reg823 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg829 = (1'h0);
  reg signed [(4'he):(1'h0)] reg828 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg827 = (1'h0);
  reg [(2'h2):(1'h0)] reg826 = (1'h0);
  reg [(4'hf):(1'h0)] reg825 = (1'h0);
  reg [(4'ha):(1'h0)] reg824 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg822 = (1'h0);
  reg [(4'hf):(1'h0)] reg821 = (1'h0);
  reg [(3'h5):(1'h0)] reg820 = (1'h0);
  reg [(2'h2):(1'h0)] reg819 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg818 = (1'h0);
  reg [(4'ha):(1'h0)] reg817 = (1'h0);
  reg [(3'h7):(1'h0)] reg812 = (1'h0);
  reg [(4'he):(1'h0)] reg811 = (1'h0);
  reg [(4'hb):(1'h0)] reg810 = (1'h0);
  reg [(4'h8):(1'h0)] reg808 = (1'h0);
  reg [(3'h7):(1'h0)] reg807 = (1'h0);
  reg [(3'h5):(1'h0)] reg806 = (1'h0);
  reg [(3'h6):(1'h0)] reg805 = (1'h0);
  reg [(3'h4):(1'h0)] reg804 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg801 = (1'h0);
  reg [(5'h10):(1'h0)] reg800 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg799 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg798 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg797 = (1'h0);
  reg signed [(4'he):(1'h0)] reg794 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg788 = (1'h0);
  reg [(4'h9):(1'h0)] reg783 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg796 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg795 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg793 = (1'h0);
  reg [(2'h2):(1'h0)] reg792 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg791 = (1'h0);
  reg [(4'ha):(1'h0)] reg790 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg789 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg787 = (1'h0);
  reg [(4'hd):(1'h0)] reg786 = (1'h0);
  reg [(3'h7):(1'h0)] reg785 = (1'h0);
  reg [(3'h5):(1'h0)] reg784 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg782 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg771 = (1'h0);
  reg [(4'ha):(1'h0)] reg770 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg781 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg780 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg779 = (1'h0);
  reg [(3'h4):(1'h0)] reg778 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg777 = (1'h0);
  reg [(4'hd):(1'h0)] reg776 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg775 = (1'h0);
  reg [(4'hb):(1'h0)] reg774 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg773 = (1'h0);
  reg [(3'h5):(1'h0)] reg772 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg769 = (1'h0);
  reg [(4'he):(1'h0)] reg768 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg767 = (1'h0);
  reg [(5'h10):(1'h0)] reg765 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg764 = (1'h0);
  reg [(3'h6):(1'h0)] reg763 = (1'h0);
  reg [(2'h2):(1'h0)] reg761 = (1'h0);
  reg [(4'hb):(1'h0)] reg760 = (1'h0);
  reg signed [(4'he):(1'h0)] reg757 = (1'h0);
  reg [(4'hd):(1'h0)] reg756 = (1'h0);
  reg [(3'h4):(1'h0)] reg755 = (1'h0);
  reg [(3'h7):(1'h0)] reg754 = (1'h0);
  reg [(4'ha):(1'h0)] reg752 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg751 = (1'h0);
  reg [(3'h4):(1'h0)] reg750 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg749 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1080 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1078 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1058 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1070 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1068 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1066 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1073 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1069 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1064 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1057 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1052 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1048 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1045 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1046 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1044 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1042 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1039 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1029 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1036 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1033 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1028 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1027 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1022 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1021 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1020 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1008 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1004 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1015 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1011 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1006 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1003 = (1'h0);
  reg [(4'h9):(1'h0)] forvar997 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar992 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar991 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar985 = (1'h0);
  reg [(4'hc):(1'h0)] forvar980 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar979 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar968 = (1'h0);
  reg [(5'h10):(1'h0)] forvar970 = (1'h0);
  reg [(4'h8):(1'h0)] forvar967 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar961 = (1'h0);
  reg [(4'h8):(1'h0)] forvar960 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar958 = (1'h0);
  reg [(4'hc):(1'h0)] forvar957 = (1'h0);
  reg [(5'h10):(1'h0)] forvar953 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar948 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar955 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar954 = (1'h0);
  reg [(3'h4):(1'h0)] forvar952 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar945 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar943 = (1'h0);
  reg [(4'h8):(1'h0)] forvar942 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar941 = (1'h0);
  reg [(5'h10):(1'h0)] forvar938 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar925 = (1'h0);
  reg [(4'hc):(1'h0)] forvar933 = (1'h0);
  reg [(4'ha):(1'h0)] forvar928 = (1'h0);
  reg [(3'h5):(1'h0)] forvar926 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar924 = (1'h0);
  reg [(4'hd):(1'h0)] forvar920 = (1'h0);
  reg [(3'h6):(1'h0)] forvar910 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar907 = (1'h0);
  reg [(4'hb):(1'h0)] forvar903 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar902 = (1'h0);
  reg [(4'hc):(1'h0)] forvar889 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar899 = (1'h0);
  reg [(4'h8):(1'h0)] forvar888 = (1'h0);
  reg [(5'h10):(1'h0)] forvar887 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar879 = (1'h0);
  reg [(4'hd):(1'h0)] forvar874 = (1'h0);
  reg [(2'h3):(1'h0)] forvar860 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar863 = (1'h0);
  reg [(3'h5):(1'h0)] forvar857 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar875 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar872 = (1'h0);
  reg [(5'h10):(1'h0)] forvar865 = (1'h0);
  reg [(2'h2):(1'h0)] forvar862 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar856 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar851 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar850 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar845 = (1'h0);
  reg [(3'h4):(1'h0)] forvar843 = (1'h0);
  reg [(3'h7):(1'h0)] forvar842 = (1'h0);
  reg [(4'he):(1'h0)] forvar841 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar839 = (1'h0);
  reg [(4'hd):(1'h0)] forvar834 = (1'h0);
  reg [(4'h9):(1'h0)] forvar831 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar830 = (1'h0);
  reg [(3'h6):(1'h0)] forvar823 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar816 = (1'h0);
  reg [(3'h5):(1'h0)] forvar815 = (1'h0);
  reg [(4'hb):(1'h0)] forvar814 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar813 = (1'h0);
  reg [(4'h9):(1'h0)] forvar809 = (1'h0);
  reg [(2'h2):(1'h0)] forvar803 = (1'h0);
  reg [(3'h4):(1'h0)] forvar802 = (1'h0);
  reg [(4'hb):(1'h0)] forvar797 = (1'h0);
  reg [(4'hc):(1'h0)] forvar791 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar794 = (1'h0);
  reg [(3'h4):(1'h0)] forvar788 = (1'h0);
  reg [(4'hd):(1'h0)] forvar783 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar772 = (1'h0);
  reg [(4'ha):(1'h0)] forvar769 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar771 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar770 = (1'h0);
  reg [(4'hb):(1'h0)] forvar766 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar762 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar759 = (1'h0);
  reg [(2'h3):(1'h0)] forvar758 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar753 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar748 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar747 = (1'h0);
  reg [(4'hc):(1'h0)] forvar746 = (1'h0);
  assign y = {wire838,
                 wire745,
                 wire744,
                 reg1084,
                 reg1083,
                 reg1082,
                 reg1081,
                 reg1079,
                 reg1057,
                 reg1069,
                 reg1077,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg1072,
                 reg1071,
                 reg1070,
                 reg1068,
                 reg1067,
                 reg1066,
                 reg1065,
                 reg1063,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 reg1056,
                 reg1055,
                 reg1054,
                 reg1053,
                 reg1051,
                 reg1046,
                 reg1044,
                 reg1042,
                 reg1050,
                 reg1049,
                 reg1048,
                 reg1047,
                 reg1045,
                 reg1043,
                 reg1041,
                 reg1040,
                 reg1038,
                 reg1037,
                 reg1035,
                 reg1034,
                 reg1032,
                 reg1031,
                 reg1030,
                 reg1029,
                 reg1026,
                 reg1025,
                 reg1024,
                 reg1023,
                 reg1011,
                 reg1006,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1016,
                 reg1014,
                 reg1013,
                 reg1012,
                 reg1003,
                 reg1010,
                 reg1009,
                 reg1008,
                 reg1007,
                 reg1005,
                 reg1004,
                 reg1002,
                 reg1001,
                 reg1000,
                 reg999,
                 reg998,
                 reg996,
                 reg995,
                 reg994,
                 reg993,
                 reg992,
                 reg990,
                 reg989,
                 reg988,
                 reg987,
                 reg985,
                 reg986,
                 reg984,
                 reg983,
                 reg982,
                 reg981,
                 reg978,
                 reg977,
                 reg976,
                 reg975,
                 reg974,
                 reg973,
                 reg970,
                 reg972,
                 reg971,
                 reg969,
                 reg968,
                 reg966,
                 reg965,
                 reg964,
                 reg963,
                 reg962,
                 reg955,
                 reg954,
                 reg952,
                 reg942,
                 reg945,
                 reg943,
                 reg960,
                 reg959,
                 reg958,
                 reg957,
                 reg956,
                 reg953,
                 reg951,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 reg946,
                 reg944,
                 reg940,
                 reg939,
                 reg938,
                 reg937,
                 reg936,
                 reg935,
                 reg934,
                 reg932,
                 reg931,
                 reg930,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 reg925,
                 reg923,
                 reg922,
                 reg921,
                 reg919,
                 reg918,
                 reg917,
                 reg916,
                 reg915,
                 reg914,
                 reg913,
                 reg910,
                 reg907,
                 reg912,
                 reg911,
                 reg909,
                 reg908,
                 reg906,
                 reg905,
                 reg904,
                 reg888,
                 reg901,
                 reg900,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 reg889,
                 reg886,
                 reg885,
                 reg884,
                 reg883,
                 reg882,
                 reg881,
                 reg880,
                 reg875,
                 reg872,
                 reg862,
                 reg878,
                 reg877,
                 reg876,
                 reg874,
                 reg873,
                 reg865,
                 reg871,
                 reg870,
                 reg869,
                 reg868,
                 reg867,
                 reg866,
                 reg864,
                 reg863,
                 reg861,
                 reg860,
                 reg859,
                 reg858,
                 reg857,
                 reg855,
                 reg854,
                 reg850,
                 reg845,
                 reg853,
                 reg852,
                 reg851,
                 reg849,
                 reg848,
                 reg847,
                 reg846,
                 reg844,
                 reg840,
                 reg837,
                 reg836,
                 reg835,
                 reg833,
                 reg832,
                 reg823,
                 reg829,
                 reg828,
                 reg827,
                 reg826,
                 reg825,
                 reg824,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 reg818,
                 reg817,
                 reg812,
                 reg811,
                 reg810,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg801,
                 reg800,
                 reg799,
                 reg798,
                 reg797,
                 reg794,
                 reg788,
                 reg783,
                 reg796,
                 reg795,
                 reg793,
                 reg792,
                 reg791,
                 reg790,
                 reg789,
                 reg787,
                 reg786,
                 reg785,
                 reg784,
                 reg782,
                 reg771,
                 reg770,
                 reg781,
                 reg780,
                 reg779,
                 reg778,
                 reg777,
                 reg776,
                 reg775,
                 reg774,
                 reg773,
                 reg772,
                 reg769,
                 reg768,
                 reg767,
                 reg765,
                 reg764,
                 reg763,
                 reg761,
                 reg760,
                 reg757,
                 reg756,
                 reg755,
                 reg754,
                 reg752,
                 reg751,
                 reg750,
                 reg749,
                 forvar1080,
                 forvar1078,
                 forvar1058,
                 forvar1070,
                 forvar1068,
                 forvar1066,
                 forvar1073,
                 forvar1069,
                 forvar1064,
                 forvar1057,
                 forvar1052,
                 forvar1048,
                 forvar1045,
                 forvar1046,
                 forvar1044,
                 forvar1042,
                 forvar1039,
                 forvar1029,
                 forvar1036,
                 forvar1033,
                 forvar1028,
                 forvar1027,
                 forvar1022,
                 forvar1021,
                 forvar1020,
                 forvar1008,
                 forvar1004,
                 forvar1015,
                 forvar1011,
                 forvar1006,
                 forvar1003,
                 forvar997,
                 forvar992,
                 forvar991,
                 forvar985,
                 forvar980,
                 forvar979,
                 forvar968,
                 forvar970,
                 forvar967,
                 forvar961,
                 forvar960,
                 forvar958,
                 forvar957,
                 forvar953,
                 forvar948,
                 forvar955,
                 forvar954,
                 forvar952,
                 forvar945,
                 forvar943,
                 forvar942,
                 forvar941,
                 forvar938,
                 forvar925,
                 forvar933,
                 forvar928,
                 forvar926,
                 forvar924,
                 forvar920,
                 forvar910,
                 forvar907,
                 forvar903,
                 forvar902,
                 forvar889,
                 forvar899,
                 forvar888,
                 forvar887,
                 forvar879,
                 forvar874,
                 forvar860,
                 forvar863,
                 forvar857,
                 forvar875,
                 forvar872,
                 forvar865,
                 forvar862,
                 forvar856,
                 forvar851,
                 forvar850,
                 forvar845,
                 forvar843,
                 forvar842,
                 forvar841,
                 forvar839,
                 forvar834,
                 forvar831,
                 forvar830,
                 forvar823,
                 forvar816,
                 forvar815,
                 forvar814,
                 forvar813,
                 forvar809,
                 forvar803,
                 forvar802,
                 forvar797,
                 forvar791,
                 forvar794,
                 forvar788,
                 forvar783,
                 forvar772,
                 forvar769,
                 forvar771,
                 forvar770,
                 forvar766,
                 forvar762,
                 forvar759,
                 forvar758,
                 forvar753,
                 forvar748,
                 forvar747,
                 forvar746,
                 (1'h0)};
  assign wire744 = wire743;
  assign wire745 = {wire744};
  always
    @(posedge clk) begin
      for (forvar746 = (1'h0); (forvar746 < (1'h0)); forvar746 = (forvar746 + (1'h1)))
        begin
          for (forvar747 = (1'h0); (forvar747 < (2'h2)); forvar747 = (forvar747 + (1'h1)))
            begin
              for (forvar748 = (1'h0); (forvar748 < (2'h2)); forvar748 = (forvar748 + (1'h1)))
                begin
                  if (wire744)
                    begin
                      reg749 <= ($unsigned(wire740[(1'h1):(1'h0)]) <= $unsigned((wire741 << wire743)));
                      reg750 <= $signed((wire743 ^ $unsigned(((8'hac) || wire742))));
                      reg751 <= ((&$signed((reg750 >= wire741))) ?
                          wire742 : $signed(($signed(forvar748) >= forvar748[(1'h0):(1'h0)])));
                      reg752 <= (forvar746[(1'h0):(1'h0)] ^~ {$unsigned({reg750})});
                    end
                  else
                    begin
                      reg749 <= ((~$unsigned($unsigned(wire742))) * $unsigned(reg750[(1'h0):(1'h0)]));
                      reg750 <= (~(^{{wire743}}));
                    end
                  for (forvar753 = (1'h0); (forvar753 < (1'h1)); forvar753 = (forvar753 + (1'h1)))
                    begin
                      reg754 <= (($signed((wire740 ?
                          wire740 : forvar753)) && (|$unsigned(reg752))) > ((wire740[(3'h4):(2'h3)] ?
                          (|forvar748) : forvar753) | $unsigned($signed(wire743))));
                      reg755 <= $unsigned(($unsigned(((8'ha4) & wire741)) >> {(wire744 ?
                              wire740 : wire744)}));
                    end
                  reg756 <= ((($signed(wire744) ?
                          $signed(forvar748) : (reg749 ? forvar748 : reg750)) ?
                      ((~^reg749) ?
                          (wire745 ?
                              reg749 : wire745) : $signed(wire745)) : (|$unsigned(reg749))) <<< wire742);
                end
              reg757 <= wire745[(3'h7):(1'h0)];
              for (forvar758 = (1'h0); (forvar758 < (1'h1)); forvar758 = (forvar758 + (1'h1)))
                begin
                  for (forvar759 = (1'h0); (forvar759 < (2'h2)); forvar759 = (forvar759 + (1'h1)))
                    begin
                      reg760 <= reg755[(2'h3):(2'h2)];
                      reg761 <= reg757;
                    end
                  for (forvar762 = (1'h0); (forvar762 < (1'h1)); forvar762 = (forvar762 + (1'h1)))
                    begin
                      reg763 <= ((($signed(reg756) >= forvar762[(1'h0):(1'h0)]) >>> $unsigned((wire741 << wire741))) & ((forvar753 ?
                          $signed(reg755) : reg760) * (|(~|wire741))));
                      reg764 <= $unsigned($signed((|reg751[(4'hb):(3'h7)])));
                      reg765 <= $signed($unsigned((reg750 ?
                          (~^wire742) : reg749)));
                    end
                end
              for (forvar766 = (1'h0); (forvar766 < (1'h0)); forvar766 = (forvar766 + (1'h1)))
                begin
                  if ($unsigned({(~(|reg756))}))
                    begin
                      reg767 <= wire743[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg767 <= (8'hb9);
                    end
                  reg768 <= ((($signed(reg754) ?
                          (&wire744) : $signed(reg763)) || wire743) ?
                      reg763[(2'h2):(1'h1)] : wire741);
                end
            end
          if ($unsigned(reg761[(1'h0):(1'h0)]))
            begin
              reg769 <= $unsigned(forvar746[(2'h2):(1'h1)]);
              for (forvar770 = (1'h0); (forvar770 < (1'h1)); forvar770 = (forvar770 + (1'h1)))
                begin
                  for (forvar771 = (1'h0); (forvar771 < (1'h0)); forvar771 = (forvar771 + (1'h1)))
                    begin
                      reg772 <= $unsigned($signed($signed($unsigned(forvar762))));
                      reg773 <= $signed(forvar753);
                      reg774 <= wire744;
                      reg775 <= (forvar770[(3'h5):(3'h4)] || (forvar746 ?
                          {(^reg752)} : forvar747[(3'h5):(1'h0)]));
                    end
                  if (((^forvar766) + {((~&wire742) ?
                          {reg750} : $unsigned(reg750))}))
                    begin
                      reg776 <= $unsigned($signed($unsigned(((8'hb2) < (8'hb6)))));
                      reg777 <= (8'hb9);
                    end
                  else
                    begin
                      reg776 <= ((((~^(8'ha9)) || forvar759[(2'h3):(2'h2)]) ?
                          ($unsigned(wire744) + ((8'hb9) ?
                              reg760 : forvar762)) : ($unsigned((8'hba)) ?
                              (wire740 ?
                                  reg767 : reg752) : $unsigned(reg763))) < forvar762[(1'h0):(1'h0)]);
                      reg777 <= (~|wire745);
                      reg778 <= $signed((+reg777));
                    end
                  reg779 <= (~wire741[(3'h5):(1'h0)]);
                  if ($unsigned($signed({reg752})))
                    begin
                      reg780 <= (wire740 ? reg757[(4'hb):(2'h2)] : forvar753);
                      reg781 <= ($unsigned($unsigned(wire741)) | (reg752 ?
                          reg764[(4'ha):(4'h8)] : {$signed(reg751)}));
                    end
                  else
                    begin
                      reg780 <= ($signed((reg769 * (reg767 + wire744))) && $signed({reg774[(4'h8):(1'h0)]}));
                    end
                end
            end
          else
            begin
              if ((|(~reg772)))
                begin
                  for (forvar769 = (1'h0); (forvar769 < (2'h2)); forvar769 = (forvar769 + (1'h1)))
                    begin
                      reg770 <= wire741;
                      reg771 <= (((+$signed(reg757)) ?
                          ((wire741 ?
                              reg760 : reg750) || $signed(reg769)) : $signed((^wire741))) - (~((~forvar759) >> $unsigned(reg760))));
                    end
                  for (forvar772 = (1'h0); (forvar772 < (2'h3)); forvar772 = (forvar772 + (1'h1)))
                    begin
                      reg773 <= (|{((forvar753 ?
                              reg776 : reg775) ^~ forvar772[(4'h9):(3'h7)])});
                      reg774 <= $signed($unsigned(reg761));
                      reg775 <= (8'ha3);
                    end
                  if (forvar753)
                    begin
                      reg776 <= wire742[(4'h8):(3'h7)];
                      reg777 <= (8'hab);
                    end
                  else
                    begin
                      reg776 <= {({$unsigned(reg763)} == $signed((wire740 ?
                              (8'haf) : reg778)))};
                      reg777 <= (8'hb3);
                      reg778 <= (($unsigned($signed(wire740)) - $signed($unsigned(reg755))) * forvar747);
                      reg779 <= $unsigned((8'ha0));
                    end
                  if ($signed((-$unsigned({reg775}))))
                    begin
                      reg780 <= {$unsigned((reg771[(3'h7):(3'h4)] ?
                              $signed(reg751) : $signed((8'ha3))))};
                      reg781 <= $unsigned($signed({$unsigned(reg772)}));
                      reg782 <= reg772;
                    end
                  else
                    begin
                      reg780 <= ($signed(reg780[(3'h6):(1'h0)]) | reg770);
                    end
                end
              else
                begin
                  if ((^~(($signed((8'hb3)) | (reg773 ?
                      reg781 : reg776)) + {$signed(reg780)})))
                    begin
                      reg769 <= $signed((&((forvar758 ?
                          (8'ha7) : forvar762) & $signed((8'hb4)))));
                      reg770 <= $signed(($signed((~|reg752)) ?
                          forvar771 : reg772));
                    end
                  else
                    begin
                      reg769 <= $signed($signed(($signed(reg780) & {forvar771})));
                      reg770 <= reg749[(3'h4):(2'h2)];
                      reg771 <= ($signed((reg770[(3'h5):(3'h5)] ?
                              {reg779} : $signed(reg777))) ?
                          wire741 : $unsigned(forvar770[(1'h1):(1'h0)]));
                      reg772 <= ((reg752 || $unsigned($signed(forvar771))) ?
                          reg771 : ((&reg757) ~^ $unsigned(forvar759)));
                    end
                  reg773 <= $unsigned(($signed(((8'ha4) ?
                      reg765 : forvar758)) >> reg775[(1'h1):(1'h1)]));
                end
              if ((&(wire742 ?
                  ($unsigned(reg754) ?
                      forvar753 : (|reg777)) : ($unsigned((8'ha2)) * $signed((8'hb6))))))
                begin
                  for (forvar783 = (1'h0); (forvar783 < (2'h3)); forvar783 = (forvar783 + (1'h1)))
                    begin
                      reg784 <= reg761[(2'h2):(1'h1)];
                      reg785 <= $signed({$unsigned($signed(reg757))});
                      reg786 <= reg769;
                      reg787 <= (8'hab);
                    end
                  for (forvar788 = (1'h0); (forvar788 < (1'h1)); forvar788 = (forvar788 + (1'h1)))
                    begin
                      reg789 <= (|(|$signed((-reg775))));
                      reg790 <= ($signed($signed((~reg774))) ^ {(reg773 ?
                              wire743 : $unsigned(reg785))});
                      reg791 <= reg757;
                      reg792 <= reg785[(3'h5):(1'h1)];
                    end
                  reg793 <= ($signed(reg751[(4'hb):(2'h3)]) < (reg780 ^~ (^reg789)));
                  for (forvar794 = (1'h0); (forvar794 < (2'h2)); forvar794 = (forvar794 + (1'h1)))
                    begin
                      reg795 <= (~&(8'hac));
                      reg796 <= (((reg780 << {reg774}) ?
                          forvar758[(2'h3):(1'h1)] : $unsigned((forvar748 ?
                              (8'hb0) : wire741))) - $signed((forvar747 ?
                          reg772 : reg791[(4'hc):(3'h4)])));
                    end
                end
              else
                begin
                  if ((forvar766 != ($unsigned((forvar753 <<< (8'h9c))) <= $signed((wire740 >= reg770)))))
                    begin
                      reg783 <= forvar758;
                      reg784 <= $signed({forvar783[(2'h3):(2'h2)]});
                      reg785 <= $unsigned(($unsigned($signed(reg764)) ?
                          reg763[(3'h6):(1'h0)] : $unsigned((forvar770 * reg757))));
                      reg786 <= (^(((~^reg755) || $unsigned(wire745)) ^~ (~&(reg774 ?
                          forvar746 : reg779))));
                    end
                  else
                    begin
                      reg783 <= (($signed(reg763[(3'h4):(1'h0)]) ?
                              $signed($unsigned(reg771)) : (reg765 <<< ((8'hab) <<< reg792))) ?
                          {reg784[(1'h0):(1'h0)]} : (-(~{forvar794})));
                      reg784 <= $unsigned($signed((-(~^(8'hb3)))));
                      reg785 <= $signed(wire745);
                    end
                  if ((wire745[(1'h1):(1'h0)] ?
                      ((^$signed(forvar788)) >= {(reg776 ?
                              reg796 : reg792)}) : ((^~$unsigned(reg787)) | ((reg749 ?
                              reg790 : forvar771) ?
                          $unsigned(reg767) : reg772[(1'h0):(1'h0)]))))
                    begin
                      reg787 <= $signed({{reg792[(2'h2):(1'h1)]}});
                      reg788 <= reg778;
                      reg789 <= $signed((!wire741[(2'h2):(2'h2)]));
                      reg790 <= ((|(wire744 ?
                              (reg764 || reg761) : reg781[(3'h7):(2'h3)])) ?
                          (((+reg795) <<< reg776) && forvar771[(1'h1):(1'h0)]) : reg788[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg787 <= reg780[(2'h2):(1'h0)];
                      reg788 <= ((~^(+(!reg796))) << {(~&$unsigned(reg776))});
                    end
                  for (forvar791 = (1'h0); (forvar791 < (1'h1)); forvar791 = (forvar791 + (1'h1)))
                    begin
                      reg792 <= (^$signed({reg785}));
                      reg793 <= $signed($signed($signed((reg787 ?
                          (8'h9c) : wire742))));
                      reg794 <= $unsigned(({reg795[(2'h2):(1'h1)]} ?
                          $unsigned($unsigned(forvar759)) : reg795));
                    end
                end
              if ($signed(((reg774 ?
                  $unsigned(forvar769) : {forvar747}) & ((reg763 == (8'hb0)) != (reg767 + reg751)))))
                begin
                  reg797 <= (reg749 ?
                      $signed((|reg784)) : {(forvar759[(2'h2):(2'h2)] ^~ (reg768 ?
                              (8'ha4) : reg795))});
                  if ($signed((((reg782 + reg756) * (reg761 ?
                          reg793 : (8'ha0))) ?
                      $signed((forvar746 < reg750)) : $signed({(8'hab)}))))
                    begin
                      reg798 <= ({wire742[(3'h5):(1'h1)]} * wire741);
                      reg799 <= $signed(({$unsigned(reg752)} ?
                          (!((8'h9f) ? reg779 : reg770)) : {(forvar748 ?
                                  (8'hb5) : wire744)}));
                      reg800 <= ($unsigned(forvar788[(2'h2):(2'h2)]) ?
                          forvar772[(3'h4):(2'h2)] : $signed((((8'hb2) ?
                              reg761 : forvar794) ^~ reg777)));
                    end
                  else
                    begin
                      reg798 <= $unsigned((forvar788[(1'h1):(1'h1)] ?
                          forvar766 : (~^$unsigned(forvar746))));
                      reg799 <= $signed($unsigned(((-reg788) && $signed(reg792))));
                      reg800 <= (^~$unsigned(reg792));
                      reg801 <= (+reg781[(3'h6):(3'h6)]);
                    end
                end
              else
                begin
                  for (forvar797 = (1'h0); (forvar797 < (2'h2)); forvar797 = (forvar797 + (1'h1)))
                    begin
                      reg798 <= reg780[(3'h4):(2'h3)];
                      reg799 <= (|($unsigned(wire744) ?
                          (forvar771 ?
                              $unsigned(reg790) : (reg774 + reg760)) : {$unsigned(reg798)}));
                    end
                end
            end
          for (forvar802 = (1'h0); (forvar802 < (1'h1)); forvar802 = (forvar802 + (1'h1)))
            begin
              for (forvar803 = (1'h0); (forvar803 < (1'h1)); forvar803 = (forvar803 + (1'h1)))
                begin
                  reg804 <= $signed((forvar753[(3'h4):(3'h4)] <<< forvar794));
                  if (wire744)
                    begin
                      reg805 <= ($signed((8'h9c)) ?
                          forvar747[(4'ha):(3'h4)] : $signed((-reg755)));
                      reg806 <= reg771;
                    end
                  else
                    begin
                      reg805 <= reg792;
                      reg806 <= (|reg779);
                      reg807 <= ($signed(wire741) > (~^wire741[(4'h9):(1'h0)]));
                      reg808 <= $signed(reg779[(3'h5):(2'h3)]);
                    end
                  for (forvar809 = (1'h0); (forvar809 < (1'h1)); forvar809 = (forvar809 + (1'h1)))
                    begin
                      reg810 <= (((&$unsigned(reg796)) ?
                              reg771[(2'h3):(2'h2)] : (&$unsigned(forvar762))) ?
                          (reg749[(3'h5):(1'h0)] ^ (8'hb3)) : (!forvar794[(3'h6):(3'h4)]));
                    end
                  if ({$signed($signed(reg764[(3'h4):(2'h2)]))})
                    begin
                      reg811 <= {$unsigned((|(reg778 ~^ reg784)))};
                    end
                  else
                    begin
                      reg811 <= (8'hb1);
                    end
                end
              reg812 <= (^($signed((~|reg789)) ?
                  forvar746[(3'h6):(3'h4)] : $signed(reg751[(2'h3):(1'h1)])));
            end
        end
      for (forvar813 = (1'h0); (forvar813 < (2'h3)); forvar813 = (forvar813 + (1'h1)))
        begin
          for (forvar814 = (1'h0); (forvar814 < (2'h2)); forvar814 = (forvar814 + (1'h1)))
            begin
              for (forvar815 = (1'h0); (forvar815 < (1'h0)); forvar815 = (forvar815 + (1'h1)))
                begin
                  for (forvar816 = (1'h0); (forvar816 < (2'h2)); forvar816 = (forvar816 + (1'h1)))
                    begin
                      reg817 <= reg804;
                    end
                  if ($unsigned($unsigned(((+reg786) + (reg777 ?
                      (8'hb7) : reg751)))))
                    begin
                      reg818 <= ({reg752[(4'ha):(3'h5)]} ?
                          wire743 : forvar813[(1'h0):(1'h0)]);
                      reg819 <= (~^{((|reg781) && (reg779 ? reg764 : reg797))});
                      reg820 <= $unsigned(wire744[(4'h9):(4'h8)]);
                      reg821 <= (((-(forvar791 && reg776)) ?
                              {$signed(forvar802)} : ((8'hb1) ?
                                  $signed(forvar753) : $signed(reg819))) ?
                          $signed((!$unsigned(reg763))) : $signed((reg786[(3'h6):(3'h5)] ?
                              forvar753 : reg819[(2'h2):(2'h2)])));
                    end
                  else
                    begin
                      reg818 <= (~^forvar788[(2'h3):(2'h2)]);
                    end
                  reg822 <= reg781[(3'h4):(2'h2)];
                end
            end
          if (($signed($unsigned((forvar783 ? reg750 : wire742))) ?
              (^((&reg795) > (forvar797 | forvar762))) : {(reg764[(3'h4):(1'h0)] >> reg783)}))
            begin
              if ((|$signed((~^(forvar747 ? reg764 : reg780)))))
                begin
                  for (forvar823 = (1'h0); (forvar823 < (1'h1)); forvar823 = (forvar823 + (1'h1)))
                    begin
                      reg824 <= $signed(reg804[(2'h3):(2'h2)]);
                      reg825 <= $unsigned($signed((^(8'hb7))));
                    end
                  if ($signed((|(!$unsigned(reg781)))))
                    begin
                      reg826 <= {(+($signed(forvar797) ?
                              (reg750 >>> reg788) : reg799[(1'h0):(1'h0)]))};
                      reg827 <= (^((^(8'ha2)) | ($signed(forvar759) ?
                          $unsigned(reg822) : reg811)));
                    end
                  else
                    begin
                      reg826 <= ({$signed((reg796 == reg780))} ?
                          $signed(reg810[(4'ha):(4'ha)]) : ((forvar753[(2'h2):(1'h1)] < reg798) ?
                              {(reg801 == reg797)} : reg796));
                      reg827 <= $signed(({reg812} ?
                          (forvar797 ?
                              {reg827} : reg756[(4'h9):(1'h0)]) : $unsigned($signed(forvar809))));
                      reg828 <= (($signed($unsigned((8'hac))) ?
                          {(reg790 << (8'ha3))} : $signed(wire742[(4'h8):(4'h8)])) || forvar816);
                      reg829 <= $unsigned((forvar770[(3'h5):(2'h2)] << reg775));
                    end
                end
              else
                begin
                  reg823 <= ({reg806[(3'h5):(3'h5)]} ?
                      reg780 : (^~$unsigned((reg783 ? reg771 : reg795))));
                  if (reg805)
                    begin
                      reg824 <= forvar747;
                      reg825 <= (-(reg786[(2'h3):(1'h0)] ^ ((~&forvar747) & $unsigned(forvar814))));
                    end
                  else
                    begin
                      reg824 <= (^$signed((~^{reg772})));
                      reg825 <= ((~^reg768) & (8'hae));
                    end
                end
            end
          else
            begin
              for (forvar823 = (1'h0); (forvar823 < (1'h1)); forvar823 = (forvar823 + (1'h1)))
                begin
                  if ($signed(reg763[(2'h2):(2'h2)]))
                    begin
                      reg824 <= (8'hac);
                    end
                  else
                    begin
                      reg824 <= (|(($signed(reg768) ?
                          forvar794[(1'h1):(1'h0)] : (+reg754)) * {(^~(8'had))}));
                      reg825 <= ($signed($unsigned(reg810[(4'hb):(2'h3)])) << $unsigned(((|forvar815) ?
                          (forvar797 ^~ forvar770) : reg820)));
                    end
                end
              if (forvar759[(3'h4):(3'h4)])
                begin
                  if ($signed({$signed((reg828 > reg812))}))
                    begin
                      reg826 <= (8'hb7);
                      reg827 <= $signed({$unsigned((forvar783 ?
                              forvar794 : (8'hba)))});
                    end
                  else
                    begin
                      reg826 <= reg781;
                      reg827 <= (({{(8'hab)}} - reg771[(3'h5):(3'h4)]) ?
                          $signed(($signed(reg778) >> (reg781 ?
                              forvar772 : reg781))) : $unsigned($signed((reg783 ?
                              reg792 : (8'hb5)))));
                    end
                end
              else
                begin
                  if ($unsigned((-reg798[(1'h1):(1'h1)])))
                    begin
                      reg826 <= (&(^~reg779[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg826 <= forvar771;
                      reg827 <= forvar797[(1'h1):(1'h1)];
                      reg828 <= (~^$unsigned(($signed(reg789) ^~ forvar791[(2'h2):(1'h0)])));
                      reg829 <= (8'hba);
                    end
                end
              for (forvar830 = (1'h0); (forvar830 < (2'h2)); forvar830 = (forvar830 + (1'h1)))
                begin
                  for (forvar831 = (1'h0); (forvar831 < (2'h3)); forvar831 = (forvar831 + (1'h1)))
                    begin
                      reg832 <= ($signed((reg812[(3'h6):(1'h1)] >> ((8'ha2) == reg752))) ?
                          (~|(!(|reg785))) : (forvar823 ?
                              (reg810[(3'h4):(2'h3)] ?
                                  reg796 : (forvar830 >>> reg751)) : (forvar814 ?
                                  $unsigned(reg752) : {reg795})));
                      reg833 <= $unsigned(((reg764 ^~ $signed((8'hb1))) ?
                          ($signed(reg797) | $unsigned(reg796)) : $unsigned(((8'hb5) ?
                              reg793 : reg769))));
                    end
                end
              for (forvar834 = (1'h0); (forvar834 < (2'h3)); forvar834 = (forvar834 + (1'h1)))
                begin
                  reg835 <= wire740[(1'h0):(1'h0)];
                end
            end
          reg836 <= {(~&$signed($signed(reg777)))};
        end
      reg837 <= ((|$unsigned((reg807 ?
          reg787 : (8'had)))) >>> reg817[(3'h5):(3'h4)]);
    end
  assign wire838 = reg750;
  always
    @(posedge clk) begin
      for (forvar839 = (1'h0); (forvar839 < (1'h0)); forvar839 = (forvar839 + (1'h1)))
        begin
          reg840 <= ($signed(($signed(reg788) ~^ ((8'h9f) <<< reg836))) ?
              {$signed((wire743 ?
                      reg757 : (8'h9f)))} : $unsigned($signed((reg799 ?
                  reg782 : (8'hb1)))));
        end
      for (forvar841 = (1'h0); (forvar841 < (2'h2)); forvar841 = (forvar841 + (1'h1)))
        begin
          for (forvar842 = (1'h0); (forvar842 < (2'h2)); forvar842 = (forvar842 + (1'h1)))
            begin
              if (reg765)
                begin
                  for (forvar843 = (1'h0); (forvar843 < (1'h1)); forvar843 = (forvar843 + (1'h1)))
                    begin
                      reg844 <= ($unsigned((-(^reg764))) ?
                          (reg808 ?
                              $signed({reg832}) : reg767) : $unsigned({(-reg764)}));
                    end
                  for (forvar845 = (1'h0); (forvar845 < (1'h0)); forvar845 = (forvar845 + (1'h1)))
                    begin
                      reg846 <= ($signed({(reg761 ?
                              reg750 : forvar843)}) >= $signed((reg761[(2'h2):(2'h2)] ?
                          ((8'ha3) == reg768) : forvar841[(1'h0):(1'h0)])));
                      reg847 <= $signed($signed(reg769));
                      reg848 <= (|$signed(reg773));
                      reg849 <= ($signed((|(reg772 ?
                          reg828 : reg812))) >>> (((8'h9f) >>> $signed(reg783)) <= $unsigned(forvar843[(1'h1):(1'h0)])));
                    end
                  for (forvar850 = (1'h0); (forvar850 < (1'h1)); forvar850 = (forvar850 + (1'h1)))
                    begin
                      reg851 <= (reg777[(2'h2):(2'h2)] ? reg756 : reg833);
                      reg852 <= (8'hb8);
                      reg853 <= ((~(reg794[(3'h6):(3'h6)] ?
                              ((8'ha3) ?
                                  forvar841 : reg820) : $unsigned(reg833))) ?
                          reg817 : (reg780[(2'h3):(1'h0)] ?
                              ((reg783 ?
                                  reg778 : (8'ha1)) || reg820[(3'h4):(1'h0)]) : (reg824 ?
                                  (~&wire741) : $unsigned(reg776))));
                    end
                end
              else
                begin
                  for (forvar843 = (1'h0); (forvar843 < (1'h0)); forvar843 = (forvar843 + (1'h1)))
                    begin
                      reg844 <= ($signed($unsigned(reg756[(4'ha):(4'h8)])) - {reg829});
                      reg845 <= reg844;
                      reg846 <= ((~(~&(reg833 ? reg770 : reg800))) ?
                          reg822 : {((reg846 ? reg771 : reg764) ?
                                  reg779 : ((8'hb8) + (8'h9d)))});
                    end
                  if ((-($unsigned((reg849 ?
                      reg768 : reg793)) * reg769[(2'h3):(1'h1)])))
                    begin
                      reg847 <= ((8'ha7) != $signed(reg752[(4'h8):(1'h1)]));
                      reg848 <= (reg788 >>> (forvar843[(2'h3):(1'h1)] ?
                          $signed($signed(reg768)) : (((8'ha1) ?
                                  reg778 : reg825) ?
                              $unsigned(reg829) : (!reg760))));
                    end
                  else
                    begin
                      reg847 <= $signed((8'ha7));
                      reg848 <= forvar845;
                      reg849 <= (forvar841[(3'h7):(2'h3)] ?
                          (reg822[(2'h2):(2'h2)] ?
                              $unsigned((wire743 ?
                                  reg847 : reg757)) : $unsigned($signed(reg772))) : (8'haf));
                      reg850 <= (+reg800[(4'hb):(3'h7)]);
                    end
                  for (forvar851 = (1'h0); (forvar851 < (1'h1)); forvar851 = (forvar851 + (1'h1)))
                    begin
                      reg852 <= $signed(($signed((reg823 ?
                          reg845 : forvar841)) <= $unsigned((reg754 ?
                          reg761 : reg782))));
                      reg853 <= ((+((~reg778) ?
                          reg806 : reg837[(4'hb):(2'h3)])) >= (reg750 ?
                          ({(8'hb8)} ^ {reg808}) : $unsigned(wire744)));
                      reg854 <= $unsigned($unsigned((reg780 ?
                          $unsigned(reg761) : $unsigned(reg799))));
                      reg855 <= forvar842;
                    end
                end
            end
          if ((~^(((reg787 ? reg767 : forvar845) << reg782) - forvar842)))
            begin
              if (reg751)
                begin
                  for (forvar856 = (1'h0); (forvar856 < (2'h3)); forvar856 = (forvar856 + (1'h1)))
                    begin
                      reg857 <= ($unsigned({{(8'hb2)}}) == $unsigned(reg773));
                      reg858 <= (8'ha5);
                      reg859 <= $unsigned($unsigned((~|(reg819 + reg791))));
                      reg860 <= {$unsigned((wire741[(4'h9):(1'h0)] ?
                              ((8'hb6) ? reg785 : reg859) : (+reg789)))};
                    end
                  reg861 <= reg789[(3'h4):(1'h1)];
                  for (forvar862 = (1'h0); (forvar862 < (2'h3)); forvar862 = (forvar862 + (1'h1)))
                    begin
                      reg863 <= $unsigned(reg827[(3'h6):(1'h1)]);
                      reg864 <= reg820;
                    end
                end
              else
                begin
                  for (forvar856 = (1'h0); (forvar856 < (2'h3)); forvar856 = (forvar856 + (1'h1)))
                    begin
                      reg857 <= $unsigned($unsigned($signed($unsigned(wire743))));
                    end
                  reg858 <= (~(~(reg749[(1'h0):(1'h0)] >= (8'h9e))));
                  reg859 <= (~&reg785[(1'h0):(1'h0)]);
                  reg860 <= ({((wire741 == reg811) ?
                              reg751[(2'h3):(1'h1)] : (reg851 ?
                                  (8'hb4) : wire838))} ?
                      $signed((^reg805[(3'h4):(2'h3)])) : (!reg780));
                end
              if ((^~reg826))
                begin
                  for (forvar865 = (1'h0); (forvar865 < (2'h3)); forvar865 = (forvar865 + (1'h1)))
                    begin
                      reg866 <= forvar862[(1'h0):(1'h0)];
                      reg867 <= $unsigned((($unsigned(reg808) ?
                          $signed(reg799) : $unsigned(reg844)) + ($signed(reg861) ?
                          reg793 : forvar865)));
                      reg868 <= ($unsigned((reg844 ?
                              $signed(reg776) : {reg837})) ?
                          {reg795[(3'h4):(2'h3)]} : $signed(forvar850[(3'h6):(2'h3)]));
                    end
                  if ((&(8'ha5)))
                    begin
                      reg869 <= reg772;
                      reg870 <= ((~&(((8'ha1) >= reg786) ?
                          {reg750} : $unsigned(reg836))) ^~ reg868);
                      reg871 <= (^wire740);
                    end
                  else
                    begin
                      reg869 <= $unsigned({(~&(~^reg781))});
                      reg870 <= ($unsigned((reg851[(1'h0):(1'h0)] ?
                              (8'hb4) : reg797[(1'h1):(1'h0)])) ?
                          reg794[(4'he):(4'he)] : (&reg789));
                    end
                end
              else
                begin
                  if (((((wire740 ? (8'hb9) : reg868) <<< $signed(reg860)) ?
                      {$signed(reg836)} : ($signed(reg858) - (^(8'ha0)))) + ($signed(reg764[(2'h3):(1'h1)]) ?
                      ((~|(8'hb4)) ?
                          (forvar851 ?
                              reg811 : reg812) : $unsigned((8'ha7))) : $unsigned({(8'hb3)}))))
                    begin
                      reg865 <= ($unsigned(((+(8'ha2)) != reg812[(2'h3):(1'h1)])) ~^ $unsigned((|(reg793 < reg784))));
                      reg866 <= $unsigned(reg765);
                      reg867 <= ((-({forvar845} != (reg820 ?
                          reg832 : forvar839))) + reg751[(3'h7):(2'h3)]);
                      reg868 <= $unsigned((forvar845 >= forvar862));
                    end
                  else
                    begin
                      reg865 <= {(^(^(wire741 - reg868)))};
                      reg866 <= (reg800[(4'ha):(3'h7)] == (~((reg852 ?
                              reg819 : reg808) ?
                          reg798[(3'h4):(1'h0)] : (8'hb7))));
                      reg867 <= {($unsigned(((8'ha6) || (8'hae))) & reg861[(1'h0):(1'h0)])};
                      reg868 <= (($signed({wire838}) || wire742) ?
                          reg828 : $unsigned(wire742[(2'h3):(2'h2)]));
                    end
                  if ((&reg781[(1'h0):(1'h0)]))
                    begin
                      reg869 <= $signed(($unsigned(forvar856[(3'h4):(2'h3)]) ?
                          (!(reg857 ?
                              reg751 : reg865)) : (+reg819[(1'h1):(1'h0)])));
                      reg870 <= (wire743[(1'h1):(1'h0)] ^ (reg784[(3'h5):(1'h1)] ?
                          $unsigned(reg844) : $unsigned({reg787})));
                    end
                  else
                    begin
                      reg869 <= {$unsigned(((reg817 ? reg848 : forvar839) ?
                              {reg780} : $signed(reg798)))};
                      reg870 <= (~^(8'ha8));
                      reg871 <= $signed(({(|reg860)} + $signed(forvar841)));
                    end
                  for (forvar872 = (1'h0); (forvar872 < (1'h0)); forvar872 = (forvar872 + (1'h1)))
                    begin
                      reg873 <= ({reg804[(2'h3):(2'h2)]} | $unsigned($signed($signed((8'hb6)))));
                    end
                  reg874 <= {reg774[(4'h9):(1'h0)]};
                end
              for (forvar875 = (1'h0); (forvar875 < (2'h2)); forvar875 = (forvar875 + (1'h1)))
                begin
                  if ({reg851[(2'h3):(1'h0)]})
                    begin
                      reg876 <= ((^~$unsigned(((8'hac) ?
                          wire745 : reg795))) | $unsigned((&(reg808 >= reg771))));
                      reg877 <= reg845;
                      reg878 <= (~$unsigned($signed($signed((8'hb0)))));
                    end
                  else
                    begin
                      reg876 <= reg835[(2'h2):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar856 = (1'h0); (forvar856 < (2'h3)); forvar856 = (forvar856 + (1'h1)))
                begin
                  for (forvar857 = (1'h0); (forvar857 < (2'h2)); forvar857 = (forvar857 + (1'h1)))
                    begin
                      reg858 <= ({$signed(reg795)} ?
                          reg773 : (~|$signed((reg836 ? reg873 : wire744))));
                      reg859 <= ((((~^reg770) ? (!reg810) : $signed((8'hb6))) ?
                              ((reg771 < forvar875) ?
                                  (reg808 ?
                                      wire745 : reg789) : (^~reg795)) : ((&forvar872) - forvar857[(3'h4):(2'h3)])) ?
                          (|((reg819 || reg774) ?
                              reg764 : (reg796 <<< (8'h9e)))) : $signed(($unsigned(reg796) ?
                              (^~forvar872) : reg769[(3'h4):(3'h4)])));
                    end
                end
              if (reg804[(2'h3):(2'h3)])
                begin
                  if ((((^~(8'hac)) ? $signed((^reg829)) : forvar851) ?
                      (($signed(reg768) ?
                          ((8'ha6) < forvar843) : (reg851 >= reg781)) + (!(8'hb5))) : $unsigned(($signed(reg779) ?
                          (wire743 ?
                              (8'h9c) : reg790) : $unsigned(forvar865)))))
                    begin
                      reg860 <= (~($signed((+reg874)) <<< {$unsigned(reg853)}));
                      reg861 <= reg851[(1'h1):(1'h0)];
                      reg862 <= $unsigned(forvar841[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg860 <= reg837;
                    end
                  for (forvar863 = (1'h0); (forvar863 < (2'h3)); forvar863 = (forvar863 + (1'h1)))
                    begin
                      reg864 <= $signed($unsigned($unsigned($unsigned(forvar841))));
                      reg865 <= reg847[(2'h3):(2'h3)];
                      reg866 <= $signed((&((reg783 ?
                          (8'ha4) : wire740) < $signed(reg853))));
                    end
                  if ({reg864})
                    begin
                      reg867 <= reg756[(3'h4):(2'h3)];
                      reg868 <= reg785;
                      reg869 <= ({((forvar875 >> (8'hb5)) + (~&reg764))} ?
                          ({(reg789 <= reg757)} - (!reg761)) : ($unsigned($signed(reg779)) <= $unsigned(reg819)));
                      reg870 <= (!$unsigned($unsigned($unsigned((8'ha2)))));
                    end
                  else
                    begin
                      reg867 <= $unsigned((reg760 < ((!reg812) | {reg820})));
                      reg868 <= (!(~^(~(+reg819))));
                    end
                  if ((~reg833[(2'h2):(2'h2)]))
                    begin
                      reg871 <= (({(reg833 ?
                              reg836 : reg811)} ^ reg865[(1'h0):(1'h0)]) - $unsigned(reg846));
                      reg872 <= (8'haa);
                    end
                  else
                    begin
                      reg871 <= $signed($signed(((8'haf) ?
                          (reg823 >> reg861) : $signed(forvar856))));
                      reg872 <= ((reg780 >= reg865) & $unsigned($unsigned((reg772 | reg832))));
                      reg873 <= ((reg770 ?
                          ($unsigned(wire742) >= ((8'hb8) ?
                              reg857 : (8'hb4))) : {$unsigned(reg855)}) ~^ ($unsigned($unsigned(reg787)) ?
                          reg822 : $unsigned((reg781 ? (8'haf) : reg765))));
                    end
                end
              else
                begin
                  for (forvar860 = (1'h0); (forvar860 < (1'h1)); forvar860 = (forvar860 + (1'h1)))
                    begin
                      reg861 <= $signed((^reg763));
                      reg862 <= reg807[(3'h7):(3'h7)];
                      reg863 <= reg790;
                      reg864 <= $signed((reg859 != reg876));
                    end
                  for (forvar865 = (1'h0); (forvar865 < (1'h0)); forvar865 = (forvar865 + (1'h1)))
                    begin
                      reg866 <= (({$signed((8'ha2))} ?
                          ($signed(reg786) > {reg825}) : (+{reg775})) > {reg824});
                      reg867 <= (^~((^~reg781[(3'h4):(1'h0)]) == $signed($signed(reg868))));
                      reg868 <= reg774;
                      reg869 <= $signed((8'ha3));
                    end
                  if (reg775[(2'h3):(2'h3)])
                    begin
                      reg870 <= (8'ha6);
                      reg871 <= {((~reg761[(1'h0):(1'h0)]) ?
                              (~|$unsigned(reg837)) : (reg794 ?
                                  {reg835} : (&(8'ha4))))};
                      reg872 <= (!reg867[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg870 <= reg757;
                    end
                end
              for (forvar874 = (1'h0); (forvar874 < (2'h2)); forvar874 = (forvar874 + (1'h1)))
                begin
                  if (reg794)
                    begin
                      reg875 <= (forvar850 ? reg837[(4'h8):(1'h1)] : wire740);
                      reg876 <= ($signed((~^$signed(reg764))) ?
                          (reg794 ?
                              $unsigned((~|reg780)) : $signed($unsigned(reg801))) : reg760);
                      reg877 <= (^($unsigned(reg749[(1'h0):(1'h0)]) ?
                          ($signed(reg787) ?
                              reg869 : reg858) : {$unsigned(reg829)}));
                      reg878 <= ($unsigned(reg851) ~^ reg846[(4'hc):(1'h1)]);
                    end
                  else
                    begin
                      reg875 <= reg770[(4'h8):(3'h5)];
                      reg876 <= (~|(!reg872));
                    end
                  for (forvar879 = (1'h0); (forvar879 < (2'h3)); forvar879 = (forvar879 + (1'h1)))
                    begin
                      reg880 <= $signed(reg829);
                      reg881 <= ((~(-(reg793 ?
                          reg846 : (8'ha3)))) >= ($signed($unsigned(reg820)) > (reg755[(3'h4):(2'h3)] ?
                          (reg806 ? (8'hb3) : wire742) : {reg756})));
                      reg882 <= reg828[(3'h4):(1'h1)];
                    end
                  if (reg792)
                    begin
                      reg883 <= ((reg782[(2'h2):(1'h0)] == $signed((reg847 >= reg861))) ?
                          (((&forvar843) ~^ $unsigned(reg866)) ?
                              {reg763[(2'h2):(1'h0)]} : $signed((!(8'h9e)))) : ((reg826 ?
                                  {reg788} : reg871) ?
                              (-$signed(reg801)) : forvar874));
                      reg884 <= $unsigned($unsigned((reg805[(3'h6):(2'h3)] ?
                          reg878 : $unsigned(reg863))));
                    end
                  else
                    begin
                      reg883 <= $signed(forvar862[(2'h2):(1'h1)]);
                      reg884 <= reg871;
                    end
                  reg885 <= $signed(reg873[(1'h1):(1'h0)]);
                end
            end
          if ((|$signed((-(~&forvar841)))))
            begin
              reg886 <= {(({reg873} ?
                      $unsigned(reg767) : (reg799 ?
                          reg767 : reg782)) ^ (8'hb1))};
            end
          else
            begin
              reg886 <= reg829[(4'ha):(2'h3)];
            end
          for (forvar887 = (1'h0); (forvar887 < (1'h0)); forvar887 = (forvar887 + (1'h1)))
            begin
              if ($signed(($signed({reg824}) >>> $signed(reg829))))
                begin
                  for (forvar888 = (1'h0); (forvar888 < (2'h2)); forvar888 = (forvar888 + (1'h1)))
                    begin
                      reg889 <= (+$signed(({forvar850} + $unsigned(wire740))));
                      reg890 <= reg850;
                      reg891 <= $unsigned((&$signed((!reg777))));
                    end
                  if (reg863[(1'h0):(1'h0)])
                    begin
                      reg892 <= (!(-$signed((reg787 - (8'hb9)))));
                      reg893 <= {(reg772[(3'h4):(2'h2)] > reg754[(1'h1):(1'h0)])};
                      reg894 <= ($signed(reg794) > (|(^(~&reg778))));
                    end
                  else
                    begin
                      reg892 <= reg771;
                      reg893 <= $signed((($unsigned(reg890) ~^ $unsigned(reg819)) ?
                          (8'hb6) : (((8'ha2) ? reg770 : forvar850) ?
                              (reg812 ? reg781 : reg769) : $unsigned(reg885))));
                      reg894 <= $unsigned(((reg756[(3'h4):(1'h1)] || $signed(wire741)) ?
                          (reg881[(1'h0):(1'h0)] ?
                              $unsigned((8'hb0)) : reg763[(1'h1):(1'h1)]) : (&$signed(reg773))));
                      reg895 <= reg763[(2'h3):(1'h0)];
                    end
                  if (($signed($signed($unsigned(reg810))) ?
                      ((!reg826) < {reg800}) : $signed($unsigned(forvar874))))
                    begin
                      reg896 <= ((~{(reg871 == forvar842)}) >> forvar857);
                      reg897 <= $signed(($signed($signed(reg874)) ?
                          reg793 : $unsigned((-(8'ha8)))));
                      reg898 <= reg789[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg896 <= reg820;
                      reg897 <= ((~|{$signed(reg897)}) ?
                          $signed(reg866) : $unsigned(wire742));
                    end
                  for (forvar899 = (1'h0); (forvar899 < (2'h2)); forvar899 = (forvar899 + (1'h1)))
                    begin
                      reg900 <= wire743;
                      reg901 <= $signed({reg866[(2'h2):(1'h1)]});
                    end
                end
              else
                begin
                  reg888 <= $unsigned((~|(!(~&reg820))));
                  for (forvar889 = (1'h0); (forvar889 < (2'h2)); forvar889 = (forvar889 + (1'h1)))
                    begin
                      reg890 <= ($signed($unsigned((reg785 ?
                              reg875 : reg819))) ?
                          $signed($signed({forvar857})) : $signed(((reg804 ?
                                  (8'ha4) : forvar839) ?
                              (forvar863 ?
                                  (8'hab) : reg782) : forvar865[(3'h5):(3'h4)])));
                      reg891 <= (&{reg837});
                      reg892 <= reg860[(1'h0):(1'h0)];
                      reg893 <= (8'hb3);
                    end
                end
              for (forvar902 = (1'h0); (forvar902 < (2'h2)); forvar902 = (forvar902 + (1'h1)))
                begin
                  for (forvar903 = (1'h0); (forvar903 < (2'h3)); forvar903 = (forvar903 + (1'h1)))
                    begin
                      reg904 <= ($unsigned(((reg760 ?
                              reg872 : reg763) || reg760[(4'h8):(1'h1)])) ?
                          forvar875 : (($unsigned(reg865) != reg761[(2'h2):(1'h1)]) ?
                              ($signed(reg806) - (-reg864)) : $signed($signed((8'ha7)))));
                      reg905 <= reg889[(1'h0):(1'h0)];
                      reg906 <= ((8'ha3) > (((reg901 & reg846) >>> reg851) ?
                          reg794 : reg844[(3'h7):(3'h6)]));
                    end
                end
              if ($signed((reg873 ^~ reg840)))
                begin
                  for (forvar907 = (1'h0); (forvar907 < (2'h3)); forvar907 = (forvar907 + (1'h1)))
                    begin
                      reg908 <= reg854;
                      reg909 <= forvar888[(2'h3):(2'h2)];
                    end
                  for (forvar910 = (1'h0); (forvar910 < (1'h1)); forvar910 = (forvar910 + (1'h1)))
                    begin
                      reg911 <= ($unsigned(($unsigned((8'hb9)) ?
                              (reg857 >>> reg881) : {reg807})) ?
                          (8'hb3) : ($unsigned(reg845[(4'ha):(4'ha)]) <= $unsigned($unsigned(reg900))));
                      reg912 <= ((reg778 ? forvar850 : $signed((~^reg792))) ?
                          reg770[(4'ha):(4'ha)] : reg755[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  if ((reg778[(1'h0):(1'h0)] < reg826[(1'h1):(1'h1)]))
                    begin
                      reg907 <= $unsigned(reg872[(3'h5):(3'h4)]);
                      reg908 <= (((reg769 ? (&reg911) : (~reg845)) ?
                              ($signed((8'hae)) >> (reg874 | wire744)) : (|reg818[(4'ha):(4'h8)])) ?
                          $unsigned((reg786[(4'hc):(4'h9)] ?
                              reg764[(4'ha):(4'h9)] : $signed(reg787))) : (^~$unsigned(forvar887)));
                      reg909 <= (8'had);
                      reg910 <= reg852;
                    end
                  else
                    begin
                      reg907 <= ({(~&(reg828 >> forvar843))} ?
                          $unsigned((|reg861[(1'h0):(1'h0)])) : (reg769 ?
                              $signed((reg865 ?
                                  (8'ha6) : reg863)) : $signed(reg820[(2'h3):(1'h1)])));
                      reg908 <= $unsigned((^~$unsigned((forvar839 ?
                          reg801 : (8'hba)))));
                    end
                end
              if (reg885[(1'h0):(1'h0)])
                begin
                  if (({$signed($signed(reg876))} >>> forvar851))
                    begin
                      reg913 <= reg765[(4'he):(4'h8)];
                      reg914 <= ($signed($signed(reg788[(3'h6):(3'h6)])) ?
                          {((~^reg764) ^ $unsigned(reg835))} : $unsigned(reg794));
                      reg915 <= reg854;
                      reg916 <= (8'hae);
                    end
                  else
                    begin
                      reg913 <= {(((~^(8'ha7)) * $unsigned(reg770)) << ((reg780 ^ reg827) ?
                              reg780 : $unsigned(reg863)))};
                      reg914 <= reg775[(3'h6):(3'h5)];
                    end
                  if ($signed(reg896[(3'h6):(1'h0)]))
                    begin
                      reg917 <= (($signed($unsigned(reg908)) & (~&forvar851[(2'h3):(2'h3)])) ?
                          reg829[(1'h1):(1'h1)] : (^~((|reg807) >= (+reg872))));
                      reg918 <= (|((&$signed(reg844)) >> ((!reg788) ?
                          {(8'ha2)} : wire741[(4'h8):(2'h3)])));
                      reg919 <= $unsigned(reg789);
                    end
                  else
                    begin
                      reg917 <= reg872[(4'ha):(3'h7)];
                      reg918 <= $signed((~^$signed({reg837})));
                      reg919 <= (($unsigned(reg819) >= ($signed(reg871) ?
                          (|(8'ha7)) : reg892)) << reg791[(4'ha):(1'h0)]);
                    end
                  for (forvar920 = (1'h0); (forvar920 < (1'h1)); forvar920 = (forvar920 + (1'h1)))
                    begin
                      reg921 <= $signed(reg819[(1'h1):(1'h0)]);
                      reg922 <= ((!$unsigned((!reg799))) && $signed(reg859));
                      reg923 <= forvar907[(3'h6):(1'h1)];
                    end
                end
              else
                begin
                  if ($unsigned((&($unsigned((8'hb4)) ?
                      $unsigned(reg828) : {reg890}))))
                    begin
                      reg913 <= (!reg884);
                      reg914 <= $signed((-(reg890[(2'h2):(2'h2)] - $unsigned(forvar842))));
                      reg915 <= $signed((((reg849 ?
                              reg870 : forvar857) >= (forvar841 ?
                              reg859 : reg828)) ?
                          $unsigned((reg773 ^ reg847)) : (8'ha3)));
                      reg916 <= (($signed((^~reg889)) ?
                              reg820 : wire743[(1'h1):(1'h1)]) ?
                          reg836[(2'h3):(1'h1)] : ($unsigned((reg898 ?
                                  reg829 : reg891)) ?
                              forvar899 : $unsigned(reg767)));
                    end
                  else
                    begin
                      reg913 <= ((((reg863 ?
                              (8'hb4) : reg870) * $unsigned(reg808)) ?
                          (reg771[(1'h0):(1'h0)] + (-forvar920)) : ((reg756 ?
                                  reg848 : (8'hb7)) ?
                              (~&reg866) : {reg866})) >> (~^$signed((8'hba))));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed(reg800))
        begin
          for (forvar924 = (1'h0); (forvar924 < (1'h0)); forvar924 = (forvar924 + (1'h1)))
            begin
              reg925 <= reg861[(1'h1):(1'h0)];
              if (reg760[(4'h9):(3'h6)])
                begin
                  if ((reg799 | (~|(((8'hb6) ? reg784 : reg895) ?
                      $unsigned((8'haf)) : $signed(reg801)))))
                    begin
                      reg926 <= reg906[(2'h3):(1'h0)];
                      reg927 <= (({reg892[(4'h8):(1'h0)]} == reg765) ?
                          reg913[(3'h7):(2'h3)] : ({((8'hb7) ?
                                  wire744 : reg773)} & (-reg862)));
                      reg928 <= (((^$signed(reg890)) ?
                              reg793[(1'h0):(1'h0)] : (~(&reg847))) ?
                          (!{reg774[(4'h8):(2'h3)]}) : $signed((reg804 * $unsigned((8'h9e)))));
                    end
                  else
                    begin
                      reg926 <= (reg925[(2'h3):(2'h3)] < ((&$unsigned((8'hb9))) >>> ({(8'hb6)} + wire838)));
                      reg927 <= $signed(reg865);
                      reg928 <= $signed($signed(reg811[(4'he):(1'h1)]));
                      reg929 <= reg917;
                    end
                end
              else
                begin
                  for (forvar926 = (1'h0); (forvar926 < (2'h2)); forvar926 = (forvar926 + (1'h1)))
                    begin
                      reg927 <= $signed(reg923);
                    end
                  for (forvar928 = (1'h0); (forvar928 < (1'h1)); forvar928 = (forvar928 + (1'h1)))
                    begin
                      reg929 <= (!(({reg757} ?
                              ((8'hba) ?
                                  reg878 : reg817) : (reg818 || reg889)) ?
                          $unsigned({reg890}) : $unsigned($signed(reg891))));
                      reg930 <= $unsigned({{$unsigned(reg901)}});
                      reg931 <= reg893;
                      reg932 <= {reg774[(1'h0):(1'h0)]};
                    end
                end
              for (forvar933 = (1'h0); (forvar933 < (1'h1)); forvar933 = (forvar933 + (1'h1)))
                begin
                  reg934 <= $signed($signed(reg751[(3'h7):(1'h1)]));
                  if (((((-reg768) ? $signed(reg922) : reg817) ^ (|(reg873 ?
                          reg805 : (8'ha1)))) ?
                      $signed((+$signed(reg921))) : (reg930[(3'h6):(2'h3)] ?
                          $unsigned((reg892 ? (8'ha5) : (8'hb9))) : reg863)))
                    begin
                      reg935 <= (~$signed(reg781));
                    end
                  else
                    begin
                      reg935 <= ($unsigned($signed(reg909)) ?
                          (~((!reg820) ?
                              (^reg862) : (forvar933 ?
                                  reg905 : (8'ha6)))) : (((~&reg935) * (&(8'h9d))) >>> {(~&reg873)}));
                      reg936 <= ((^~reg897[(3'h5):(1'h0)]) ?
                          reg859[(2'h3):(1'h0)] : ($unsigned($unsigned(reg850)) & ($unsigned(reg847) ?
                              (reg932 ?
                                  reg869 : (8'ha8)) : $unsigned(reg799))));
                    end
                  reg937 <= ($unsigned((+reg853[(2'h3):(1'h0)])) ?
                      reg892 : (8'haf));
                end
              reg938 <= (reg804[(3'h4):(1'h1)] ?
                  ($signed(((8'hb4) >>> reg849)) > reg851[(3'h4):(3'h4)]) : (((^~(8'hab)) >>> $signed((8'h9d))) >>> (reg929 >= forvar924[(2'h2):(1'h0)])));
            end
        end
      else
        begin
          for (forvar924 = (1'h0); (forvar924 < (2'h2)); forvar924 = (forvar924 + (1'h1)))
            begin
              for (forvar925 = (1'h0); (forvar925 < (2'h3)); forvar925 = (forvar925 + (1'h1)))
                begin
                  for (forvar926 = (1'h0); (forvar926 < (1'h0)); forvar926 = (forvar926 + (1'h1)))
                    begin
                      reg927 <= {$signed(wire838[(1'h0):(1'h0)])};
                    end
                  for (forvar928 = (1'h0); (forvar928 < (1'h0)); forvar928 = (forvar928 + (1'h1)))
                    begin
                      reg929 <= reg806;
                      reg930 <= (reg912 ?
                          (&reg796) : ($signed((|reg932)) ?
                              (((8'ha7) ^~ reg768) <= reg811) : {$unsigned(reg797)}));
                      reg931 <= ((reg927 ?
                              reg852[(3'h7):(1'h1)] : ((-reg891) ?
                                  reg935 : reg884)) ?
                          {(^$signed(reg775))} : (!(reg789 ~^ reg872[(1'h0):(1'h0)])));
                      reg932 <= ($unsigned((^(!(8'hb1)))) ?
                          (($unsigned((8'ha5)) >> (reg751 ? (8'hb6) : reg775)) ?
                              reg761 : reg845) : reg912);
                    end
                end
            end
          for (forvar933 = (1'h0); (forvar933 < (1'h0)); forvar933 = (forvar933 + (1'h1)))
            begin
              if ($signed($unsigned(($signed(reg807) >> $signed(reg870)))))
                begin
                  if (reg861[(2'h2):(2'h2)])
                    begin
                      reg934 <= ($signed((~^{reg788})) ?
                          reg886 : (^~{$unsigned(reg752)}));
                      reg935 <= ((8'hb3) ?
                          $unsigned((8'h9f)) : reg919[(4'h9):(3'h4)]);
                      reg936 <= reg812;
                      reg937 <= forvar933[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg934 <= wire742;
                      reg935 <= ($unsigned({$signed(reg811)}) ?
                          (($signed((8'hb8)) - (reg819 ^~ (8'hb0))) * reg787) : (reg767 ?
                              ($unsigned(reg910) >>> reg894) : ((reg885 > (8'ha5)) ?
                                  ((8'ha2) ?
                                      reg937 : reg799) : reg897[(1'h0):(1'h0)])));
                      reg936 <= ($unsigned(reg774) - (8'hb1));
                    end
                  for (forvar938 = (1'h0); (forvar938 < (2'h2)); forvar938 = (forvar938 + (1'h1)))
                    begin
                      reg939 <= $signed($unsigned((~&reg875)));
                      reg940 <= $unsigned($signed((~|$signed((8'hb1)))));
                    end
                end
              else
                begin
                  reg934 <= reg897[(3'h6):(1'h0)];
                  reg935 <= reg888;
                end
            end
        end
      if ((((|(reg861 > reg867)) >= ((forvar928 >> reg894) >>> $unsigned((8'hb5)))) - $unsigned($unsigned((&reg825)))))
        begin
          for (forvar941 = (1'h0); (forvar941 < (2'h3)); forvar941 = (forvar941 + (1'h1)))
            begin
              for (forvar942 = (1'h0); (forvar942 < (2'h2)); forvar942 = (forvar942 + (1'h1)))
                begin
                  for (forvar943 = (1'h0); (forvar943 < (2'h3)); forvar943 = (forvar943 + (1'h1)))
                    begin
                      reg944 <= {$signed((8'hb8))};
                    end
                  for (forvar945 = (1'h0); (forvar945 < (1'h0)); forvar945 = (forvar945 + (1'h1)))
                    begin
                      reg946 <= $signed(forvar942);
                      reg947 <= $unsigned(reg863[(3'h5):(3'h5)]);
                      reg948 <= ((reg783[(3'h4):(1'h1)] ?
                              {$unsigned(reg749)} : $signed(reg937[(3'h5):(1'h0)])) ?
                          $unsigned(((~^reg781) ?
                              {reg765} : (reg914 >>> (8'ha4)))) : (($unsigned(reg882) | $signed(reg866)) ?
                              ($unsigned(reg852) || (reg756 << (8'haa))) : $signed(reg804)));
                      reg949 <= ({reg851[(2'h3):(1'h0)]} ?
                          (|(((8'hae) ? reg800 : reg862) ?
                              (reg765 ?
                                  reg835 : reg774) : $unsigned(reg792))) : $unsigned(((reg864 - reg888) ?
                              $signed(reg822) : reg790[(3'h5):(2'h3)])));
                    end
                  if (reg922)
                    begin
                      reg950 <= (reg792 >= $unsigned($unsigned($unsigned(reg791))));
                      reg951 <= (|($signed(((8'hab) ?
                          reg761 : reg846)) + ((reg791 ? reg761 : reg946) ?
                          (~&(8'had)) : reg938[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg950 <= ($unsigned(reg896[(1'h0):(1'h0)]) & (reg847 || (~|reg871)));
                    end
                end
            end
          for (forvar952 = (1'h0); (forvar952 < (2'h3)); forvar952 = (forvar952 + (1'h1)))
            begin
              reg953 <= reg901[(4'h8):(3'h6)];
              for (forvar954 = (1'h0); (forvar954 < (2'h3)); forvar954 = (forvar954 + (1'h1)))
                begin
                  for (forvar955 = (1'h0); (forvar955 < (2'h2)); forvar955 = (forvar955 + (1'h1)))
                    begin
                      reg956 <= (&$signed(((|forvar955) ?
                          ((8'hba) * forvar942) : {reg925})));
                      reg957 <= $unsigned(reg777[(1'h0):(1'h0)]);
                      reg958 <= {reg859};
                      reg959 <= (~&($unsigned(forvar933[(4'ha):(4'ha)]) + reg779[(3'h6):(2'h2)]));
                    end
                end
              reg960 <= (reg794 << ($unsigned(reg840) < {(8'ha3)}));
            end
        end
      else
        begin
          for (forvar941 = (1'h0); (forvar941 < (1'h1)); forvar941 = (forvar941 + (1'h1)))
            begin
              if (reg754[(2'h2):(1'h1)])
                begin
                  for (forvar942 = (1'h0); (forvar942 < (2'h3)); forvar942 = (forvar942 + (1'h1)))
                    begin
                      reg943 <= (^~$signed(($signed(reg812) >= reg889)));
                      reg944 <= reg861[(1'h0):(1'h0)];
                      reg945 <= $signed(($unsigned((~^reg828)) && $signed((8'ha0))));
                    end
                  reg946 <= (^~$signed(({reg912} - reg761)));
                  if ((~^reg847[(2'h2):(1'h1)]))
                    begin
                      reg947 <= $unsigned((+$unsigned((~^reg782))));
                      reg948 <= reg906[(2'h2):(1'h0)];
                      reg949 <= (8'hb3);
                    end
                  else
                    begin
                      reg947 <= $unsigned((^~(&reg888[(4'ha):(2'h3)])));
                      reg948 <= ({(~&forvar926[(2'h2):(1'h1)])} <<< (^~((reg757 ^~ reg888) ?
                          $signed((8'ha9)) : (reg936 && reg959))));
                      reg949 <= $signed({({reg863} + reg949)});
                    end
                end
              else
                begin
                  if ($unsigned(reg917[(4'h8):(2'h3)]))
                    begin
                      reg942 <= $unsigned({((8'haa) ?
                              $unsigned(reg911) : {reg932})});
                      reg943 <= reg819;
                      reg944 <= $unsigned(reg750);
                    end
                  else
                    begin
                      reg942 <= $unsigned(((~reg796[(2'h3):(1'h0)]) <= ((|(8'ha6)) ?
                          (reg946 >>> (8'hb1)) : $unsigned(forvar942))));
                      reg943 <= ($unsigned($signed((8'hba))) ?
                          $unsigned({reg958[(4'ha):(4'h9)]}) : $unsigned((reg912 ?
                              (reg805 << reg779) : (^reg825))));
                      reg944 <= (!$signed((reg817 + (8'hb1))));
                      reg945 <= {(~&((reg869 ? reg757 : reg914) << (8'hb5)))};
                    end
                  if (((~reg958) >>> ($signed(reg908[(3'h6):(3'h5)]) ?
                      (~&{reg875}) : reg878)))
                    begin
                      reg946 <= $signed((!reg797[(2'h3):(2'h3)]));
                      reg947 <= reg770;
                    end
                  else
                    begin
                      reg946 <= (wire740 | ((|$signed(wire838)) ?
                          $signed($unsigned(reg878)) : forvar924));
                    end
                  for (forvar948 = (1'h0); (forvar948 < (1'h0)); forvar948 = (forvar948 + (1'h1)))
                    begin
                      reg949 <= reg835[(2'h3):(1'h1)];
                      reg950 <= $unsigned(($unsigned(wire745) <<< ((!wire743) == $signed(reg921))));
                      reg951 <= reg795[(2'h2):(1'h1)];
                      reg952 <= (8'hb9);
                    end
                  for (forvar953 = (1'h0); (forvar953 < (2'h3)); forvar953 = (forvar953 + (1'h1)))
                    begin
                      reg954 <= (reg877[(2'h3):(1'h1)] ?
                          $unsigned(reg891[(4'h8):(3'h7)]) : ((+$signed(reg781)) ?
                              reg819 : reg857[(3'h5):(2'h2)]));
                      reg955 <= $unsigned((-reg946));
                      reg956 <= reg888[(3'h6):(3'h4)];
                    end
                end
              for (forvar957 = (1'h0); (forvar957 < (1'h0)); forvar957 = (forvar957 + (1'h1)))
                begin
                  for (forvar958 = (1'h0); (forvar958 < (2'h2)); forvar958 = (forvar958 + (1'h1)))
                    begin
                      reg959 <= reg889[(3'h5):(1'h1)];
                    end
                end
              for (forvar960 = (1'h0); (forvar960 < (1'h1)); forvar960 = (forvar960 + (1'h1)))
                begin
                  for (forvar961 = (1'h0); (forvar961 < (2'h3)); forvar961 = (forvar961 + (1'h1)))
                    begin
                      reg962 <= ({((reg786 >>> (8'haa)) * (~&reg948))} && $signed($signed(reg907[(2'h2):(1'h0)])));
                      reg963 <= (+(^$signed({reg949})));
                      reg964 <= ((reg761[(1'h0):(1'h0)] > reg788[(1'h1):(1'h0)]) ?
                          ((|reg960[(3'h7):(3'h6)]) ~^ $unsigned($signed(reg919))) : reg923);
                      reg965 <= ($unsigned(reg791[(4'hc):(4'hc)]) ?
                          {$signed((8'hab))} : (-((reg917 ^~ reg760) ?
                              ((8'haa) ? reg868 : reg855) : (|reg886))));
                    end
                  reg966 <= $signed($unsigned(reg787));
                end
            end
          for (forvar967 = (1'h0); (forvar967 < (1'h0)); forvar967 = (forvar967 + (1'h1)))
            begin
              if ({wire741})
                begin
                  if ($unsigned($unsigned(reg754[(2'h3):(1'h0)])))
                    begin
                      reg968 <= {reg905[(2'h2):(2'h2)]};
                      reg969 <= reg907;
                    end
                  else
                    begin
                      reg968 <= (reg968[(2'h2):(1'h0)] ?
                          (($unsigned(reg863) & (reg878 >> reg881)) || reg826[(1'h0):(1'h0)]) : reg953);
                    end
                  for (forvar970 = (1'h0); (forvar970 < (2'h3)); forvar970 = (forvar970 + (1'h1)))
                    begin
                      reg971 <= (8'hb2);
                      reg972 <= (~(wire744[(1'h0):(1'h0)] && (~^{reg794})));
                    end
                end
              else
                begin
                  for (forvar968 = (1'h0); (forvar968 < (1'h1)); forvar968 = (forvar968 + (1'h1)))
                    begin
                      reg969 <= reg938[(2'h2):(1'h1)];
                      reg970 <= (reg783 ?
                          $signed(reg832[(2'h2):(2'h2)]) : {reg934});
                      reg971 <= ((|($signed(reg861) ?
                              reg833 : $signed((8'had)))) ?
                          {(&$unsigned(reg878))} : $unsigned($unsigned({(8'haf)})));
                    end
                  if (({$unsigned($signed(reg958))} ?
                      reg928[(3'h5):(3'h5)] : $unsigned((8'h9e))))
                    begin
                      reg972 <= reg954;
                      reg973 <= $signed(($unsigned($unsigned(forvar953)) & (8'hac)));
                    end
                  else
                    begin
                      reg972 <= (|$signed(($signed(forvar958) ^ (8'hb4))));
                      reg973 <= (($signed((8'ha3)) & (reg971 ^ (^reg960))) ?
                          ($unsigned($unsigned(reg846)) ?
                              ($signed((8'hb8)) >= $signed(reg959)) : forvar948[(3'h5):(3'h5)]) : (|$unsigned((reg905 != reg840))));
                      reg974 <= (~^forvar942);
                    end
                  if ((($signed((^reg864)) ?
                      (+(wire742 ?
                          reg752 : reg891)) : {{reg756}}) * (^~(reg884 ?
                      (8'h9f) : reg795))))
                    begin
                      reg975 <= $signed((|({reg880} + reg780[(3'h4):(2'h3)])));
                      reg976 <= ((({reg959} != $signed(reg957)) ?
                          {reg882[(2'h2):(1'h1)]} : forvar954) & $unsigned((reg874 - reg929[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg975 <= ((8'h9f) ?
                          $unsigned(reg959) : {$signed(reg840)});
                      reg976 <= $signed((-(reg872 ?
                          $signed(reg874) : $signed(forvar941))));
                      reg977 <= (~(((reg823 ? wire838 : reg850) ?
                              reg976 : (reg867 & reg868)) ?
                          ((reg756 ? forvar952 : reg844) + (reg890 ?
                              forvar967 : reg751)) : $signed((reg797 > (8'haf)))));
                      reg978 <= ({reg796[(3'h5):(3'h4)]} ^~ $unsigned($signed($signed((8'h9d)))));
                    end
                end
              for (forvar979 = (1'h0); (forvar979 < (1'h1)); forvar979 = (forvar979 + (1'h1)))
                begin
                  for (forvar980 = (1'h0); (forvar980 < (2'h3)); forvar980 = (forvar980 + (1'h1)))
                    begin
                      reg981 <= $signed($signed($unsigned(reg947[(1'h0):(1'h0)])));
                      reg982 <= ((reg939[(2'h2):(1'h0)] + (reg965 ?
                          reg769[(2'h2):(1'h1)] : $unsigned(reg880))) ^ ((^$signed(reg949)) ^ (reg828 ?
                          {reg778} : (reg923 > reg796))));
                      reg983 <= forvar954;
                      reg984 <= {reg837[(2'h3):(2'h2)]};
                    end
                end
              if (($unsigned($unsigned((-(8'hb9)))) ?
                  reg947 : $unsigned(reg792)))
                begin
                  for (forvar985 = (1'h0); (forvar985 < (1'h0)); forvar985 = (forvar985 + (1'h1)))
                    begin
                      reg986 <= $signed(reg901);
                    end
                end
              else
                begin
                  reg985 <= $unsigned(reg775);
                  reg986 <= (~|$signed((^~(~^reg770))));
                  if ($signed($signed($signed({reg965}))))
                    begin
                      reg987 <= reg880[(1'h1):(1'h0)];
                      reg988 <= (-(~({(8'h9d)} << (&reg935))));
                      reg989 <= $unsigned((((reg799 ?
                          (8'ha4) : reg912) ~^ (reg817 >> reg969)) | {reg953}));
                      reg990 <= ($unsigned(reg883[(4'h9):(2'h2)]) ?
                          $signed(reg858) : $unsigned((reg785 && reg845)));
                    end
                  else
                    begin
                      reg987 <= (reg832 - $signed(reg783));
                      reg988 <= $signed(reg988);
                      reg989 <= (^(((forvar958 ? reg916 : reg935) ?
                          (reg893 <<< reg873) : (^reg931)) ^~ ($unsigned(reg950) ?
                          {reg866} : ((8'hab) ? reg836 : (8'hba)))));
                    end
                end
            end
          for (forvar991 = (1'h0); (forvar991 < (2'h3)); forvar991 = (forvar991 + (1'h1)))
            begin
              if ($unsigned(($unsigned($unsigned(reg934)) || reg794)))
                begin
                  reg992 <= ({((reg963 ?
                          reg956 : reg871) < $signed(forvar961))} >> ($signed($signed(forvar957)) && ($unsigned(reg956) >>> (reg763 <<< reg874))));
                end
              else
                begin
                  for (forvar992 = (1'h0); (forvar992 < (1'h0)); forvar992 = (forvar992 + (1'h1)))
                    begin
                      reg993 <= reg791;
                      reg994 <= $signed({($signed(forvar952) ~^ forvar960[(1'h1):(1'h1)])});
                      reg995 <= (|reg958);
                      reg996 <= ($signed(($signed(reg958) ?
                              reg752 : (|reg784))) ?
                          $signed(reg988[(1'h1):(1'h1)]) : forvar992);
                    end
                end
              for (forvar997 = (1'h0); (forvar997 < (1'h0)); forvar997 = (forvar997 + (1'h1)))
                begin
                  if (reg884[(3'h6):(2'h3)])
                    begin
                      reg998 <= $signed(reg772[(2'h2):(1'h1)]);
                      reg999 <= forvar925;
                    end
                  else
                    begin
                      reg998 <= (|($unsigned($signed(forvar991)) ^ $unsigned((reg943 ^~ forvar985))));
                      reg999 <= {(8'hb3)};
                      reg1000 <= $signed((~|((reg888 >>> reg858) ?
                          reg855 : $signed(reg784))));
                    end
                  reg1001 <= (~$unsigned(reg925));
                end
              reg1002 <= ((reg994 ?
                  (|(reg772 ?
                      reg845 : reg829)) : reg763) < forvar968[(2'h2):(1'h1)]);
            end
          if ({reg750})
            begin
              if ({reg818})
                begin
                  for (forvar1003 = (1'h0); (forvar1003 < (2'h3)); forvar1003 = (forvar1003 + (1'h1)))
                    begin
                      reg1004 <= reg859;
                      reg1005 <= $signed($signed((((8'haf) | reg808) ?
                          (^~reg977) : $signed((8'haf)))));
                    end
                  for (forvar1006 = (1'h0); (forvar1006 < (1'h1)); forvar1006 = (forvar1006 + (1'h1)))
                    begin
                      reg1007 <= ((reg995 | (reg867[(1'h0):(1'h0)] ?
                          (wire740 ? reg755 : reg808) : forvar952)) ^ (8'hab));
                      reg1008 <= $unsigned({($signed(reg825) != $unsigned(reg761))});
                      reg1009 <= $unsigned({reg950});
                      reg1010 <= (8'hb1);
                    end
                end
              else
                begin
                  if ($signed(($signed($unsigned(reg993)) ?
                      ($signed((8'ha9)) > $signed(reg877)) : reg878)))
                    begin
                      reg1003 <= (|{($unsigned(reg858) ?
                              reg777[(1'h0):(1'h0)] : $signed(reg845))});
                      reg1004 <= $unsigned(reg987);
                      reg1005 <= ((({reg1007} ?
                              reg824[(1'h1):(1'h0)] : reg883[(3'h5):(3'h5)]) || ($unsigned(reg889) ?
                              ((8'ha2) * reg947) : $unsigned((8'ha5)))) ?
                          $signed($unsigned((reg951 + reg911))) : $signed({(-reg853)}));
                    end
                  else
                    begin
                      reg1003 <= $unsigned(($unsigned(reg874) ?
                          forvar961[(1'h0):(1'h0)] : (+reg931[(2'h2):(2'h2)])));
                      reg1004 <= ({((|reg915) <<< (-reg888))} && reg859);
                      reg1005 <= (8'hb4);
                    end
                  for (forvar1006 = (1'h0); (forvar1006 < (1'h1)); forvar1006 = (forvar1006 + (1'h1)))
                    begin
                      reg1007 <= $unsigned((|{reg798}));
                      reg1008 <= $signed(($unsigned((reg893 ?
                              reg960 : reg893)) ?
                          ($unsigned(reg882) < (reg904 ?
                              reg946 : reg976)) : reg750[(2'h3):(2'h2)]));
                      reg1009 <= $signed($unsigned($signed((reg820 ?
                          reg871 : (8'hae)))));
                      reg1010 <= reg952[(3'h4):(2'h3)];
                    end
                  for (forvar1011 = (1'h0); (forvar1011 < (1'h1)); forvar1011 = (forvar1011 + (1'h1)))
                    begin
                      reg1012 <= $signed($unsigned($unsigned(reg827)));
                      reg1013 <= $unsigned(reg800);
                      reg1014 <= $unsigned(reg776[(4'ha):(1'h1)]);
                    end
                  for (forvar1015 = (1'h0); (forvar1015 < (1'h1)); forvar1015 = (forvar1015 + (1'h1)))
                    begin
                      reg1016 <= $signed($signed($unsigned($unsigned(reg788))));
                      reg1017 <= $signed(reg761);
                      reg1018 <= ($unsigned($unsigned((reg936 ?
                          reg959 : forvar960))) ^~ reg825);
                      reg1019 <= $signed($signed($unsigned(((8'ha3) ?
                          reg779 : (8'hb3)))));
                    end
                end
            end
          else
            begin
              for (forvar1003 = (1'h0); (forvar1003 < (2'h3)); forvar1003 = (forvar1003 + (1'h1)))
                begin
                  for (forvar1004 = (1'h0); (forvar1004 < (2'h3)); forvar1004 = (forvar1004 + (1'h1)))
                    begin
                      reg1005 <= {($unsigned(reg932) ?
                              reg824 : (~&(reg927 ? reg837 : reg811)))};
                    end
                  if (((reg840[(1'h0):(1'h0)] ?
                      reg969 : {(~&reg765)}) & ((!(+reg750)) ?
                      (|(&reg939)) : $unsigned({forvar970}))))
                    begin
                      reg1006 <= (!($unsigned({(8'had)}) | (!((8'ha7) - reg810))));
                      reg1007 <= $unsigned($signed(reg999));
                    end
                  else
                    begin
                      reg1006 <= reg982[(4'hd):(2'h3)];
                      reg1007 <= (8'ha0);
                    end
                  for (forvar1008 = (1'h0); (forvar1008 < (2'h2)); forvar1008 = (forvar1008 + (1'h1)))
                    begin
                      reg1009 <= $signed(reg1004[(2'h3):(2'h2)]);
                      reg1010 <= ((^$unsigned((forvar953 ~^ reg915))) ?
                          $signed(reg1004) : ($unsigned(reg757) ?
                              ($signed(forvar954) ^ (^reg763)) : (&$signed(reg972))));
                    end
                end
              reg1011 <= $unsigned({forvar925[(1'h1):(1'h0)]});
            end
        end
      for (forvar1020 = (1'h0); (forvar1020 < (1'h0)); forvar1020 = (forvar1020 + (1'h1)))
        begin
          for (forvar1021 = (1'h0); (forvar1021 < (2'h3)); forvar1021 = (forvar1021 + (1'h1)))
            begin
              for (forvar1022 = (1'h0); (forvar1022 < (2'h3)); forvar1022 = (forvar1022 + (1'h1)))
                begin
                  if ({(8'hba)})
                    begin
                      reg1023 <= $signed({(|((8'ha3) ? reg918 : forvar991))});
                      reg1024 <= (+$signed($unsigned(reg754)));
                      reg1025 <= ((reg861[(2'h3):(2'h2)] ?
                              $unsigned((reg858 ? reg818 : reg926)) : reg764) ?
                          $signed({(reg970 ?
                                  (8'hb9) : reg901)}) : {(~|(reg807 * reg951))});
                    end
                  else
                    begin
                      reg1023 <= (&reg877[(1'h1):(1'h1)]);
                    end
                end
            end
        end
      reg1026 <= $signed((^~(&(^reg969))));
    end
  always
    @(posedge clk) begin
      for (forvar1027 = (1'h0); (forvar1027 < (1'h1)); forvar1027 = (forvar1027 + (1'h1)))
        begin
          for (forvar1028 = (1'h0); (forvar1028 < (1'h0)); forvar1028 = (forvar1028 + (1'h1)))
            begin
              if ($unsigned(($signed(reg926) < reg910[(3'h6):(3'h4)])))
                begin
                  if (($signed(reg962) ?
                      $unsigned($signed(reg883[(1'h1):(1'h0)])) : $signed((^~(reg891 ?
                          reg784 : (8'ha1))))))
                    begin
                      reg1029 <= $unsigned(reg949);
                      reg1030 <= (~|reg1001[(3'h6):(1'h0)]);
                      reg1031 <= ($unsigned($signed({(8'ha1)})) ?
                          (~(reg797[(1'h0):(1'h0)] ?
                              reg772 : (wire741 ?
                                  reg782 : reg998))) : $signed(($unsigned((8'hb9)) && $signed(reg761))));
                      reg1032 <= (reg951 ~^ (~|(&(reg781 ?
                          reg880 : forvar1027))));
                    end
                  else
                    begin
                      reg1029 <= reg988[(2'h2):(1'h1)];
                      reg1030 <= (~|($unsigned($signed(reg857)) ?
                          $unsigned($unsigned((8'ha3))) : (^reg822)));
                      reg1031 <= reg888[(1'h1):(1'h0)];
                      reg1032 <= reg828;
                    end
                  for (forvar1033 = (1'h0); (forvar1033 < (1'h0)); forvar1033 = (forvar1033 + (1'h1)))
                    begin
                      reg1034 <= reg929;
                      reg1035 <= reg988[(3'h4):(2'h2)];
                    end
                  for (forvar1036 = (1'h0); (forvar1036 < (2'h3)); forvar1036 = (forvar1036 + (1'h1)))
                    begin
                      reg1037 <= $unsigned({reg1006});
                      reg1038 <= {$unsigned(((8'hb7) != $signed(reg791)))};
                    end
                end
              else
                begin
                  for (forvar1029 = (1'h0); (forvar1029 < (1'h0)); forvar1029 = (forvar1029 + (1'h1)))
                    begin
                      reg1030 <= {reg822[(4'h9):(4'h8)]};
                      reg1031 <= ((~&($unsigned(reg848) >= $signed(reg761))) ^ (reg1005 < $signed((reg824 ?
                          reg894 : reg749))));
                      reg1032 <= $signed($unsigned($signed(reg990[(4'h8):(1'h1)])));
                    end
                end
            end
          if ((reg817 ?
              (($unsigned(reg1017) ^ $signed(reg767)) ?
                  ($unsigned(reg799) | ((8'hb1) <= (8'haa))) : ((reg984 + reg750) ?
                      {reg819} : ((8'hb5) ? reg905 : reg972))) : reg922))
            begin
              for (forvar1039 = (1'h0); (forvar1039 < (1'h1)); forvar1039 = (forvar1039 + (1'h1)))
                begin
                  if (reg1007[(4'h8):(3'h5)])
                    begin
                      reg1040 <= {$unsigned(((8'ha6) || $unsigned(reg993)))};
                    end
                  else
                    begin
                      reg1040 <= {$unsigned(reg859[(1'h1):(1'h0)])};
                      reg1041 <= ((|(reg952[(3'h5):(2'h3)] == reg797)) ~^ (-(forvar1039 != {reg876})));
                    end
                end
              for (forvar1042 = (1'h0); (forvar1042 < (1'h0)); forvar1042 = (forvar1042 + (1'h1)))
                begin
                  reg1043 <= $signed($signed((~((8'ha2) ? (8'h9e) : reg858))));
                  for (forvar1044 = (1'h0); (forvar1044 < (1'h1)); forvar1044 = (forvar1044 + (1'h1)))
                    begin
                      reg1045 <= ({reg950} || (8'hb9));
                    end
                end
              for (forvar1046 = (1'h0); (forvar1046 < (1'h1)); forvar1046 = (forvar1046 + (1'h1)))
                begin
                  if ((($signed($signed((8'hac))) && {reg751}) ?
                      ((reg779[(1'h0):(1'h0)] != reg880) | (~(reg811 ?
                          reg820 : (8'h9c)))) : $signed((&$signed(reg895)))))
                    begin
                      reg1047 <= $unsigned(($unsigned($signed(reg900)) ?
                          ({reg940} < $unsigned(reg926)) : (reg811 ?
                              (+reg850) : $unsigned(reg882))));
                      reg1048 <= ((~&reg1007) >> reg806);
                      reg1049 <= reg894[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg1047 <= (8'haa);
                      reg1048 <= ($unsigned(reg798) ?
                          $unsigned(reg825) : reg993);
                    end
                  reg1050 <= reg822;
                end
            end
          else
            begin
              for (forvar1039 = (1'h0); (forvar1039 < (1'h0)); forvar1039 = (forvar1039 + (1'h1)))
                begin
                  reg1040 <= {(|(reg944 ?
                          ((8'hb1) ? reg1049 : reg767) : forvar1029))};
                  if ({((~^(reg950 - reg917)) | $signed((+reg750)))})
                    begin
                      reg1041 <= ($signed($unsigned($signed((8'hb7)))) ?
                          reg855 : $signed($signed(reg944[(3'h5):(2'h2)])));
                      reg1042 <= ((^((wire744 || (8'ha4)) ?
                          $unsigned((8'hb7)) : $unsigned(reg790))) - reg1029[(1'h0):(1'h0)]);
                      reg1043 <= $unsigned(reg939[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg1041 <= (^$signed(($signed(reg801) - (reg914 ?
                          reg889 : reg756))));
                      reg1042 <= reg929;
                      reg1043 <= $unsigned(($unsigned(reg1017[(1'h0):(1'h0)]) ?
                          reg863 : ((reg1019 ? reg987 : reg897) ?
                              (reg849 >= reg862) : (8'ha7))));
                      reg1044 <= (-{(&reg981)});
                    end
                  for (forvar1045 = (1'h0); (forvar1045 < (2'h2)); forvar1045 = (forvar1045 + (1'h1)))
                    begin
                      reg1046 <= reg765;
                      reg1047 <= (reg1001[(3'h5):(3'h5)] ~^ reg761[(1'h1):(1'h1)]);
                    end
                  for (forvar1048 = (1'h0); (forvar1048 < (1'h1)); forvar1048 = (forvar1048 + (1'h1)))
                    begin
                      reg1049 <= (reg794 ?
                          reg774 : {((reg976 && reg910) >> (reg827 != reg869))});
                      reg1050 <= $signed((^~$signed($unsigned(forvar1028))));
                    end
                end
              reg1051 <= reg992[(1'h0):(1'h0)];
            end
          if (((^~(reg799[(3'h7):(1'h1)] ?
              reg853[(1'h0):(1'h0)] : (8'ha9))) <= $signed($unsigned(reg1016))))
            begin
              for (forvar1052 = (1'h0); (forvar1052 < (2'h2)); forvar1052 = (forvar1052 + (1'h1)))
                begin
                  if (({wire745} ^~ reg972))
                    begin
                      reg1053 <= ((reg948 ?
                          $signed(reg851[(1'h1):(1'h0)]) : reg914) ^ reg848);
                      reg1054 <= (^~($unsigned(reg785[(2'h2):(1'h1)]) ?
                          {(8'ha1)} : ($signed(reg1049) ?
                              reg893 : ((8'ha4) ? reg1001 : reg849))));
                      reg1055 <= (8'hb8);
                      reg1056 <= (-($unsigned((8'hb3)) ?
                          (8'ha8) : ({reg789} ?
                              $unsigned(reg889) : reg1030[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg1053 <= reg858[(2'h3):(1'h0)];
                      reg1054 <= $signed(reg775[(2'h2):(1'h1)]);
                      reg1055 <= $signed(($signed(reg959[(2'h2):(2'h2)]) * ($signed(reg1030) || $signed(forvar1052))));
                    end
                end
              for (forvar1057 = (1'h0); (forvar1057 < (2'h2)); forvar1057 = (forvar1057 + (1'h1)))
                begin
                  if ((reg918[(4'hb):(1'h0)] ?
                      $unsigned({(wire743 & (8'ha4))}) : (^~({reg882} ^ {reg950}))))
                    begin
                      reg1058 <= (reg847 * (((~|reg978) ? (~reg954) : reg1005) ?
                          ((reg848 ?
                              reg956 : reg1006) & (^reg861)) : (^(reg811 ?
                              reg931 : reg1019))));
                      reg1059 <= reg973[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg1058 <= (+reg749);
                      reg1059 <= {{$unsigned(reg817[(2'h3):(1'h1)])}};
                      reg1060 <= ((($signed(wire740) ?
                                  reg829[(3'h5):(2'h3)] : $signed(reg1003)) ?
                              ($signed(reg982) <<< (wire740 <= reg1012)) : $signed((reg866 ?
                                  reg840 : reg785))) ?
                          (^$signed((~(8'haf)))) : (($signed(reg846) ?
                                  (reg931 > (8'h9c)) : reg905[(1'h0):(1'h0)]) ?
                              ($unsigned(reg942) ?
                                  (reg864 <= (8'had)) : (wire745 ?
                                      reg1001 : reg1041)) : reg1018[(2'h3):(2'h3)]));
                      reg1061 <= reg892;
                    end
                  if (((-$signed({reg960})) ^ $signed((reg965[(3'h7):(3'h7)] ?
                      (&reg1016) : reg846))))
                    begin
                      reg1062 <= $signed(({$signed(reg849)} ~^ ($signed(reg1004) ?
                          $signed((8'hb3)) : (forvar1027 * forvar1036))));
                    end
                  else
                    begin
                      reg1062 <= $signed((~^{$signed(reg889)}));
                      reg1063 <= reg807;
                    end
                  for (forvar1064 = (1'h0); (forvar1064 < (1'h1)); forvar1064 = (forvar1064 + (1'h1)))
                    begin
                      reg1065 <= {$signed((reg804 ? reg773 : (-reg955)))};
                    end
                end
              if ($unsigned((($signed((8'ha7)) != (reg817 ? (8'hae) : reg773)) ?
                  (8'hab) : {(~^reg804)})))
                begin
                  if (($signed((|((8'hb2) ? reg1062 : reg999))) ?
                      (!($signed(reg782) ?
                          reg770[(1'h0):(1'h0)] : (reg820 ?
                              reg858 : reg872))) : (reg835[(4'h8):(3'h5)] ?
                          reg925[(4'hb):(2'h3)] : $signed((~^forvar1042)))))
                    begin
                      reg1066 <= reg886;
                      reg1067 <= (((&(reg1031 ?
                          reg966 : reg1004)) >> forvar1048) << ((reg754 && {reg827}) || $signed((-reg994))));
                    end
                  else
                    begin
                      reg1066 <= ($signed(reg1013[(3'h5):(3'h5)]) ?
                          reg785[(3'h5):(1'h1)] : $unsigned((~|((8'ha7) ~^ reg867))));
                      reg1067 <= forvar1048[(2'h2):(1'h1)];
                      reg1068 <= $unsigned(((reg1007[(4'h9):(3'h7)] ?
                              $signed(reg938) : (~&reg780)) ?
                          ($unsigned((8'hae)) ?
                              $signed(reg812) : $signed(reg956)) : (8'hae)));
                    end
                  for (forvar1069 = (1'h0); (forvar1069 < (2'h2)); forvar1069 = (forvar1069 + (1'h1)))
                    begin
                      reg1070 <= reg925[(3'h6):(2'h2)];
                      reg1071 <= (reg799[(2'h3):(1'h0)] ? reg836 : reg817);
                      reg1072 <= (~|((reg810[(3'h4):(1'h1)] & $unsigned(reg800)) ~^ $signed(reg886)));
                    end
                  for (forvar1073 = (1'h0); (forvar1073 < (1'h1)); forvar1073 = (forvar1073 + (1'h1)))
                    begin
                      reg1074 <= {reg777};
                      reg1075 <= $unsigned((($signed(reg1003) + $unsigned(reg940)) ?
                          $unsigned($unsigned((8'had))) : $signed(reg760[(1'h0):(1'h0)])));
                      reg1076 <= (|(~&((reg1062 ?
                          reg996 : reg818) ^ $signed(reg926))));
                      reg1077 <= ($unsigned($signed($unsigned(reg810))) > (^~reg1016));
                    end
                end
              else
                begin
                  for (forvar1066 = (1'h0); (forvar1066 < (1'h0)); forvar1066 = (forvar1066 + (1'h1)))
                    begin
                      reg1067 <= ($unsigned(reg975[(4'hb):(3'h5)]) & (8'ha1));
                    end
                  for (forvar1068 = (1'h0); (forvar1068 < (2'h3)); forvar1068 = (forvar1068 + (1'h1)))
                    begin
                      reg1069 <= (&reg1051[(3'h4):(3'h4)]);
                    end
                  for (forvar1070 = (1'h0); (forvar1070 < (1'h0)); forvar1070 = (forvar1070 + (1'h1)))
                    begin
                      reg1071 <= reg893;
                    end
                end
            end
          else
            begin
              if ($signed($unsigned(reg993[(3'h4):(2'h3)])))
                begin
                  for (forvar1052 = (1'h0); (forvar1052 < (2'h3)); forvar1052 = (forvar1052 + (1'h1)))
                    begin
                      reg1053 <= (8'ha0);
                      reg1054 <= (-reg995[(2'h2):(1'h0)]);
                      reg1055 <= (~^(^reg878[(3'h4):(3'h4)]));
                    end
                  reg1056 <= $unsigned(($unsigned((8'hac)) - (((8'h9c) >>> (8'ha8)) ?
                      reg983[(3'h7):(2'h2)] : (reg969 >>> reg948))));
                  reg1057 <= reg1032;
                  for (forvar1058 = (1'h0); (forvar1058 < (2'h3)); forvar1058 = (forvar1058 + (1'h1)))
                    begin
                      reg1059 <= ($unsigned(($unsigned(reg790) ?
                              reg846[(4'hb):(4'h9)] : $unsigned(reg800))) ?
                          reg1045 : {(~|(~&reg925))});
                    end
                end
              else
                begin
                  for (forvar1052 = (1'h0); (forvar1052 < (2'h2)); forvar1052 = (forvar1052 + (1'h1)))
                    begin
                      reg1053 <= $unsigned($signed(reg818));
                      reg1054 <= forvar1033[(4'h9):(4'h8)];
                      reg1055 <= reg818;
                      reg1056 <= $unsigned(reg807);
                    end
                  for (forvar1057 = (1'h0); (forvar1057 < (1'h1)); forvar1057 = (forvar1057 + (1'h1)))
                    begin
                      reg1058 <= ($signed(reg823) + ((!(!reg981)) ?
                          reg1034 : ((forvar1029 ?
                              reg914 : reg901) || ((8'haf) ?
                              reg756 : reg1032))));
                      reg1059 <= (reg801[(1'h1):(1'h0)] * reg876[(4'h8):(2'h2)]);
                    end
                end
              reg1060 <= $unsigned(((forvar1042[(3'h4):(2'h2)] ?
                  $unsigned(reg976) : $unsigned(wire743)) <= reg932[(4'hd):(3'h6)]));
            end
          for (forvar1078 = (1'h0); (forvar1078 < (1'h0)); forvar1078 = (forvar1078 + (1'h1)))
            begin
              reg1079 <= (~|{reg964});
              if ({reg888})
                begin
                  for (forvar1080 = (1'h0); (forvar1080 < (2'h3)); forvar1080 = (forvar1080 + (1'h1)))
                    begin
                      reg1081 <= ((~^(~reg801)) ?
                          (+(((8'h9c) <= reg824) << (~^reg981))) : ($signed({reg919}) ^ (~|reg787)));
                      reg1082 <= reg1037;
                      reg1083 <= (($unsigned($unsigned(reg1040)) | $signed((^reg996))) ?
                          (~reg993[(1'h0):(1'h0)]) : (({reg1050} * $unsigned(reg889)) ?
                              reg1040 : reg937));
                    end
                end
              else
                begin
                  for (forvar1080 = (1'h0); (forvar1080 < (2'h3)); forvar1080 = (forvar1080 + (1'h1)))
                    begin
                      reg1081 <= reg1061;
                      reg1082 <= $signed((reg828 < (^~$signed(reg940))));
                      reg1083 <= forvar1033[(3'h6):(2'h2)];
                      reg1084 <= reg956[(1'h1):(1'h0)];
                    end
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module5
#(parameter param628 = ((~|(&(+(8'ha1)))) ? ((((8'h9e) || (8'hba)) + {(8'hba)}) ? ((^(8'had)) ? {(8'hae)} : (~&(8'hb1))) : {(~&(8'ha9))}) : ((((8'hae) ? (8'hb4) : (8'haa)) ? (8'ha5) : ((8'hac) ? (8'hae) : (8'ha4))) ? (|((8'hb5) ? (8'hac) : (8'hb6))) : {((8'hb3) ? (8'hba) : (8'ha1))})))
(y, clk, wire10, wire9, wire8, wire7, wire6);
  output wire [(32'h1455):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire10;
  input wire signed [(3'h5):(1'h0)] wire9;
  input wire [(3'h6):(1'h0)] wire8;
  input wire [(4'he):(1'h0)] wire7;
  input wire [(4'hb):(1'h0)] wire6;
  wire [(4'hf):(1'h0)] wire627;
  wire [(4'hc):(1'h0)] wire535;
  wire signed [(2'h2):(1'h0)] wire268;
  wire [(4'ha):(1'h0)] wire267;
  wire [(4'h8):(1'h0)] wire266;
  wire signed [(4'h8):(1'h0)] wire265;
  wire [(3'h5):(1'h0)] wire11;
  reg signed [(4'h9):(1'h0)] reg626 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg625 = (1'h0);
  reg [(4'h9):(1'h0)] reg624 = (1'h0);
  reg [(4'h8):(1'h0)] reg622 = (1'h0);
  reg [(2'h2):(1'h0)] reg621 = (1'h0);
  reg [(4'ha):(1'h0)] reg620 = (1'h0);
  reg [(4'h8):(1'h0)] reg619 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg618 = (1'h0);
  reg [(4'h8):(1'h0)] reg617 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg616 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg615 = (1'h0);
  reg [(3'h5):(1'h0)] reg613 = (1'h0);
  reg [(4'ha):(1'h0)] reg611 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg608 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg607 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg606 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg604 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg603 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg602 = (1'h0);
  reg [(4'hb):(1'h0)] reg601 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg600 = (1'h0);
  reg [(4'ha):(1'h0)] reg599 = (1'h0);
  reg [(4'hd):(1'h0)] reg597 = (1'h0);
  reg [(4'h8):(1'h0)] reg595 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg592 = (1'h0);
  reg [(5'h10):(1'h0)] reg587 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg572 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg567 = (1'h0);
  reg [(3'h6):(1'h0)] reg551 = (1'h0);
  reg [(4'hd):(1'h0)] reg542 = (1'h0);
  reg [(4'hd):(1'h0)] reg540 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg591 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg590 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg589 = (1'h0);
  reg signed [(4'he):(1'h0)] reg588 = (1'h0);
  reg [(2'h3):(1'h0)] reg586 = (1'h0);
  reg [(3'h4):(1'h0)] reg585 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg584 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg583 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg581 = (1'h0);
  reg [(3'h4):(1'h0)] reg580 = (1'h0);
  reg [(4'hb):(1'h0)] reg579 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg578 = (1'h0);
  reg signed [(4'he):(1'h0)] reg576 = (1'h0);
  reg [(4'hc):(1'h0)] reg575 = (1'h0);
  reg [(2'h2):(1'h0)] reg574 = (1'h0);
  reg [(4'he):(1'h0)] reg573 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg571 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg570 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg569 = (1'h0);
  reg [(4'he):(1'h0)] reg568 = (1'h0);
  reg [(4'hd):(1'h0)] reg566 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg565 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg564 = (1'h0);
  reg [(4'hf):(1'h0)] reg563 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg562 = (1'h0);
  reg [(4'hb):(1'h0)] reg561 = (1'h0);
  reg [(2'h2):(1'h0)] reg560 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg559 = (1'h0);
  reg [(4'hd):(1'h0)] reg558 = (1'h0);
  reg [(4'h9):(1'h0)] reg557 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg556 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg555 = (1'h0);
  reg [(2'h2):(1'h0)] reg554 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg553 = (1'h0);
  reg [(4'hb):(1'h0)] reg552 = (1'h0);
  reg [(3'h7):(1'h0)] reg549 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg548 = (1'h0);
  reg [(3'h5):(1'h0)] reg547 = (1'h0);
  reg [(5'h10):(1'h0)] reg546 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg545 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg544 = (1'h0);
  reg [(3'h4):(1'h0)] reg543 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg541 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg538 = (1'h0);
  reg [(4'hf):(1'h0)] reg537 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg384 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg378 = (1'h0);
  reg [(4'ha):(1'h0)] reg382 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg381 = (1'h0);
  reg [(4'h9):(1'h0)] reg380 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg379 = (1'h0);
  reg [(5'h10):(1'h0)] reg377 = (1'h0);
  reg [(4'ha):(1'h0)] reg374 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg370 = (1'h0);
  reg [(4'h9):(1'h0)] reg366 = (1'h0);
  reg [(4'hb):(1'h0)] reg373 = (1'h0);
  reg [(2'h2):(1'h0)] reg372 = (1'h0);
  reg [(5'h10):(1'h0)] reg371 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg369 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg368 = (1'h0);
  reg [(3'h5):(1'h0)] reg367 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg365 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg363 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg362 = (1'h0);
  reg [(3'h4):(1'h0)] reg348 = (1'h0);
  reg [(4'hc):(1'h0)] reg343 = (1'h0);
  reg [(4'hc):(1'h0)] reg341 = (1'h0);
  reg [(2'h3):(1'h0)] reg336 = (1'h0);
  reg [(4'ha):(1'h0)] reg335 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg333 = (1'h0);
  reg [(3'h4):(1'h0)] reg329 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg318 = (1'h0);
  reg [(2'h3):(1'h0)] reg321 = (1'h0);
  reg [(4'h9):(1'h0)] reg320 = (1'h0);
  reg [(3'h4):(1'h0)] reg360 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg359 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg358 = (1'h0);
  reg [(4'h9):(1'h0)] reg357 = (1'h0);
  reg [(2'h3):(1'h0)] reg355 = (1'h0);
  reg [(4'h9):(1'h0)] reg354 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg353 = (1'h0);
  reg [(4'he):(1'h0)] reg352 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg351 = (1'h0);
  reg [(3'h7):(1'h0)] reg350 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg347 = (1'h0);
  reg [(4'ha):(1'h0)] reg346 = (1'h0);
  reg [(4'hb):(1'h0)] reg345 = (1'h0);
  reg [(3'h4):(1'h0)] reg344 = (1'h0);
  reg [(3'h5):(1'h0)] reg342 = (1'h0);
  reg [(4'ha):(1'h0)] reg340 = (1'h0);
  reg [(5'h10):(1'h0)] reg339 = (1'h0);
  reg [(2'h3):(1'h0)] reg338 = (1'h0);
  reg [(4'hb):(1'h0)] reg337 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg334 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg332 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg331 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg328 = (1'h0);
  reg [(4'hd):(1'h0)] reg327 = (1'h0);
  reg [(4'h8):(1'h0)] reg326 = (1'h0);
  reg [(4'ha):(1'h0)] reg325 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg324 = (1'h0);
  reg [(4'ha):(1'h0)] reg323 = (1'h0);
  reg [(4'hd):(1'h0)] reg322 = (1'h0);
  reg [(2'h2):(1'h0)] reg319 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg317 = (1'h0);
  reg [(4'hb):(1'h0)] reg314 = (1'h0);
  reg [(3'h5):(1'h0)] reg311 = (1'h0);
  reg [(4'ha):(1'h0)] reg299 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg300 = (1'h0);
  reg signed [(4'he):(1'h0)] reg316 = (1'h0);
  reg signed [(4'he):(1'h0)] reg315 = (1'h0);
  reg [(2'h2):(1'h0)] reg313 = (1'h0);
  reg [(4'h9):(1'h0)] reg312 = (1'h0);
  reg [(4'h9):(1'h0)] reg310 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg309 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg308 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg307 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg306 = (1'h0);
  reg [(4'h9):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg303 = (1'h0);
  reg [(4'hc):(1'h0)] reg302 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg301 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg298 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg297 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg285 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg280 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg294 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg293 = (1'h0);
  reg [(4'hb):(1'h0)] reg292 = (1'h0);
  reg [(4'hf):(1'h0)] reg291 = (1'h0);
  reg [(2'h3):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg289 = (1'h0);
  reg [(4'hd):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg287 = (1'h0);
  reg signed [(4'he):(1'h0)] reg286 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg284 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg283 = (1'h0);
  reg [(4'ha):(1'h0)] reg282 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg281 = (1'h0);
  reg [(3'h5):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg273 = (1'h0);
  reg [(4'hc):(1'h0)] reg270 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg277 = (1'h0);
  reg [(3'h5):(1'h0)] reg276 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg275 = (1'h0);
  reg [(3'h7):(1'h0)] reg274 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg272 = (1'h0);
  reg [(4'h8):(1'h0)] reg271 = (1'h0);
  reg [(4'hf):(1'h0)] reg254 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg252 = (1'h0);
  reg [(4'h9):(1'h0)] reg247 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg263 = (1'h0);
  reg [(4'hc):(1'h0)] reg262 = (1'h0);
  reg [(4'hf):(1'h0)] reg261 = (1'h0);
  reg [(5'h10):(1'h0)] reg260 = (1'h0);
  reg [(4'h9):(1'h0)] reg259 = (1'h0);
  reg signed [(4'he):(1'h0)] reg258 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg257 = (1'h0);
  reg [(5'h10):(1'h0)] reg256 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg255 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg253 = (1'h0);
  reg [(4'he):(1'h0)] reg251 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg250 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg249 = (1'h0);
  reg [(3'h6):(1'h0)] reg248 = (1'h0);
  reg [(4'hf):(1'h0)] reg246 = (1'h0);
  reg [(4'hb):(1'h0)] reg245 = (1'h0);
  reg [(5'h10):(1'h0)] reg244 = (1'h0);
  reg [(4'hb):(1'h0)] reg242 = (1'h0);
  reg [(4'h8):(1'h0)] reg240 = (1'h0);
  reg [(4'hc):(1'h0)] reg234 = (1'h0);
  reg [(2'h3):(1'h0)] reg233 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg241 = (1'h0);
  reg [(2'h2):(1'h0)] reg239 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg238 = (1'h0);
  reg [(3'h6):(1'h0)] reg237 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg236 = (1'h0);
  reg [(2'h3):(1'h0)] reg235 = (1'h0);
  reg [(4'h8):(1'h0)] reg231 = (1'h0);
  reg [(2'h2):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg227 = (1'h0);
  reg [(4'hf):(1'h0)] reg226 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg221 = (1'h0);
  reg [(2'h3):(1'h0)] reg219 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg215 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg225 = (1'h0);
  reg [(4'hf):(1'h0)] reg224 = (1'h0);
  reg [(4'he):(1'h0)] reg223 = (1'h0);
  reg [(3'h7):(1'h0)] reg222 = (1'h0);
  reg [(3'h7):(1'h0)] reg220 = (1'h0);
  reg [(5'h10):(1'h0)] reg218 = (1'h0);
  reg [(5'h10):(1'h0)] reg217 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg216 = (1'h0);
  reg [(4'hf):(1'h0)] reg214 = (1'h0);
  reg [(4'hb):(1'h0)] reg203 = (1'h0);
  reg [(2'h3):(1'h0)] reg213 = (1'h0);
  reg [(4'h9):(1'h0)] reg212 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg210 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg209 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg208 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg207 = (1'h0);
  reg [(4'hf):(1'h0)] reg206 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg205 = (1'h0);
  reg signed [(4'he):(1'h0)] reg204 = (1'h0);
  reg [(4'hb):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg198 = (1'h0);
  reg [(4'h9):(1'h0)] reg197 = (1'h0);
  reg [(5'h10):(1'h0)] reg196 = (1'h0);
  reg [(4'h9):(1'h0)] reg195 = (1'h0);
  reg signed [(4'he):(1'h0)] reg193 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg191 = (1'h0);
  reg [(3'h4):(1'h0)] reg190 = (1'h0);
  reg [(4'hb):(1'h0)] reg189 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg188 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg186 = (1'h0);
  reg [(4'h9):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg184 = (1'h0);
  reg [(4'hc):(1'h0)] reg182 = (1'h0);
  reg [(3'h7):(1'h0)] reg181 = (1'h0);
  reg signed [(4'he):(1'h0)] reg174 = (1'h0);
  reg [(4'hd):(1'h0)] reg167 = (1'h0);
  reg [(2'h3):(1'h0)] reg180 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg179 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg178 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg177 = (1'h0);
  reg [(4'hd):(1'h0)] reg176 = (1'h0);
  reg [(4'hc):(1'h0)] reg175 = (1'h0);
  reg [(5'h10):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg172 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg171 = (1'h0);
  reg [(4'hc):(1'h0)] reg170 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg169 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg168 = (1'h0);
  reg [(3'h5):(1'h0)] reg165 = (1'h0);
  reg [(4'he):(1'h0)] reg164 = (1'h0);
  reg [(4'hc):(1'h0)] reg163 = (1'h0);
  reg [(4'ha):(1'h0)] reg162 = (1'h0);
  reg [(5'h10):(1'h0)] reg153 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg160 = (1'h0);
  reg [(3'h7):(1'h0)] reg159 = (1'h0);
  reg [(4'he):(1'h0)] reg158 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg156 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg155 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg154 = (1'h0);
  reg [(5'h10):(1'h0)] reg152 = (1'h0);
  reg [(4'hb):(1'h0)] reg151 = (1'h0);
  reg [(2'h2):(1'h0)] reg149 = (1'h0);
  reg [(4'hb):(1'h0)] reg148 = (1'h0);
  reg [(2'h2):(1'h0)] reg147 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg144 = (1'h0);
  reg [(4'ha):(1'h0)] reg143 = (1'h0);
  reg [(5'h10):(1'h0)] reg142 = (1'h0);
  reg [(4'ha):(1'h0)] reg141 = (1'h0);
  reg [(3'h4):(1'h0)] reg140 = (1'h0);
  reg [(4'hf):(1'h0)] reg139 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg136 = (1'h0);
  reg [(3'h6):(1'h0)] reg134 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg133 = (1'h0);
  reg signed [(4'he):(1'h0)] reg132 = (1'h0);
  reg [(4'hf):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg130 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg129 = (1'h0);
  reg signed [(4'he):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg126 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg125 = (1'h0);
  reg [(4'h8):(1'h0)] reg124 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg123 = (1'h0);
  reg [(3'h7):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg121 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg120 = (1'h0);
  reg [(5'h10):(1'h0)] reg118 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg117 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg115 = (1'h0);
  reg [(3'h4):(1'h0)] reg114 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg113 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg112 = (1'h0);
  reg [(4'hd):(1'h0)] reg100 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg96 = (1'h0);
  reg [(4'ha):(1'h0)] reg109 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg107 = (1'h0);
  reg [(4'h8):(1'h0)] reg106 = (1'h0);
  reg signed [(4'he):(1'h0)] reg104 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg101 = (1'h0);
  reg [(3'h6):(1'h0)] reg99 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg98 = (1'h0);
  reg [(4'h9):(1'h0)] reg97 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg95 = (1'h0);
  reg [(2'h2):(1'h0)] reg94 = (1'h0);
  reg [(4'hd):(1'h0)] reg90 = (1'h0);
  reg signed [(4'he):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg88 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg84 = (1'h0);
  reg [(3'h6):(1'h0)] reg83 = (1'h0);
  reg [(4'ha):(1'h0)] reg82 = (1'h0);
  reg [(3'h4):(1'h0)] reg81 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg77 = (1'h0);
  reg signed [(4'he):(1'h0)] reg76 = (1'h0);
  reg [(4'hb):(1'h0)] reg75 = (1'h0);
  reg [(5'h10):(1'h0)] reg73 = (1'h0);
  reg [(3'h5):(1'h0)] reg69 = (1'h0);
  reg [(2'h2):(1'h0)] reg66 = (1'h0);
  reg [(4'hd):(1'h0)] reg72 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg71 = (1'h0);
  reg [(5'h10):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg67 = (1'h0);
  reg [(2'h2):(1'h0)] reg65 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg64 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg63 = (1'h0);
  reg [(4'ha):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg52 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg58 = (1'h0);
  reg [(3'h4):(1'h0)] reg62 = (1'h0);
  reg [(4'he):(1'h0)] reg61 = (1'h0);
  reg [(4'hd):(1'h0)] reg59 = (1'h0);
  reg [(4'h9):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg56 = (1'h0);
  reg [(3'h6):(1'h0)] reg44 = (1'h0);
  reg signed [(4'he):(1'h0)] reg54 = (1'h0);
  reg [(4'hd):(1'h0)] reg53 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg51 = (1'h0);
  reg [(4'hd):(1'h0)] reg50 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg49 = (1'h0);
  reg [(3'h4):(1'h0)] reg48 = (1'h0);
  reg [(3'h7):(1'h0)] reg46 = (1'h0);
  reg [(4'ha):(1'h0)] reg45 = (1'h0);
  reg [(4'ha):(1'h0)] reg43 = (1'h0);
  reg [(2'h2):(1'h0)] reg42 = (1'h0);
  reg [(5'h10):(1'h0)] reg41 = (1'h0);
  reg [(3'h7):(1'h0)] reg40 = (1'h0);
  reg [(4'h9):(1'h0)] reg39 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg37 = (1'h0);
  reg [(4'h8):(1'h0)] reg36 = (1'h0);
  reg signed [(4'he):(1'h0)] reg35 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg33 = (1'h0);
  reg [(2'h3):(1'h0)] reg32 = (1'h0);
  reg [(5'h10):(1'h0)] reg31 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg30 = (1'h0);
  reg [(4'hd):(1'h0)] reg29 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg28 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg27 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg26 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg23 = (1'h0);
  reg [(4'hb):(1'h0)] reg22 = (1'h0);
  reg [(4'hd):(1'h0)] reg20 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg18 = (1'h0);
  reg [(5'h10):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg16 = (1'h0);
  reg [(2'h3):(1'h0)] forvar623 = (1'h0);
  reg [(3'h5):(1'h0)] forvar619 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar617 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar614 = (1'h0);
  reg [(3'h7):(1'h0)] forvar612 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar610 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar609 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar605 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar598 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar596 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar594 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar593 = (1'h0);
  reg [(2'h2):(1'h0)] forvar588 = (1'h0);
  reg [(2'h2):(1'h0)] forvar575 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar565 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar561 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar554 = (1'h0);
  reg [(4'hb):(1'h0)] forvar546 = (1'h0);
  reg [(4'he):(1'h0)] forvar541 = (1'h0);
  reg [(3'h6):(1'h0)] forvar587 = (1'h0);
  reg [(4'h9):(1'h0)] forvar582 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar577 = (1'h0);
  reg [(4'hd):(1'h0)] forvar572 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar567 = (1'h0);
  reg [(4'ha):(1'h0)] forvar564 = (1'h0);
  reg [(4'hd):(1'h0)] forvar559 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar551 = (1'h0);
  reg [(5'h10):(1'h0)] forvar550 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar542 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar540 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar539 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar379 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar365 = (1'h0);
  reg [(5'h10):(1'h0)] forvar378 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar376 = (1'h0);
  reg [(4'he):(1'h0)] forvar375 = (1'h0);
  reg [(2'h3):(1'h0)] forvar370 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar366 = (1'h0);
  reg [(4'he):(1'h0)] forvar364 = (1'h0);
  reg [(3'h6):(1'h0)] forvar361 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar346 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar344 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar340 = (1'h0);
  reg [(3'h5):(1'h0)] forvar326 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar317 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar356 = (1'h0);
  reg [(4'ha):(1'h0)] forvar354 = (1'h0);
  reg [(2'h3):(1'h0)] forvar350 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar348 = (1'h0);
  reg [(3'h5):(1'h0)] forvar343 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar341 = (1'h0);
  reg [(4'hc):(1'h0)] forvar336 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar335 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar333 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar329 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar321 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar320 = (1'h0);
  reg [(4'hf):(1'h0)] forvar318 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar310 = (1'h0);
  reg [(2'h3):(1'h0)] forvar314 = (1'h0);
  reg [(2'h2):(1'h0)] forvar311 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar304 = (1'h0);
  reg [(4'hc):(1'h0)] forvar300 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar299 = (1'h0);
  reg [(4'h9):(1'h0)] forvar296 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar295 = (1'h0);
  reg [(3'h5):(1'h0)] forvar290 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar286 = (1'h0);
  reg [(4'hc):(1'h0)] forvar277 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar292 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar285 = (1'h0);
  reg [(4'h8):(1'h0)] forvar280 = (1'h0);
  reg [(5'h10):(1'h0)] forvar279 = (1'h0);
  reg [(4'he):(1'h0)] forvar271 = (1'h0);
  reg [(2'h3):(1'h0)] forvar273 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar270 = (1'h0);
  reg [(4'h9):(1'h0)] forvar269 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar249 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar248 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar254 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar252 = (1'h0);
  reg [(3'h5):(1'h0)] forvar247 = (1'h0);
  reg [(5'h10):(1'h0)] forvar243 = (1'h0);
  reg [(4'hb):(1'h0)] forvar241 = (1'h0);
  reg [(4'he):(1'h0)] forvar237 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar240 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar234 = (1'h0);
  reg [(4'h9):(1'h0)] forvar233 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar232 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar229 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar228 = (1'h0);
  reg [(4'h8):(1'h0)] forvar220 = (1'h0);
  reg [(4'hf):(1'h0)] forvar214 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar221 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar219 = (1'h0);
  reg [(4'hb):(1'h0)] forvar215 = (1'h0);
  reg [(4'h9):(1'h0)] forvar208 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar203 = (1'h0);
  reg [(4'ha):(1'h0)] forvar202 = (1'h0);
  reg [(3'h7):(1'h0)] forvar201 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar199 = (1'h0);
  reg [(4'hb):(1'h0)] forvar194 = (1'h0);
  reg [(3'h7):(1'h0)] forvar192 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar187 = (1'h0);
  reg [(4'hd):(1'h0)] forvar183 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar178 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar177 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar176 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar171 = (1'h0);
  reg [(5'h10):(1'h0)] forvar170 = (1'h0);
  reg [(2'h3):(1'h0)] forvar168 = (1'h0);
  reg [(3'h5):(1'h0)] forvar174 = (1'h0);
  reg [(3'h4):(1'h0)] forvar167 = (1'h0);
  reg [(3'h4):(1'h0)] forvar166 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar161 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar157 = (1'h0);
  reg [(4'h9):(1'h0)] forvar153 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar150 = (1'h0);
  reg [(4'hd):(1'h0)] forvar146 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar145 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar138 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar137 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar135 = (1'h0);
  reg [(4'h9):(1'h0)] forvar130 = (1'h0);
  reg [(3'h6):(1'h0)] forvar128 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar127 = (1'h0);
  reg [(4'hd):(1'h0)] forvar122 = (1'h0);
  reg [(4'hd):(1'h0)] forvar117 = (1'h0);
  reg [(3'h4):(1'h0)] forvar119 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar116 = (1'h0);
  reg [(4'h8):(1'h0)] forvar111 = (1'h0);
  reg [(3'h6):(1'h0)] forvar110 = (1'h0);
  reg [(3'h6):(1'h0)] forvar99 = (1'h0);
  reg [(3'h6):(1'h0)] forvar108 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar105 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar100 = (1'h0);
  reg [(3'h4):(1'h0)] forvar96 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar93 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar92 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar89 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar90 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar87 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar86 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar80 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar79 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar74 = (1'h0);
  reg [(3'h7):(1'h0)] forvar65 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar69 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar66 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar54 = (1'h0);
  reg [(4'h9):(1'h0)] forvar42 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar60 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar58 = (1'h0);
  reg [(3'h6):(1'h0)] forvar55 = (1'h0);
  reg [(4'h8):(1'h0)] forvar45 = (1'h0);
  reg [(4'h8):(1'h0)] forvar52 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar47 = (1'h0);
  reg [(4'he):(1'h0)] forvar44 = (1'h0);
  reg [(4'h8):(1'h0)] forvar38 = (1'h0);
  reg [(4'hb):(1'h0)] forvar34 = (1'h0);
  reg [(3'h5):(1'h0)] forvar32 = (1'h0);
  reg [(2'h2):(1'h0)] forvar25 = (1'h0);
  reg [(4'hb):(1'h0)] forvar21 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar15 = (1'h0);
  reg [(4'hc):(1'h0)] forvar14 = (1'h0);
  reg [(3'h4):(1'h0)] forvar13 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar12 = (1'h0);
  assign y = {wire627,
                 wire535,
                 wire268,
                 wire267,
                 wire266,
                 wire265,
                 wire11,
                 reg626,
                 reg625,
                 reg624,
                 reg622,
                 reg621,
                 reg620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 reg615,
                 reg613,
                 reg611,
                 reg608,
                 reg607,
                 reg606,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 reg597,
                 reg595,
                 reg592,
                 reg587,
                 reg582,
                 reg572,
                 reg567,
                 reg551,
                 reg542,
                 reg540,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg581,
                 reg580,
                 reg579,
                 reg578,
                 reg576,
                 reg575,
                 reg574,
                 reg573,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 reg566,
                 reg565,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 reg549,
                 reg548,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 reg543,
                 reg541,
                 reg538,
                 reg537,
                 reg384,
                 reg383,
                 reg378,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg377,
                 reg374,
                 reg370,
                 reg366,
                 reg373,
                 reg372,
                 reg371,
                 reg369,
                 reg368,
                 reg367,
                 reg365,
                 reg363,
                 reg362,
                 reg348,
                 reg343,
                 reg341,
                 reg336,
                 reg335,
                 reg333,
                 reg329,
                 reg318,
                 reg321,
                 reg320,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg342,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg334,
                 reg332,
                 reg331,
                 reg330,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg319,
                 reg317,
                 reg314,
                 reg311,
                 reg299,
                 reg300,
                 reg316,
                 reg315,
                 reg313,
                 reg312,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg303,
                 reg302,
                 reg301,
                 reg298,
                 reg297,
                 reg285,
                 reg280,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg278,
                 reg273,
                 reg270,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg272,
                 reg271,
                 reg254,
                 reg252,
                 reg247,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg253,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg246,
                 reg245,
                 reg244,
                 reg242,
                 reg240,
                 reg234,
                 reg233,
                 reg241,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg231,
                 reg230,
                 reg227,
                 reg226,
                 reg221,
                 reg219,
                 reg215,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg220,
                 reg218,
                 reg217,
                 reg216,
                 reg214,
                 reg203,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg200,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg193,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg186,
                 reg185,
                 reg184,
                 reg182,
                 reg181,
                 reg174,
                 reg167,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg153,
                 reg160,
                 reg159,
                 reg158,
                 reg156,
                 reg155,
                 reg154,
                 reg152,
                 reg151,
                 reg149,
                 reg148,
                 reg147,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg136,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg118,
                 reg117,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg100,
                 reg96,
                 reg109,
                 reg107,
                 reg106,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg99,
                 reg98,
                 reg97,
                 reg95,
                 reg94,
                 reg90,
                 reg91,
                 reg89,
                 reg88,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg73,
                 reg69,
                 reg66,
                 reg72,
                 reg71,
                 reg70,
                 reg68,
                 reg67,
                 reg65,
                 reg64,
                 reg63,
                 reg55,
                 reg52,
                 reg58,
                 reg62,
                 reg61,
                 reg59,
                 reg57,
                 reg56,
                 reg44,
                 reg54,
                 reg53,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg46,
                 reg45,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg37,
                 reg36,
                 reg35,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg24,
                 reg23,
                 reg22,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 forvar623,
                 forvar619,
                 forvar617,
                 forvar614,
                 forvar612,
                 forvar610,
                 forvar609,
                 forvar605,
                 forvar598,
                 forvar596,
                 forvar594,
                 forvar593,
                 forvar588,
                 forvar575,
                 forvar565,
                 forvar561,
                 forvar554,
                 forvar546,
                 forvar541,
                 forvar587,
                 forvar582,
                 forvar577,
                 forvar572,
                 forvar567,
                 forvar564,
                 forvar559,
                 forvar551,
                 forvar550,
                 forvar542,
                 forvar540,
                 forvar539,
                 forvar379,
                 forvar365,
                 forvar378,
                 forvar376,
                 forvar375,
                 forvar370,
                 forvar366,
                 forvar364,
                 forvar361,
                 forvar346,
                 forvar344,
                 forvar340,
                 forvar326,
                 forvar317,
                 forvar356,
                 forvar354,
                 forvar350,
                 forvar348,
                 forvar343,
                 forvar341,
                 forvar336,
                 forvar335,
                 forvar333,
                 forvar329,
                 forvar321,
                 forvar320,
                 forvar318,
                 forvar310,
                 forvar314,
                 forvar311,
                 forvar304,
                 forvar300,
                 forvar299,
                 forvar296,
                 forvar295,
                 forvar290,
                 forvar286,
                 forvar277,
                 forvar292,
                 forvar285,
                 forvar280,
                 forvar279,
                 forvar271,
                 forvar273,
                 forvar270,
                 forvar269,
                 forvar249,
                 forvar248,
                 forvar254,
                 forvar252,
                 forvar247,
                 forvar243,
                 forvar241,
                 forvar237,
                 forvar240,
                 forvar234,
                 forvar233,
                 forvar232,
                 forvar229,
                 forvar228,
                 forvar220,
                 forvar214,
                 forvar221,
                 forvar219,
                 forvar215,
                 forvar208,
                 forvar203,
                 forvar202,
                 forvar201,
                 forvar199,
                 forvar194,
                 forvar192,
                 forvar187,
                 forvar183,
                 forvar178,
                 forvar177,
                 forvar176,
                 forvar171,
                 forvar170,
                 forvar168,
                 forvar174,
                 forvar167,
                 forvar166,
                 forvar161,
                 forvar157,
                 forvar153,
                 forvar150,
                 forvar146,
                 forvar145,
                 forvar138,
                 forvar137,
                 forvar135,
                 forvar130,
                 forvar128,
                 forvar127,
                 forvar122,
                 forvar117,
                 forvar119,
                 forvar116,
                 forvar111,
                 forvar110,
                 forvar99,
                 forvar108,
                 forvar105,
                 forvar100,
                 forvar96,
                 forvar93,
                 forvar92,
                 forvar89,
                 forvar90,
                 forvar87,
                 forvar86,
                 forvar80,
                 forvar79,
                 forvar74,
                 forvar65,
                 forvar69,
                 forvar66,
                 forvar54,
                 forvar42,
                 forvar60,
                 forvar58,
                 forvar55,
                 forvar45,
                 forvar52,
                 forvar47,
                 forvar44,
                 forvar38,
                 forvar34,
                 forvar32,
                 forvar25,
                 forvar21,
                 forvar15,
                 forvar14,
                 forvar13,
                 forvar12,
                 (1'h0)};
  assign wire11 = $signed(((~wire7) ?
                      wire9[(3'h4):(3'h4)] : {(wire7 ? wire10 : wire9)}));
  always
    @(posedge clk) begin
      for (forvar12 = (1'h0); (forvar12 < (2'h2)); forvar12 = (forvar12 + (1'h1)))
        begin
          for (forvar13 = (1'h0); (forvar13 < (2'h2)); forvar13 = (forvar13 + (1'h1)))
            begin
              for (forvar14 = (1'h0); (forvar14 < (2'h3)); forvar14 = (forvar14 + (1'h1)))
                begin
                  for (forvar15 = (1'h0); (forvar15 < (2'h2)); forvar15 = (forvar15 + (1'h1)))
                    begin
                      reg16 <= (-forvar14[(4'h9):(2'h3)]);
                      reg17 <= $unsigned((-$unsigned((+wire9))));
                      reg18 <= forvar14[(2'h2):(1'h1)];
                      reg19 <= wire11;
                    end
                  reg20 <= $signed((((wire11 ^~ reg18) ?
                      wire7 : reg17[(4'hf):(3'h7)]) && wire9));
                  for (forvar21 = (1'h0); (forvar21 < (1'h0)); forvar21 = (forvar21 + (1'h1)))
                    begin
                      reg22 <= reg16;
                      reg23 <= (&(reg17 != wire9));
                      reg24 <= (reg22[(3'h7):(1'h1)] ?
                          forvar14[(4'h8):(2'h2)] : wire8[(3'h4):(1'h0)]);
                    end
                  for (forvar25 = (1'h0); (forvar25 < (2'h2)); forvar25 = (forvar25 + (1'h1)))
                    begin
                      reg26 <= ((+$unsigned((reg19 * reg19))) ?
                          $unsigned((-reg23)) : wire8);
                      reg27 <= reg18[(1'h0):(1'h0)];
                      reg28 <= {forvar13[(2'h2):(1'h1)]};
                      reg29 <= $signed($unsigned({wire11}));
                    end
                end
              if (forvar12[(4'h9):(4'h8)])
                begin
                  reg30 <= (((((8'ha8) ? (8'hb5) : forvar15) >>> reg18) ?
                      {(reg18 && forvar12)} : wire6) ~^ reg26[(4'h8):(3'h4)]);
                  if ($unsigned((reg16 ? reg29[(3'h7):(1'h0)] : (8'haa))))
                    begin
                      reg31 <= ((-reg30[(4'ha):(3'h7)]) <= {$unsigned($unsigned(reg28))});
                      reg32 <= $signed({(reg22 ^~ reg28)});
                      reg33 <= {{wire8}};
                    end
                  else
                    begin
                      reg31 <= (~|{(^reg26)});
                      reg32 <= reg30[(1'h1):(1'h1)];
                      reg33 <= $signed(((forvar14 ?
                          (wire6 && reg22) : (reg19 ?
                              (8'haf) : forvar25)) - (forvar21 | reg16)));
                    end
                end
              else
                begin
                  if (forvar15)
                    begin
                      reg30 <= $unsigned($signed(reg20));
                    end
                  else
                    begin
                      reg30 <= {reg23[(3'h7):(1'h0)]};
                      reg31 <= (8'had);
                    end
                  for (forvar32 = (1'h0); (forvar32 < (2'h3)); forvar32 = (forvar32 + (1'h1)))
                    begin
                      reg33 <= ($unsigned({{reg30}}) & (^forvar14));
                    end
                  for (forvar34 = (1'h0); (forvar34 < (2'h2)); forvar34 = (forvar34 + (1'h1)))
                    begin
                      reg35 <= $unsigned(reg29[(2'h3):(2'h2)]);
                      reg36 <= ({(~^$signed((8'haa)))} + (&$unsigned((reg32 ~^ reg17))));
                      reg37 <= $unsigned((&(~^wire8)));
                    end
                  for (forvar38 = (1'h0); (forvar38 < (1'h0)); forvar38 = (forvar38 + (1'h1)))
                    begin
                      reg39 <= (($unsigned(wire10) ? reg27 : {{reg35}}) ?
                          forvar34[(4'h8):(3'h6)] : forvar14);
                      reg40 <= (((-(+reg22)) << $unsigned($unsigned((8'haa)))) ?
                          (!($unsigned(reg32) ?
                              reg20[(3'h7):(1'h1)] : $signed(reg28))) : $signed(forvar14[(3'h5):(2'h3)]));
                      reg41 <= $unsigned((~&wire11));
                    end
                end
            end
          if (reg27)
            begin
              reg42 <= $unsigned($signed(((forvar25 | forvar25) >>> (^forvar13))));
              reg43 <= (^~(((+(8'ha6)) <<< (|forvar25)) || {(~&reg39)}));
              if ({reg28})
                begin
                  for (forvar44 = (1'h0); (forvar44 < (2'h2)); forvar44 = (forvar44 + (1'h1)))
                    begin
                      reg45 <= (^~(8'ha9));
                      reg46 <= {$signed(reg40[(2'h3):(1'h0)])};
                    end
                  for (forvar47 = (1'h0); (forvar47 < (1'h1)); forvar47 = (forvar47 + (1'h1)))
                    begin
                      reg48 <= $signed((|($signed(wire8) ?
                          {forvar14} : (wire7 - forvar32))));
                      reg49 <= ($signed((8'ha9)) ?
                          reg31[(4'he):(4'h8)] : ({$unsigned(reg22)} ?
                              reg26[(3'h5):(1'h0)] : ($signed(forvar47) ?
                                  $signed((8'hb2)) : (reg30 || wire10))));
                      reg50 <= ((+{(forvar13 > reg42)}) ?
                          $signed(reg16) : $signed($signed((forvar21 >>> wire8))));
                      reg51 <= reg46[(1'h0):(1'h0)];
                    end
                  for (forvar52 = (1'h0); (forvar52 < (2'h2)); forvar52 = (forvar52 + (1'h1)))
                    begin
                      reg53 <= (((|(reg19 ? reg51 : (8'ha6))) ?
                              ((8'hb5) ?
                                  $unsigned((8'ha0)) : {reg36}) : (!(~forvar21))) ?
                          (reg36[(3'h5):(2'h3)] ?
                              (~^(~wire11)) : $signed(reg26[(4'ha):(2'h3)])) : reg29);
                      reg54 <= {reg35};
                    end
                end
              else
                begin
                  reg44 <= wire10[(2'h3):(2'h3)];
                  for (forvar45 = (1'h0); (forvar45 < (1'h0)); forvar45 = (forvar45 + (1'h1)))
                    begin
                      reg46 <= $signed((|(~^$signed((8'had)))));
                    end
                end
              if (reg45)
                begin
                  for (forvar55 = (1'h0); (forvar55 < (2'h3)); forvar55 = (forvar55 + (1'h1)))
                    begin
                      reg56 <= {forvar13[(1'h0):(1'h0)]};
                      reg57 <= $unsigned(((^(forvar13 || reg31)) ?
                          wire11[(2'h3):(2'h2)] : $signed($unsigned(wire8))));
                    end
                  for (forvar58 = (1'h0); (forvar58 < (1'h0)); forvar58 = (forvar58 + (1'h1)))
                    begin
                      reg59 <= forvar21[(3'h5):(2'h2)];
                    end
                  for (forvar60 = (1'h0); (forvar60 < (1'h1)); forvar60 = (forvar60 + (1'h1)))
                    begin
                      reg61 <= forvar34;
                      reg62 <= $unsigned(reg46);
                    end
                end
              else
                begin
                  for (forvar55 = (1'h0); (forvar55 < (1'h1)); forvar55 = (forvar55 + (1'h1)))
                    begin
                      reg56 <= reg17[(4'hf):(3'h7)];
                      reg57 <= {reg57[(3'h4):(3'h4)]};
                      reg58 <= (^~((forvar13 ?
                          (forvar32 ?
                              reg17 : forvar55) : wire9) > ((forvar45 <<< forvar13) ?
                          (reg46 ? reg16 : (8'ha6)) : $unsigned(wire7))));
                      reg59 <= ((forvar15[(2'h2):(1'h1)] ?
                          (~|(wire9 <<< reg48)) : reg48) || $signed((~reg17[(4'he):(1'h0)])));
                    end
                end
            end
          else
            begin
              for (forvar42 = (1'h0); (forvar42 < (2'h3)); forvar42 = (forvar42 + (1'h1)))
                begin
                  if ($unsigned({(((8'hb2) ?
                          forvar12 : reg57) >>> $signed(reg16))}))
                    begin
                      reg43 <= $signed(($signed({forvar44}) & $unsigned($unsigned(reg26))));
                      reg44 <= ((|((reg54 ? reg56 : (8'hb6)) ?
                              (8'haa) : $signed((8'haa)))) ?
                          $signed(($unsigned(reg40) == (reg40 - reg35))) : reg30[(3'h5):(1'h0)]);
                      reg45 <= reg50;
                    end
                  else
                    begin
                      reg43 <= reg59;
                    end
                  reg46 <= reg59[(3'h6):(1'h1)];
                end
              for (forvar47 = (1'h0); (forvar47 < (2'h2)); forvar47 = (forvar47 + (1'h1)))
                begin
                  if (reg48[(1'h0):(1'h0)])
                    begin
                      reg48 <= reg49[(2'h3):(2'h3)];
                      reg49 <= reg54[(4'ha):(2'h3)];
                      reg50 <= reg42;
                    end
                  else
                    begin
                      reg48 <= (forvar21 ?
                          $signed((wire9[(3'h5):(1'h0)] <= reg50)) : reg42);
                      reg49 <= {($unsigned((wire10 <= reg46)) && $signed(reg20[(3'h5):(3'h4)]))};
                      reg50 <= (!$unsigned(wire6));
                    end
                  if ($signed($unsigned({{reg28}})))
                    begin
                      reg51 <= reg44;
                      reg52 <= ($signed(wire10) >>> ($signed((wire9 && reg19)) ?
                          reg27[(4'hc):(2'h3)] : ((~reg53) ?
                              $signed(forvar13) : (8'ha8))));
                      reg53 <= reg49[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg51 <= $unsigned((8'ha9));
                      reg52 <= forvar44[(4'hc):(3'h4)];
                      reg53 <= $signed(forvar45);
                    end
                  for (forvar54 = (1'h0); (forvar54 < (1'h0)); forvar54 = (forvar54 + (1'h1)))
                    begin
                      reg55 <= (+$signed(forvar60));
                      reg56 <= (|(|(((8'haa) ? (8'hb6) : reg58) >>> (reg36 ?
                          reg61 : reg44))));
                    end
                end
            end
          if (($unsigned(($unsigned(reg20) >= wire11)) <<< reg53[(3'h5):(2'h3)]))
            begin
              if (reg31)
                begin
                  if (($unsigned({(+reg40)}) * reg44[(3'h6):(1'h1)]))
                    begin
                      reg63 <= wire11[(1'h1):(1'h1)];
                      reg64 <= ($signed(reg58) & forvar34[(3'h4):(2'h3)]);
                      reg65 <= reg46;
                    end
                  else
                    begin
                      reg63 <= $unsigned($signed((-(forvar38 * reg16))));
                      reg64 <= (^forvar38[(1'h1):(1'h1)]);
                      reg65 <= (~|reg40[(3'h5):(3'h4)]);
                    end
                  for (forvar66 = (1'h0); (forvar66 < (2'h3)); forvar66 = (forvar66 + (1'h1)))
                    begin
                      reg67 <= $signed($signed($unsigned((~reg52))));
                      reg68 <= $unsigned(((&reg37[(3'h5):(3'h4)]) ?
                          forvar38 : ((~&reg54) >> $unsigned(reg63))));
                    end
                  for (forvar69 = (1'h0); (forvar69 < (2'h3)); forvar69 = (forvar69 + (1'h1)))
                    begin
                      reg70 <= reg32[(1'h1):(1'h1)];
                      reg71 <= reg54;
                      reg72 <= (8'haa);
                    end
                end
              else
                begin
                  if ((&(($signed(reg44) ? {reg58} : forvar45[(1'h0):(1'h0)]) ?
                      {$signed((8'hb5))} : (reg33 - {reg37}))))
                    begin
                      reg63 <= (((&{reg27}) <= (8'haa)) ?
                          reg24 : $signed(reg28));
                    end
                  else
                    begin
                      reg63 <= reg42[(1'h0):(1'h0)];
                    end
                  reg64 <= ((reg18 << ($unsigned(reg36) - {reg64})) == $unsigned((~(&forvar69))));
                  for (forvar65 = (1'h0); (forvar65 < (1'h1)); forvar65 = (forvar65 + (1'h1)))
                    begin
                      reg66 <= $signed(((&$unsigned(reg67)) ?
                          reg63 : ($signed(reg20) ?
                              $unsigned(reg24) : {(8'ha8)})));
                    end
                  if (($signed(forvar44) ?
                      ((-(~^forvar69)) ?
                          ($signed(reg41) != $unsigned(forvar65)) : (((8'hb9) ^~ reg40) ?
                              forvar47 : (~|reg24))) : reg36[(1'h0):(1'h0)]))
                    begin
                      reg67 <= $unsigned(forvar32[(1'h0):(1'h0)]);
                      reg68 <= ((~&reg18) != {wire11[(2'h2):(1'h1)]});
                      reg69 <= $signed(reg42);
                      reg70 <= $signed(forvar47);
                    end
                  else
                    begin
                      reg67 <= (forvar34 <<< $unsigned(($unsigned(reg40) ?
                          $unsigned(reg54) : $unsigned(forvar12))));
                      reg68 <= (!$unsigned($unsigned($signed(reg17))));
                      reg69 <= ($signed((reg35[(4'hd):(3'h7)] ?
                          ((8'ha7) + reg72) : (reg45 & reg58))) >>> reg65);
                    end
                end
            end
          else
            begin
              reg63 <= reg48;
              reg64 <= reg68;
              if (((~|$signed($signed(reg24))) ^~ ($signed((+reg52)) ^ $unsigned((reg40 <<< reg56)))))
                begin
                  for (forvar65 = (1'h0); (forvar65 < (2'h2)); forvar65 = (forvar65 + (1'h1)))
                    begin
                      reg66 <= ($unsigned(($unsigned(reg57) ?
                              reg24 : $signed(reg31))) ?
                          $unsigned(reg18[(3'h6):(1'h0)]) : (&(reg30 & $signed(reg30))));
                      reg67 <= (reg29[(4'ha):(1'h0)] ?
                          forvar55[(2'h3):(2'h3)] : (reg63[(3'h4):(2'h2)] ?
                              ($signed((8'hb2)) ?
                                  (+forvar47) : ((8'ha7) ?
                                      reg66 : reg32)) : {reg50[(2'h2):(1'h0)]}));
                    end
                end
              else
                begin
                  for (forvar65 = (1'h0); (forvar65 < (1'h0)); forvar65 = (forvar65 + (1'h1)))
                    begin
                      reg66 <= $unsigned(((|(reg52 ?
                          reg72 : reg53)) ~^ $signed($unsigned(wire11))));
                      reg67 <= forvar47[(2'h2):(1'h0)];
                      reg68 <= {$signed(((forvar47 > (8'hb4)) ?
                              (reg71 << (8'hac)) : reg63))};
                    end
                  for (forvar69 = (1'h0); (forvar69 < (1'h0)); forvar69 = (forvar69 + (1'h1)))
                    begin
                      reg70 <= $unsigned({$unsigned(((8'ha2) ?
                              (8'hb2) : forvar32))});
                      reg71 <= forvar45[(3'h6):(1'h0)];
                      reg72 <= $signed((reg57 ?
                          ($unsigned(forvar14) ?
                              reg59 : wire11) : (-(~(8'hac)))));
                      reg73 <= $unsigned(($unsigned((^forvar42)) ?
                          (!forvar14[(4'ha):(3'h4)]) : $signed(((8'h9f) ?
                              reg32 : forvar54))));
                    end
                  for (forvar74 = (1'h0); (forvar74 < (2'h3)); forvar74 = (forvar74 + (1'h1)))
                    begin
                      reg75 <= $unsigned($unsigned(($unsigned(forvar45) ?
                          (^reg69) : (forvar47 ? forvar47 : reg72))));
                      reg76 <= forvar14;
                      reg77 <= $signed(({wire9} ?
                          (~^$signed(forvar21)) : reg65[(2'h2):(1'h0)]));
                    end
                  reg78 <= ((!(reg77[(3'h4):(1'h0)] + $unsigned(reg51))) == ($unsigned($signed(reg39)) ?
                      {$signed(reg66)} : reg73));
                end
            end
          for (forvar79 = (1'h0); (forvar79 < (2'h3)); forvar79 = (forvar79 + (1'h1)))
            begin
              for (forvar80 = (1'h0); (forvar80 < (1'h1)); forvar80 = (forvar80 + (1'h1)))
                begin
                  if ($signed((|forvar65)))
                    begin
                      reg81 <= (^$signed(((|wire6) ?
                          ((8'ha8) >> forvar15) : reg71)));
                      reg82 <= $signed(reg45);
                      reg83 <= ($unsigned((8'haf)) ?
                          ($signed(reg32[(1'h0):(1'h0)]) << $signed($unsigned(reg66))) : (^((forvar38 + reg81) ?
                              {forvar13} : reg58)));
                      reg84 <= reg57[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg81 <= (^{(reg39 - $unsigned(forvar65))});
                    end
                  reg85 <= $signed($signed(($unsigned(forvar12) ^ reg44[(3'h5):(2'h2)])));
                end
            end
        end
      for (forvar86 = (1'h0); (forvar86 < (1'h1)); forvar86 = (forvar86 + (1'h1)))
        begin
          for (forvar87 = (1'h0); (forvar87 < (2'h3)); forvar87 = (forvar87 + (1'h1)))
            begin
              reg88 <= (8'ha0);
              if (($unsigned(reg22) || (({reg88} || reg83) ?
                  $signed($signed(reg76)) : $unsigned((^reg75)))))
                begin
                  reg89 <= $unsigned(wire7[(3'h4):(1'h0)]);
                  for (forvar90 = (1'h0); (forvar90 < (2'h2)); forvar90 = (forvar90 + (1'h1)))
                    begin
                      reg91 <= (&(8'hb1));
                    end
                end
              else
                begin
                  for (forvar89 = (1'h0); (forvar89 < (2'h3)); forvar89 = (forvar89 + (1'h1)))
                    begin
                      reg90 <= (8'hb1);
                      reg91 <= $unsigned(reg72);
                    end
                end
              for (forvar92 = (1'h0); (forvar92 < (2'h3)); forvar92 = (forvar92 + (1'h1)))
                begin
                  for (forvar93 = (1'h0); (forvar93 < (1'h0)); forvar93 = (forvar93 + (1'h1)))
                    begin
                      reg94 <= $signed(reg53[(4'hd):(2'h3)]);
                      reg95 <= reg46;
                    end
                end
              if (forvar47[(3'h4):(2'h3)])
                begin
                  for (forvar96 = (1'h0); (forvar96 < (2'h3)); forvar96 = (forvar96 + (1'h1)))
                    begin
                      reg97 <= $signed((-$unsigned((reg88 ? reg51 : reg37))));
                      reg98 <= (($signed((!(8'hae))) <= {(reg19 ?
                              wire11 : (8'hb2))}) > {wire11});
                      reg99 <= reg31;
                    end
                  for (forvar100 = (1'h0); (forvar100 < (1'h0)); forvar100 = (forvar100 + (1'h1)))
                    begin
                      reg101 <= $signed({reg43[(3'h5):(2'h2)]});
                      reg102 <= $unsigned(($signed((8'ha8)) == $signed($unsigned(reg91))));
                      reg103 <= reg59;
                      reg104 <= $signed(((reg54 ?
                              (reg57 > reg44) : (forvar54 > reg39)) ?
                          reg85[(3'h5):(2'h2)] : (-$signed(reg98))));
                    end
                  for (forvar105 = (1'h0); (forvar105 < (2'h3)); forvar105 = (forvar105 + (1'h1)))
                    begin
                      reg106 <= (($unsigned((reg40 <<< forvar100)) ^ $signed($signed(reg41))) - (-(&(wire8 ?
                          reg27 : reg63))));
                      reg107 <= ((+wire9) ? reg57 : $signed(wire10));
                    end
                  for (forvar108 = (1'h0); (forvar108 < (1'h1)); forvar108 = (forvar108 + (1'h1)))
                    begin
                      reg109 <= (forvar32[(2'h3):(2'h3)] ^ (((reg89 ?
                          (8'ha1) : (8'h9d)) == (+reg68)) > (forvar47 < reg19)));
                    end
                end
              else
                begin
                  if ($unsigned((((reg29 <= reg53) + {reg63}) >>> $unsigned((reg109 - forvar44)))))
                    begin
                      reg96 <= $unsigned({{reg23}});
                      reg97 <= (&(((^~reg84) <<< $unsigned(forvar100)) < $unsigned((reg70 ?
                          wire8 : wire7))));
                      reg98 <= forvar100[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg96 <= (forvar89[(1'h0):(1'h0)] ?
                          {$unsigned((forvar74 ?
                                  forvar45 : reg18))} : $unsigned(reg102[(3'h6):(3'h6)]));
                      reg97 <= $signed(reg53[(4'hc):(4'h9)]);
                    end
                  for (forvar99 = (1'h0); (forvar99 < (2'h3)); forvar99 = (forvar99 + (1'h1)))
                    begin
                      reg100 <= (reg35 == $unsigned($unsigned(reg69)));
                    end
                  reg101 <= forvar21[(4'h8):(1'h0)];
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar110 = (1'h0); (forvar110 < (2'h2)); forvar110 = (forvar110 + (1'h1)))
        begin
          if ($unsigned(((|(reg32 ? reg56 : reg53)) ~^ {(reg62 ?
                  reg89 : reg45)})))
            begin
              for (forvar111 = (1'h0); (forvar111 < (1'h1)); forvar111 = (forvar111 + (1'h1)))
                begin
                  if ({(^~$signed((^(8'hae))))})
                    begin
                      reg112 <= $signed({(((8'hb3) <= (8'had)) ?
                              ((8'ha6) >> reg19) : (8'hb7))});
                      reg113 <= (({(reg70 && reg39)} >> (((8'hb1) ?
                          (8'h9d) : reg48) && $signed(reg88))) | (reg76[(1'h0):(1'h0)] != {(reg83 | reg40)}));
                      reg114 <= (~&$unsigned((+$unsigned(reg17))));
                      reg115 <= $unsigned((~|({reg56} ? reg39 : reg16)));
                    end
                  else
                    begin
                      reg112 <= $signed($signed($unsigned((~|reg71))));
                    end
                  for (forvar116 = (1'h0); (forvar116 < (1'h1)); forvar116 = (forvar116 + (1'h1)))
                    begin
                      reg117 <= reg98;
                      reg118 <= (reg23[(1'h0):(1'h0)] ?
                          {($unsigned(reg52) == reg35)} : $unsigned(((reg85 ?
                              reg99 : reg76) != (reg72 ? reg61 : reg73))));
                    end
                end
              for (forvar119 = (1'h0); (forvar119 < (2'h3)); forvar119 = (forvar119 + (1'h1)))
                begin
                  if ($unsigned((($unsigned(reg30) < (reg40 >> reg43)) ?
                      ((^~forvar110) * (reg104 == (8'hb8))) : $signed((!reg63)))))
                    begin
                      reg120 <= (reg44[(3'h5):(2'h3)] >= (|{(&reg48)}));
                      reg121 <= (reg40 >>> {reg19});
                    end
                  else
                    begin
                      reg120 <= $signed($unsigned(((~&(8'had)) * (reg42 ?
                          reg69 : reg102))));
                      reg121 <= (^$unsigned(($signed(reg94) ?
                          forvar110 : (!(8'hb5)))));
                      reg122 <= $unsigned($signed($signed(reg18[(3'h4):(2'h3)])));
                    end
                  if (((reg97 ^~ reg55) ? (!$signed(reg106)) : {{reg76}}))
                    begin
                      reg123 <= (($signed((reg26 << reg45)) ?
                          reg20[(4'hd):(2'h3)] : ((wire9 ?
                              reg94 : reg81) || $signed(reg109))) & reg84);
                      reg124 <= reg88[(1'h0):(1'h0)];
                      reg125 <= $signed($signed((((8'had) <= (8'hac)) ?
                          reg90[(4'ha):(3'h7)] : (reg113 ?
                              reg73 : forvar119))));
                    end
                  else
                    begin
                      reg123 <= (~|$unsigned(($unsigned((8'h9c)) ?
                          $signed(reg17) : reg46)));
                      reg124 <= $signed((+$signed(reg103)));
                      reg125 <= $signed((reg124[(1'h0):(1'h0)] ?
                          $unsigned($signed(wire8)) : ((reg81 == reg51) ?
                              {reg109} : reg31[(3'h4):(3'h4)])));
                      reg126 <= (~^reg29[(2'h3):(1'h0)]);
                    end
                end
            end
          else
            begin
              if ((&(^~(^$signed(reg68)))))
                begin
                  for (forvar111 = (1'h0); (forvar111 < (2'h3)); forvar111 = (forvar111 + (1'h1)))
                    begin
                      reg112 <= {$signed(reg61[(1'h1):(1'h0)])};
                      reg113 <= $unsigned((!reg54));
                      reg114 <= (!(|reg50));
                    end
                end
              else
                begin
                  for (forvar111 = (1'h0); (forvar111 < (1'h0)); forvar111 = (forvar111 + (1'h1)))
                    begin
                      reg112 <= (~^reg44[(2'h2):(1'h0)]);
                      reg113 <= (reg51[(4'h8):(3'h7)] ?
                          ((^(~^(8'hab))) || ($signed(reg94) >= $unsigned(reg125))) : ($unsigned($unsigned((8'hb8))) == reg99));
                      reg114 <= $signed(((reg73 <= $signed(reg19)) ?
                          $signed(reg66) : $unsigned(reg72)));
                      reg115 <= $signed(reg57[(1'h1):(1'h0)]);
                    end
                end
              for (forvar116 = (1'h0); (forvar116 < (1'h0)); forvar116 = (forvar116 + (1'h1)))
                begin
                  for (forvar117 = (1'h0); (forvar117 < (1'h1)); forvar117 = (forvar117 + (1'h1)))
                    begin
                      reg118 <= $unsigned($unsigned(((|reg29) * {reg54})));
                    end
                  for (forvar119 = (1'h0); (forvar119 < (2'h2)); forvar119 = (forvar119 + (1'h1)))
                    begin
                      reg120 <= (^(((^reg64) ? {reg102} : (reg28 * reg115)) ?
                          reg62[(1'h0):(1'h0)] : $signed($unsigned(reg27))));
                      reg121 <= (~&(($unsigned(reg52) ? reg59 : wire6) ?
                          wire10[(3'h6):(2'h2)] : $signed((~(8'hb0)))));
                    end
                  for (forvar122 = (1'h0); (forvar122 < (1'h1)); forvar122 = (forvar122 + (1'h1)))
                    begin
                      reg123 <= (reg72[(1'h0):(1'h0)] ?
                          $unsigned((^~$unsigned(reg99))) : (|$signed(((8'hb0) >= reg51))));
                      reg124 <= ((&(forvar111 ?
                          $signed(reg97) : (^reg28))) * (~|reg28[(1'h0):(1'h0)]));
                      reg125 <= $signed((!(!reg64[(2'h3):(2'h2)])));
                      reg126 <= $signed((8'ha3));
                    end
                end
            end
          for (forvar127 = (1'h0); (forvar127 < (2'h2)); forvar127 = (forvar127 + (1'h1)))
            begin
              if ((forvar116 ?
                  (^~reg50[(2'h3):(2'h3)]) : ({(-reg75)} ?
                      ((8'hb7) <<< reg51) : reg99)))
                begin
                  reg128 <= {(reg72 ~^ (reg83[(3'h4):(1'h0)] >>> (reg18 ?
                          reg68 : reg19)))};
                  if (((({(8'ha8)} ?
                              reg29[(3'h4):(2'h3)] : reg56[(4'h8):(3'h6)]) ?
                          $signed(reg57[(1'h1):(1'h0)]) : (&reg18)) ?
                      $signed(((wire6 != reg31) ?
                          forvar116 : (~|wire6))) : $signed(reg19)))
                    begin
                      reg129 <= (reg39[(3'h6):(3'h6)] << (($unsigned((8'ha4)) <= {reg112}) | reg100[(2'h2):(2'h2)]));
                      reg130 <= (reg103[(2'h3):(2'h2)] && $signed($unsigned(((8'h9f) >= reg103))));
                    end
                  else
                    begin
                      reg129 <= $unsigned(($signed($unsigned(reg28)) || (8'ha0)));
                      reg130 <= $signed((+({forvar111} ?
                          (reg123 ^ (8'hb8)) : ((8'hb4) ^ reg109))));
                    end
                  if ($signed(reg64))
                    begin
                      reg131 <= ($signed((reg130[(5'h10):(4'hc)] || $unsigned(forvar116))) ?
                          reg44 : reg114);
                      reg132 <= $unsigned($signed((|$signed((8'ha5)))));
                    end
                  else
                    begin
                      reg131 <= (({$unsigned(reg121)} ?
                          ((reg69 ? reg16 : reg85) ?
                              $unsigned(reg37) : reg98) : $signed((~^forvar111))) ~^ $signed($unsigned(wire6[(4'ha):(1'h1)])));
                      reg132 <= $signed(reg97[(4'h8):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar128 = (1'h0); (forvar128 < (1'h0)); forvar128 = (forvar128 + (1'h1)))
                    begin
                      reg129 <= (8'hb7);
                    end
                  for (forvar130 = (1'h0); (forvar130 < (2'h2)); forvar130 = (forvar130 + (1'h1)))
                    begin
                      reg131 <= reg18;
                      reg132 <= ((8'hb7) ~^ $unsigned(reg49[(2'h3):(2'h3)]));
                      reg133 <= (!(((8'hb8) + reg39) ?
                          {(forvar111 * reg90)} : reg53[(3'h7):(3'h5)]));
                      reg134 <= (-$signed((|(-(8'hba)))));
                    end
                end
            end
          for (forvar135 = (1'h0); (forvar135 < (2'h3)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 <= (^~reg17);
            end
          for (forvar137 = (1'h0); (forvar137 < (2'h2)); forvar137 = (forvar137 + (1'h1)))
            begin
              for (forvar138 = (1'h0); (forvar138 < (1'h1)); forvar138 = (forvar138 + (1'h1)))
                begin
                  if ($signed($unsigned(reg94[(2'h2):(1'h1)])))
                    begin
                      reg139 <= (^~(^(reg117[(3'h4):(2'h3)] >> reg31[(3'h6):(2'h3)])));
                      reg140 <= (~(-(8'h9e)));
                      reg141 <= ($unsigned(reg85) | $unsigned((reg90 ~^ (8'had))));
                      reg142 <= {reg128[(2'h3):(1'h1)]};
                    end
                  else
                    begin
                      reg139 <= $signed(($signed((reg118 ? reg114 : reg45)) ?
                          reg139[(1'h0):(1'h0)] : $unsigned($unsigned(reg35))));
                    end
                  reg143 <= {(+((^~reg17) ?
                          ((8'ha4) >>> (8'hb7)) : ((8'h9e) ? reg50 : reg99)))};
                  reg144 <= {$signed(reg141)};
                end
              for (forvar145 = (1'h0); (forvar145 < (2'h3)); forvar145 = (forvar145 + (1'h1)))
                begin
                  for (forvar146 = (1'h0); (forvar146 < (2'h2)); forvar146 = (forvar146 + (1'h1)))
                    begin
                      reg147 <= ($signed((~^{reg78})) ?
                          reg42[(1'h0):(1'h0)] : (~reg94[(2'h2):(1'h0)]));
                      reg148 <= (^(8'h9d));
                      reg149 <= reg81;
                    end
                  for (forvar150 = (1'h0); (forvar150 < (2'h3)); forvar150 = (forvar150 + (1'h1)))
                    begin
                      reg151 <= (~forvar130);
                      reg152 <= ((8'ha1) + ((((8'hba) ? reg69 : reg54) ?
                          reg100 : $unsigned(reg117)) > {$signed(reg124)}));
                    end
                end
              if ((($signed((forvar128 ?
                  reg101 : reg106)) == ($unsigned((8'hb7)) ?
                  reg143[(3'h4):(3'h4)] : $unsigned(wire8))) || forvar116))
                begin
                  for (forvar153 = (1'h0); (forvar153 < (2'h2)); forvar153 = (forvar153 + (1'h1)))
                    begin
                      reg154 <= reg22[(4'hb):(4'ha)];
                      reg155 <= ($unsigned(({reg82} ?
                          reg97 : (reg23 && reg24))) <= (~&((reg99 ?
                              wire9 : reg114) ?
                          $signed(forvar130) : $unsigned(reg94))));
                      reg156 <= {forvar137[(3'h4):(1'h1)]};
                    end
                  for (forvar157 = (1'h0); (forvar157 < (1'h0)); forvar157 = (forvar157 + (1'h1)))
                    begin
                      reg158 <= {$signed((!$signed(reg154)))};
                      reg159 <= ($unsigned(((8'ha4) && (reg121 <= reg133))) ?
                          $unsigned(wire6[(4'h9):(3'h5)]) : reg154[(3'h7):(1'h1)]);
                      reg160 <= reg142;
                    end
                end
              else
                begin
                  if ((|wire8))
                    begin
                      reg153 <= reg136;
                    end
                  else
                    begin
                      reg153 <= (($signed(reg133) ?
                          reg66[(1'h0):(1'h0)] : $unsigned($signed(reg68))) != (reg118[(3'h7):(1'h1)] ?
                          $unsigned($signed(reg63)) : reg156));
                      reg154 <= (~&($unsigned((reg43 ?
                          reg35 : (8'ha2))) & ((~^(8'hae)) ?
                          (reg101 ? reg151 : wire10) : reg32)));
                      reg155 <= (!($signed((~^reg100)) ?
                          $signed(wire6[(1'h1):(1'h1)]) : {$signed(reg99)}));
                      reg156 <= $signed(reg82);
                    end
                end
              for (forvar161 = (1'h0); (forvar161 < (2'h2)); forvar161 = (forvar161 + (1'h1)))
                begin
                  if (((^~{reg126[(3'h6):(3'h6)]}) << ((~^{reg26}) << reg156)))
                    begin
                      reg162 <= {$unsigned((reg48[(1'h0):(1'h0)] + (reg55 ?
                              reg22 : (8'had))))};
                      reg163 <= {(8'h9c)};
                      reg164 <= {((+{reg148}) ?
                              reg67 : ((^forvar117) < (8'hb1)))};
                      reg165 <= $signed((reg94[(1'h0):(1'h0)] ?
                          ($unsigned(reg20) ?
                              $signed(reg88) : $unsigned(forvar150)) : forvar117[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg162 <= ((~^reg147[(2'h2):(1'h0)]) ? reg69 : (8'hb9));
                      reg163 <= $unsigned(reg99);
                      reg164 <= (~^(((reg24 ? reg63 : reg41) - (reg42 ?
                              (8'ha1) : reg136)) ?
                          ($unsigned(forvar146) || (8'hb9)) : reg17[(3'h7):(2'h2)]));
                      reg165 <= $unsigned(((~&(reg125 && reg70)) ?
                          ((reg42 ?
                              reg136 : reg132) == (~|reg113)) : ((|reg158) << (8'hb9))));
                    end
                end
            end
        end
      if ($unsigned(($signed($unsigned(wire6)) ? reg156 : {reg65})))
        begin
          for (forvar166 = (1'h0); (forvar166 < (2'h2)); forvar166 = (forvar166 + (1'h1)))
            begin
              for (forvar167 = (1'h0); (forvar167 < (2'h2)); forvar167 = (forvar167 + (1'h1)))
                begin
                  if (forvar127[(4'ha):(4'ha)])
                    begin
                      reg168 <= (reg44 != {$signed(forvar166[(2'h2):(1'h1)])});
                    end
                  else
                    begin
                      reg168 <= $unsigned({(+(reg71 & (8'hb2)))});
                      reg169 <= $signed((^reg53));
                      reg170 <= ((forvar138[(3'h5):(1'h0)] + ((~&reg45) | (forvar161 + reg46))) << reg29);
                      reg171 <= {forvar166};
                    end
                  if ($signed({$signed((8'ha6))}))
                    begin
                      reg172 <= reg91[(3'h5):(2'h2)];
                      reg173 <= reg46;
                    end
                  else
                    begin
                      reg172 <= reg35[(4'h8):(1'h1)];
                    end
                  for (forvar174 = (1'h0); (forvar174 < (2'h2)); forvar174 = (forvar174 + (1'h1)))
                    begin
                      reg175 <= $signed(forvar116[(3'h6):(2'h2)]);
                      reg176 <= (8'ha2);
                    end
                  if (reg121)
                    begin
                      reg177 <= $signed($signed(((reg132 ? reg27 : wire11) ?
                          {reg37} : {(8'hb6)})));
                    end
                  else
                    begin
                      reg177 <= (reg41 ? reg35 : $signed(reg50));
                      reg178 <= reg17[(4'hc):(3'h6)];
                    end
                end
              reg179 <= $unsigned(({(reg48 > reg94)} <<< {reg78[(1'h1):(1'h1)]}));
            end
          reg180 <= (!{reg20[(1'h1):(1'h0)]});
        end
      else
        begin
          for (forvar166 = (1'h0); (forvar166 < (1'h0)); forvar166 = (forvar166 + (1'h1)))
            begin
              reg167 <= $unsigned($unsigned((reg101[(1'h1):(1'h0)] <= (^reg162))));
            end
          for (forvar168 = (1'h0); (forvar168 < (1'h1)); forvar168 = (forvar168 + (1'h1)))
            begin
              reg169 <= $unsigned((~&forvar127[(4'hc):(4'hc)]));
              for (forvar170 = (1'h0); (forvar170 < (2'h2)); forvar170 = (forvar170 + (1'h1)))
                begin
                  for (forvar171 = (1'h0); (forvar171 < (2'h2)); forvar171 = (forvar171 + (1'h1)))
                    begin
                      reg172 <= reg20;
                      reg173 <= reg39[(2'h2):(1'h0)];
                    end
                  reg174 <= forvar153[(3'h4):(2'h2)];
                end
              reg175 <= reg159;
            end
          for (forvar176 = (1'h0); (forvar176 < (1'h0)); forvar176 = (forvar176 + (1'h1)))
            begin
              for (forvar177 = (1'h0); (forvar177 < (1'h1)); forvar177 = (forvar177 + (1'h1)))
                begin
                  for (forvar178 = (1'h0); (forvar178 < (2'h3)); forvar178 = (forvar178 + (1'h1)))
                    begin
                      reg179 <= (+forvar145[(3'h6):(2'h2)]);
                      reg180 <= (!(-(~|reg89[(4'he):(3'h6)])));
                      reg181 <= $unsigned(($unsigned((reg59 ? reg134 : wire8)) ?
                          ((reg100 ?
                              reg128 : forvar171) ~^ reg141[(1'h0):(1'h0)]) : $unsigned(wire11)));
                    end
                  reg182 <= (8'hb2);
                end
              for (forvar183 = (1'h0); (forvar183 < (2'h2)); forvar183 = (forvar183 + (1'h1)))
                begin
                  if ((|(-$signed(reg50))))
                    begin
                      reg184 <= forvar146;
                      reg185 <= ((|{((8'ha9) ? forvar127 : reg100)}) ?
                          (forvar117 ?
                              reg184 : (+((8'ha2) ?
                                  reg98 : forvar137))) : (reg122[(1'h1):(1'h1)] ?
                              $unsigned(reg96) : (|(^(8'ha3)))));
                      reg186 <= (reg180 << {reg153[(4'he):(4'h9)]});
                    end
                  else
                    begin
                      reg184 <= (^~($signed((~|reg48)) ~^ reg125));
                      reg185 <= $signed((((reg133 + forvar110) ?
                              reg174 : $signed(reg152)) ?
                          forvar167[(2'h2):(1'h0)] : $signed(reg152)));
                    end
                  for (forvar187 = (1'h0); (forvar187 < (1'h0)); forvar187 = (forvar187 + (1'h1)))
                    begin
                      reg188 <= $signed($unsigned({(reg170 > reg168)}));
                      reg189 <= $unsigned(reg88);
                      reg190 <= {reg28[(2'h2):(2'h2)]};
                      reg191 <= reg17[(1'h1):(1'h1)];
                    end
                  for (forvar192 = (1'h0); (forvar192 < (2'h2)); forvar192 = (forvar192 + (1'h1)))
                    begin
                      reg193 <= $signed($signed(reg147));
                    end
                end
              for (forvar194 = (1'h0); (forvar194 < (1'h1)); forvar194 = (forvar194 + (1'h1)))
                begin
                  if ($unsigned((&{$signed(reg32)})))
                    begin
                      reg195 <= (^~$signed((^~(+reg134))));
                      reg196 <= reg190[(3'h4):(2'h3)];
                      reg197 <= {forvar192};
                    end
                  else
                    begin
                      reg195 <= $signed({reg66[(1'h0):(1'h0)]});
                    end
                  reg198 <= ($unsigned($unsigned((reg149 ?
                      reg41 : reg153))) - $unsigned(((^reg140) - (!forvar117))));
                end
            end
          for (forvar199 = (1'h0); (forvar199 < (2'h3)); forvar199 = (forvar199 + (1'h1)))
            begin
              reg200 <= $signed(({$signed(reg154)} > ((~&(8'ha3)) ^ (reg48 ?
                  reg88 : reg112))));
            end
        end
      for (forvar201 = (1'h0); (forvar201 < (2'h2)); forvar201 = (forvar201 + (1'h1)))
        begin
          for (forvar202 = (1'h0); (forvar202 < (2'h2)); forvar202 = (forvar202 + (1'h1)))
            begin
              if ($unsigned($unsigned(reg130)))
                begin
                  for (forvar203 = (1'h0); (forvar203 < (1'h0)); forvar203 = (forvar203 + (1'h1)))
                    begin
                      reg204 <= ($signed((-reg113)) ? reg189 : wire7);
                      reg205 <= $signed((reg29[(3'h4):(1'h0)] ^ $unsigned((reg40 ?
                          forvar128 : reg136))));
                      reg206 <= $unsigned(reg147);
                      reg207 <= ($signed($signed($unsigned(reg29))) - reg51[(1'h0):(1'h0)]);
                    end
                  reg208 <= $unsigned((&(reg50[(4'hb):(4'h9)] ?
                      (reg123 & (8'ha1)) : reg37)));
                  reg209 <= ($signed(((!reg160) ?
                          $signed(forvar183) : ((8'hb1) ? forvar153 : reg29))) ?
                      {({wire10} << {forvar150})} : $unsigned(((reg197 * reg37) ?
                          forvar199[(4'h8):(2'h3)] : (~forvar117))));
                  if (((({reg53} ?
                      (reg22 ?
                          forvar178 : reg50) : forvar157) >> (forvar176[(2'h3):(2'h2)] > (reg32 ?
                      reg63 : reg139))) >= forvar202))
                    begin
                      reg210 <= ((((reg164 * (8'ha2)) ?
                              forvar119[(2'h2):(2'h2)] : (~reg172)) ?
                          forvar119 : ($unsigned(reg120) ?
                              $unsigned(reg101) : (reg98 & reg55))) >>> (+reg44[(2'h2):(1'h1)]));
                      reg211 <= (!reg19);
                      reg212 <= ({($unsigned(forvar157) ?
                                  reg83[(2'h3):(1'h1)] : $unsigned(reg207))} ?
                          $signed(reg70) : (~^($signed(reg125) ?
                              reg186[(2'h2):(2'h2)] : (reg144 ?
                                  reg197 : reg177))));
                      reg213 <= reg49;
                    end
                  else
                    begin
                      reg210 <= reg30;
                    end
                end
              else
                begin
                  reg203 <= {reg139[(3'h7):(1'h1)]};
                  if ((-reg73))
                    begin
                      reg204 <= $unsigned(((reg45[(4'ha):(2'h3)] ?
                          (reg85 ? forvar145 : forvar110) : (reg124 ?
                              reg205 : reg109)) != (reg148[(1'h0):(1'h0)] ?
                          (^~(8'h9e)) : (reg27 ? reg174 : reg83))));
                      reg205 <= $signed(reg142);
                      reg206 <= $unsigned(reg66);
                    end
                  else
                    begin
                      reg204 <= ((reg204[(3'h5):(3'h4)] ?
                          reg131[(4'h9):(4'h9)] : reg52[(3'h6):(3'h4)]) >> {(reg155[(2'h2):(2'h2)] != (!reg148))});
                      reg205 <= ((&reg44[(3'h5):(1'h0)]) || ((((8'hb9) ^~ reg76) ?
                          (reg156 ?
                              reg200 : (8'hab)) : $signed(reg176)) >> $signed(reg90[(3'h5):(3'h5)])));
                      reg206 <= ((|reg107) ?
                          reg69[(3'h4):(2'h3)] : (reg204 <<< ($signed(reg168) || {reg83})));
                      reg207 <= (!$unsigned({forvar176[(4'hb):(4'hb)]}));
                    end
                  for (forvar208 = (1'h0); (forvar208 < (1'h0)); forvar208 = (forvar208 + (1'h1)))
                    begin
                      reg209 <= reg130[(3'h4):(1'h1)];
                      reg210 <= $unsigned(wire10[(3'h5):(2'h2)]);
                      reg211 <= (((^{forvar135}) ?
                              (reg112[(1'h1):(1'h1)] ?
                                  (~reg52) : (8'haf)) : $signed(reg56)) ?
                          forvar146 : ((((8'ha2) ? (8'ha0) : reg117) ?
                              $unsigned(reg167) : (forvar128 ?
                                  forvar171 : reg107)) != (reg209 ?
                              reg69 : $unsigned((8'ha0)))));
                    end
                end
              if ($signed(reg149[(1'h1):(1'h0)]))
                begin
                  reg214 <= ((~(reg63[(3'h6):(1'h0)] <<< (forvar171 || forvar192))) ^ $unsigned((|$signed(reg109))));
                  for (forvar215 = (1'h0); (forvar215 < (2'h2)); forvar215 = (forvar215 + (1'h1)))
                    begin
                      reg216 <= reg198;
                      reg217 <= $unsigned(($signed(reg147) ?
                          reg62[(2'h3):(2'h2)] : reg151));
                      reg218 <= (((wire7 ?
                                  $unsigned(reg23) : reg27[(3'h7):(3'h4)]) ?
                              $signed((~^(8'hab))) : $unsigned(reg19)) ?
                          forvar192 : reg104[(2'h3):(2'h3)]);
                    end
                  for (forvar219 = (1'h0); (forvar219 < (2'h2)); forvar219 = (forvar219 + (1'h1)))
                    begin
                      reg220 <= ((forvar215 >> reg155[(2'h3):(2'h2)]) > {reg144[(3'h4):(2'h3)]});
                    end
                  for (forvar221 = (1'h0); (forvar221 < (2'h2)); forvar221 = (forvar221 + (1'h1)))
                    begin
                      reg222 <= (^~$unsigned({reg115}));
                      reg223 <= reg214;
                      reg224 <= reg152;
                      reg225 <= {reg99[(2'h2):(2'h2)]};
                    end
                end
              else
                begin
                  for (forvar214 = (1'h0); (forvar214 < (1'h1)); forvar214 = (forvar214 + (1'h1)))
                    begin
                      reg215 <= (($unsigned({(8'hb6)}) ?
                          {reg61} : forvar127[(2'h2):(1'h0)]) >>> reg214[(4'h8):(1'h0)]);
                      reg216 <= $signed($signed(reg101[(4'h9):(3'h4)]));
                      reg217 <= reg147;
                      reg218 <= ((~&(~^(reg26 ? reg109 : (8'hb0)))) ?
                          ((forvar170[(4'h9):(4'h8)] ?
                              reg23 : $signed(reg117)) * $signed(reg81[(3'h4):(1'h1)])) : $signed((reg169 >= $signed(reg41))));
                    end
                  reg219 <= (reg125 ^ $unsigned({(~|reg72)}));
                  for (forvar220 = (1'h0); (forvar220 < (1'h0)); forvar220 = (forvar220 + (1'h1)))
                    begin
                      reg221 <= (forvar220[(3'h5):(1'h1)] ?
                          $unsigned({$signed(forvar176)}) : $signed(reg170[(3'h4):(1'h1)]));
                      reg222 <= (((8'h9d) > $signed(reg144)) <<< (((8'h9c) ?
                          (reg39 && reg56) : (|forvar221)) & ((~reg216) ?
                          {forvar192} : (reg124 <= reg44))));
                      reg223 <= ((~|$unsigned((reg225 ? reg113 : reg156))) ?
                          (reg51[(1'h1):(1'h0)] ?
                              forvar145 : ({(8'hba)} ~^ $unsigned((8'haa)))) : reg17);
                      reg224 <= reg73;
                    end
                  if ({$signed(reg200[(4'h8):(1'h1)])})
                    begin
                      reg225 <= $signed({(reg115[(1'h1):(1'h0)] ?
                              reg31[(3'h6):(2'h2)] : (reg65 <<< forvar199))});
                      reg226 <= $signed(reg98);
                      reg227 <= reg142;
                    end
                  else
                    begin
                      reg225 <= reg131[(4'he):(4'hc)];
                      reg226 <= ((reg112[(4'h8):(4'h8)] ?
                              {$signed((8'ha7))} : $unsigned({(8'ha8)})) ?
                          (reg216 < (|$signed(reg70))) : reg117[(3'h4):(2'h2)]);
                      reg227 <= $unsigned(((^reg153[(3'h6):(3'h6)]) > (reg154[(1'h0):(1'h0)] == reg51)));
                    end
                end
            end
          for (forvar228 = (1'h0); (forvar228 < (1'h1)); forvar228 = (forvar228 + (1'h1)))
            begin
              for (forvar229 = (1'h0); (forvar229 < (2'h3)); forvar229 = (forvar229 + (1'h1)))
                begin
                  reg230 <= reg82;
                  reg231 <= ($unsigned($unsigned((reg226 ?
                          reg214 : forvar146))) ?
                      (wire11[(2'h3):(2'h2)] || (reg132[(4'h9):(1'h0)] ?
                          {forvar117} : (forvar194 ^~ reg17))) : reg225);
                end
            end
        end
      for (forvar232 = (1'h0); (forvar232 < (2'h3)); forvar232 = (forvar232 + (1'h1)))
        begin
          if (reg144)
            begin
              for (forvar233 = (1'h0); (forvar233 < (2'h3)); forvar233 = (forvar233 + (1'h1)))
                begin
                  for (forvar234 = (1'h0); (forvar234 < (2'h2)); forvar234 = (forvar234 + (1'h1)))
                    begin
                      reg235 <= ($signed({$signed(forvar153)}) > (~|$signed($unsigned(reg68))));
                    end
                  if ((!(-(!$signed(reg104)))))
                    begin
                      reg236 <= {reg124};
                    end
                  else
                    begin
                      reg236 <= $unsigned(($unsigned((reg20 == (8'ha6))) ?
                          (reg158[(4'ha):(2'h2)] | reg55[(2'h3):(2'h2)]) : ($signed(reg77) + ((8'ha3) >>> reg142))));
                      reg237 <= {$unsigned(forvar138)};
                      reg238 <= forvar170[(4'he):(3'h7)];
                      reg239 <= $unsigned(wire10);
                    end
                  for (forvar240 = (1'h0); (forvar240 < (1'h0)); forvar240 = (forvar240 + (1'h1)))
                    begin
                      reg241 <= forvar228[(3'h5):(3'h4)];
                    end
                end
            end
          else
            begin
              if ((~$signed(({forvar116} ? {forvar240} : (!forvar187)))))
                begin
                  if ((!$unsigned((forvar146 ? {(8'ha2)} : reg168))))
                    begin
                      reg233 <= reg68[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg233 <= ({reg94[(2'h2):(1'h1)]} ?
                          $unsigned(((~|forvar146) ?
                              $signed(forvar240) : reg101)) : (8'h9c));
                      reg234 <= $signed((|reg43));
                      reg235 <= ((~|((reg33 ? forvar215 : reg200) ?
                              {reg43} : reg209[(2'h2):(1'h1)])) ?
                          (~&$signed(reg88[(4'ha):(4'h9)])) : (&(-(~|reg164))));
                      reg236 <= (-(reg129 ? reg172 : reg211));
                    end
                  if (((reg126[(1'h1):(1'h1)] * ((forvar202 ?
                      forvar202 : reg143) <<< reg18)) + (($signed(reg175) < ((8'h9c) ?
                          reg17 : reg70)) ?
                      forvar177 : (reg57[(1'h0):(1'h0)] ?
                          (^forvar219) : (reg241 + reg88)))))
                    begin
                      reg237 <= $signed((~^(reg106 ?
                          reg24[(2'h2):(1'h0)] : reg162)));
                      reg238 <= (~^($unsigned({forvar194}) ?
                          reg176[(3'h5):(3'h5)] : $signed((-reg227))));
                      reg239 <= $signed($signed($unsigned(((8'hb4) ?
                          reg76 : reg91))));
                    end
                  else
                    begin
                      reg237 <= ($signed(reg204) >>> $unsigned($unsigned((^~reg151))));
                      reg238 <= reg43;
                      reg239 <= $signed((^{(reg100 ? reg88 : reg169)}));
                      reg240 <= (reg65 == (reg162 ?
                          (reg78[(1'h1):(1'h1)] + $signed(reg89)) : ({wire10} & $unsigned((8'ha9)))));
                    end
                end
              else
                begin
                  for (forvar233 = (1'h0); (forvar233 < (2'h2)); forvar233 = (forvar233 + (1'h1)))
                    begin
                      reg234 <= $unsigned(((8'hab) << reg49));
                      reg235 <= $signed({forvar170[(3'h6):(1'h0)]});
                      reg236 <= reg76;
                    end
                  for (forvar237 = (1'h0); (forvar237 < (1'h1)); forvar237 = (forvar237 + (1'h1)))
                    begin
                      reg238 <= (!($unsigned(reg57[(4'h9):(4'h8)]) ~^ ((forvar232 >> (8'hb7)) << {reg77})));
                      reg239 <= $unsigned((+forvar178));
                    end
                end
              for (forvar241 = (1'h0); (forvar241 < (2'h2)); forvar241 = (forvar241 + (1'h1)))
                begin
                  reg242 <= (reg71 ?
                      $unsigned((8'ha6)) : ($unsigned((reg131 ?
                              reg217 : forvar130)) ?
                          ($signed(reg175) ?
                              (reg52 ^ reg102) : $unsigned(reg49)) : (8'hb6)));
                  for (forvar243 = (1'h0); (forvar243 < (1'h0)); forvar243 = (forvar243 + (1'h1)))
                    begin
                      reg244 <= $unsigned({{forvar232[(4'ha):(4'ha)]}});
                      reg245 <= ((~(forvar214 != $unsigned(reg122))) || (reg234[(4'h9):(4'h9)] ?
                          reg219[(1'h0):(1'h0)] : ({reg131} ~^ $signed(reg139))));
                      reg246 <= $unsigned(({$unsigned(reg23)} <= reg167[(4'ha):(3'h5)]));
                    end
                end
            end
          if ($signed($unsigned(forvar150[(1'h0):(1'h0)])))
            begin
              for (forvar247 = (1'h0); (forvar247 < (2'h3)); forvar247 = (forvar247 + (1'h1)))
                begin
                  if ($unsigned(reg162[(2'h3):(1'h1)]))
                    begin
                      reg248 <= reg94[(2'h2):(1'h1)];
                      reg249 <= {$unsigned(((&reg41) ?
                              $unsigned(reg65) : reg158))};
                      reg250 <= (($unsigned($unsigned(reg124)) == reg33[(2'h2):(1'h0)]) | $unsigned($signed(reg189)));
                      reg251 <= (+reg233);
                    end
                  else
                    begin
                      reg248 <= (-$unsigned($unsigned($signed((8'ha6)))));
                      reg249 <= (+$signed($unsigned((8'hb4))));
                      reg250 <= (-(reg117 ?
                          $unsigned(reg234) : (~|wire7[(1'h0):(1'h0)])));
                    end
                  for (forvar252 = (1'h0); (forvar252 < (2'h3)); forvar252 = (forvar252 + (1'h1)))
                    begin
                      reg253 <= (^((!(reg209 >>> reg197)) ?
                          reg152[(1'h0):(1'h0)] : $unsigned($signed(reg73))));
                    end
                end
              for (forvar254 = (1'h0); (forvar254 < (2'h2)); forvar254 = (forvar254 + (1'h1)))
                begin
                  if ((forvar201[(1'h0):(1'h0)] && ((~^(reg123 ?
                      reg94 : reg58)) << {(+reg213)})))
                    begin
                      reg255 <= {(-$unsigned($unsigned(reg129)))};
                      reg256 <= $unsigned($signed(reg51));
                      reg257 <= ($unsigned((reg218[(1'h0):(1'h0)] ?
                              (~&(8'haf)) : $signed(forvar221))) ?
                          (&(|((8'hb2) >= reg244))) : (reg65[(1'h0):(1'h0)] >> ((reg133 <= reg27) ?
                              (forvar153 ? (8'hb4) : reg197) : (reg100 ?
                                  reg94 : reg224))));
                    end
                  else
                    begin
                      reg255 <= forvar241[(2'h2):(1'h1)];
                      reg256 <= $unsigned((reg207 ?
                          reg172[(4'hb):(1'h0)] : $signed($signed((8'ha5)))));
                      reg257 <= $signed(($signed(forvar176) ?
                          reg102 : $signed($unsigned(reg32))));
                      reg258 <= $signed(($unsigned($signed(forvar192)) == (reg57[(4'h8):(1'h1)] ?
                          {reg227} : (reg193 && reg241))));
                    end
                end
              if ($signed(((|$signed(reg142)) ?
                  $unsigned(((8'hb2) ?
                      reg32 : reg236)) : (reg164 * reg203[(1'h0):(1'h0)]))))
                begin
                  if ((8'ha8))
                    begin
                      reg259 <= $unsigned(({$unsigned(reg170)} && (8'hb9)));
                      reg260 <= $unsigned(reg259);
                      reg261 <= reg140[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg259 <= $unsigned((reg251 > $signed((forvar117 >>> reg217))));
                      reg260 <= forvar138;
                      reg261 <= (|$unsigned(reg131));
                    end
                end
              else
                begin
                  if (reg213)
                    begin
                      reg259 <= reg100[(4'hb):(1'h1)];
                      reg260 <= $unsigned({reg100[(4'hc):(2'h2)]});
                      reg261 <= reg249;
                      reg262 <= {($unsigned((forvar201 <<< (8'hb3))) ~^ $unsigned($signed(reg71)))};
                    end
                  else
                    begin
                      reg259 <= $signed((8'h9c));
                    end
                  if (reg198[(4'hb):(4'ha)])
                    begin
                      reg263 <= wire6;
                    end
                  else
                    begin
                      reg263 <= $signed({reg143[(4'h9):(3'h6)]});
                      reg264 <= forvar199;
                    end
                end
            end
          else
            begin
              reg247 <= ((reg219[(2'h3):(2'h2)] || reg26) & reg133[(4'h8):(3'h7)]);
              for (forvar248 = (1'h0); (forvar248 < (2'h2)); forvar248 = (forvar248 + (1'h1)))
                begin
                  for (forvar249 = (1'h0); (forvar249 < (2'h3)); forvar249 = (forvar249 + (1'h1)))
                    begin
                      reg250 <= {(reg241 > ({(8'hac)} ?
                              $signed(forvar243) : (~(8'hb5))))};
                      reg251 <= reg180[(1'h0):(1'h0)];
                      reg252 <= ((^(|(^reg170))) ?
                          ($signed(reg117) != $signed(reg190[(1'h1):(1'h0)])) : reg261);
                    end
                  reg253 <= {(~(~^$unsigned(reg158)))};
                  reg254 <= (((~&(reg141 ?
                      forvar153 : reg248)) & $unsigned((^(8'hae)))) * (|({reg164} ?
                      (forvar130 ? reg168 : reg185) : $signed(reg99))));
                end
            end
        end
    end
  assign wire265 = $signed((-(reg42[(1'h0):(1'h0)] ?
                       $signed(wire10) : (reg122 != reg136))));
  assign wire266 = reg44[(3'h4):(2'h2)];
  assign wire267 = reg153;
  assign wire268 = ($signed(reg122) ?
                       reg209[(2'h3):(2'h2)] : ({(reg76 ? reg249 : reg95)} ?
                           $unsigned($unsigned(reg230)) : ((8'haf) + reg162[(4'h9):(3'h6)])));
  always
    @(posedge clk) begin
      if ($signed(($unsigned($signed(reg240)) ?
          reg149 : ({reg129} < {reg225}))))
        begin
          if ({($signed(reg124) <= reg67)})
            begin
              for (forvar269 = (1'h0); (forvar269 < (2'h3)); forvar269 = (forvar269 + (1'h1)))
                begin
                  for (forvar270 = (1'h0); (forvar270 < (2'h3)); forvar270 = (forvar270 + (1'h1)))
                    begin
                      reg271 <= {(reg224 - reg33[(3'h5):(3'h5)])};
                    end
                  reg272 <= reg176;
                  for (forvar273 = (1'h0); (forvar273 < (2'h3)); forvar273 = (forvar273 + (1'h1)))
                    begin
                      reg274 <= {reg186};
                      reg275 <= $signed(({$signed(reg109)} + $unsigned(reg224[(4'he):(4'hc)])));
                      reg276 <= $signed((~&(wire7 ^ (reg195 ?
                          reg261 : (8'hb8)))));
                      reg277 <= reg96;
                    end
                end
            end
          else
            begin
              for (forvar269 = (1'h0); (forvar269 < (2'h3)); forvar269 = (forvar269 + (1'h1)))
                begin
                  reg270 <= {{($signed(reg184) ? reg237 : (~^(8'hb9)))}};
                  for (forvar271 = (1'h0); (forvar271 < (1'h1)); forvar271 = (forvar271 + (1'h1)))
                    begin
                      reg272 <= reg54;
                      reg273 <= reg85;
                      reg274 <= wire10[(3'h7):(3'h7)];
                      reg275 <= $signed((&reg141[(3'h5):(2'h2)]));
                    end
                  if ((wire9[(1'h0):(1'h0)] ?
                      (reg275 ?
                          {$unsigned((8'hb3))} : $signed($unsigned((8'had)))) : {(reg30 > (reg214 ?
                              reg48 : reg227))}))
                    begin
                      reg276 <= {$unsigned($signed((^reg64)))};
                      reg277 <= reg106[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg276 <= reg121[(3'h7):(1'h1)];
                      reg277 <= ((+$unsigned(reg128[(4'hc):(4'hc)])) + $signed($unsigned(reg88)));
                      reg278 <= reg41;
                    end
                end
            end
          for (forvar279 = (1'h0); (forvar279 < (1'h1)); forvar279 = (forvar279 + (1'h1)))
            begin
              for (forvar280 = (1'h0); (forvar280 < (2'h3)); forvar280 = (forvar280 + (1'h1)))
                begin
                  if ($unsigned($signed($signed((reg219 ? (8'hae) : reg241)))))
                    begin
                      reg281 <= ($unsigned($signed((reg121 ?
                          reg238 : reg52))) >= reg100[(1'h0):(1'h0)]);
                      reg282 <= (~|$unsigned($signed(((8'haf) <= reg48))));
                      reg283 <= reg171[(3'h7):(3'h4)];
                    end
                  else
                    begin
                      reg281 <= $unsigned($signed(reg143[(3'h4):(1'h1)]));
                    end
                  reg284 <= {($signed($unsigned(reg88)) >> $unsigned($signed(reg88)))};
                  for (forvar285 = (1'h0); (forvar285 < (1'h0)); forvar285 = (forvar285 + (1'h1)))
                    begin
                      reg286 <= reg103;
                      reg287 <= ((8'hb3) >> reg174);
                      reg288 <= $signed(reg198[(4'h9):(2'h2)]);
                    end
                end
              if (reg195)
                begin
                  reg289 <= (^~{$signed((wire6 >>> reg249))});
                  if (($unsigned(reg33[(4'h9):(2'h2)]) ?
                      ($unsigned(reg176[(2'h3):(1'h1)]) - reg133) : (+(reg109 * reg52))))
                    begin
                      reg290 <= reg179[(4'h8):(2'h2)];
                      reg291 <= reg149;
                      reg292 <= ($signed({(reg122 ?
                              reg261 : reg261)}) >= reg283);
                      reg293 <= (~|{reg59});
                    end
                  else
                    begin
                      reg290 <= reg275[(2'h3):(2'h3)];
                      reg291 <= (reg70[(5'h10):(4'hf)] && ({reg70} < reg83[(2'h3):(2'h3)]));
                      reg292 <= reg284[(2'h2):(1'h0)];
                      reg293 <= {reg35};
                    end
                end
              else
                begin
                  if (reg20)
                    begin
                      reg289 <= {reg237};
                      reg290 <= ({$signed(reg101)} * (~^{(!(8'ha2))}));
                    end
                  else
                    begin
                      reg289 <= ((($signed(reg59) ? {wire10} : $signed(reg30)) ?
                              $unsigned(reg144[(1'h0):(1'h0)]) : $signed((reg149 * reg236))) ?
                          {(reg273 == (reg24 ? reg23 : reg51))} : (reg125 ?
                              {$signed(wire267)} : $unsigned(((8'hba) ?
                                  reg70 : reg225))));
                      reg290 <= reg182[(4'ha):(3'h7)];
                    end
                  reg291 <= ((~|($unsigned(reg57) & $unsigned(reg155))) ?
                      ({$signed(reg179)} + {reg128}) : (+{$signed(wire9)}));
                  for (forvar292 = (1'h0); (forvar292 < (2'h3)); forvar292 = (forvar292 + (1'h1)))
                    begin
                      reg293 <= $signed(($signed($unsigned(reg78)) & reg203));
                      reg294 <= $unsigned(reg23[(3'h7):(1'h1)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar269 = (1'h0); (forvar269 < (2'h2)); forvar269 = (forvar269 + (1'h1)))
            begin
              reg270 <= reg275[(1'h0):(1'h0)];
              for (forvar271 = (1'h0); (forvar271 < (2'h2)); forvar271 = (forvar271 + (1'h1)))
                begin
                  if (reg154[(3'h7):(3'h4)])
                    begin
                      reg272 <= reg159[(1'h0):(1'h0)];
                      reg273 <= reg37;
                      reg274 <= (($unsigned($unsigned(reg89)) ?
                          $signed(reg262) : ($signed(reg68) ?
                              reg19[(3'h7):(3'h7)] : ((8'ha5) <= forvar269))) == reg274[(1'h1):(1'h1)]);
                      reg275 <= (-(&((-reg113) & reg164)));
                    end
                  else
                    begin
                      reg272 <= (8'ha5);
                      reg273 <= (((-reg216) ^ (8'hb0)) ?
                          ({$unsigned((8'ha8))} || (!(^~(8'haa)))) : (((reg274 == reg181) ?
                                  $unsigned(reg48) : reg222) ?
                              $unsigned(reg19) : (~|(^forvar280))));
                      reg274 <= $signed(reg177[(3'h4):(2'h3)]);
                      reg275 <= ((~|(^~$signed(reg142))) ?
                          ($unsigned(reg286) ?
                              {(reg260 ?
                                      reg272 : reg55)} : $unsigned(reg236)) : $signed(($unsigned(reg253) ?
                              (wire267 ?
                                  (8'hb0) : reg270) : wire266[(2'h3):(2'h3)])));
                    end
                  if (((~^($signed(forvar270) ?
                      $signed((8'ha4)) : (reg242 ?
                          reg275 : reg84))) << ((~^{reg102}) ?
                      $unsigned({reg235}) : (~|(~|(8'hb1))))))
                    begin
                      reg276 <= $signed((wire7 << $signed($signed(reg49))));
                    end
                  else
                    begin
                      reg276 <= ((+((reg179 ?
                              (8'ha2) : forvar279) << forvar273)) ?
                          ((reg224[(3'h7):(2'h3)] | reg281) ?
                              wire267[(3'h7):(2'h3)] : $signed($unsigned(reg209))) : {{{reg250}}});
                    end
                  for (forvar277 = (1'h0); (forvar277 < (2'h3)); forvar277 = (forvar277 + (1'h1)))
                    begin
                      reg278 <= reg101[(4'ha):(1'h0)];
                    end
                  for (forvar279 = (1'h0); (forvar279 < (1'h0)); forvar279 = (forvar279 + (1'h1)))
                    begin
                      reg280 <= (8'h9d);
                      reg281 <= (&reg294);
                      reg282 <= $signed($signed($unsigned($unsigned(wire265))));
                    end
                end
              reg283 <= $signed($signed($signed((reg154 ? reg56 : reg104))));
              if (($signed(reg289[(4'he):(3'h7)]) ?
                  (reg57[(2'h3):(1'h0)] ?
                      wire11 : $signed((wire10 ?
                          reg230 : reg41))) : {((^~reg240) < (~&reg82))}))
                begin
                  reg284 <= (((reg217[(4'h9):(3'h6)] ?
                              reg198[(1'h1):(1'h1)] : (reg242 ?
                                  reg162 : (8'ha0))) ?
                          reg220[(3'h4):(1'h0)] : (&$unsigned(wire8))) ?
                      reg147 : {((reg57 - forvar285) ~^ (~^wire6))});
                  reg285 <= wire7;
                  for (forvar286 = (1'h0); (forvar286 < (2'h3)); forvar286 = (forvar286 + (1'h1)))
                    begin
                      reg287 <= reg282;
                      reg288 <= $unsigned(reg84[(4'h9):(3'h7)]);
                      reg289 <= reg246;
                    end
                  for (forvar290 = (1'h0); (forvar290 < (1'h1)); forvar290 = (forvar290 + (1'h1)))
                    begin
                      reg291 <= (({{reg275}} ?
                          ((~(8'hab)) & (&reg237)) : (~&$unsigned((8'ha7)))) && $signed(($signed(reg179) ?
                          ((8'ha6) ^~ reg130) : $unsigned(reg66))));
                      reg292 <= $signed(wire9[(3'h5):(1'h1)]);
                      reg293 <= $unsigned((reg52 ?
                          $unsigned((!wire9)) : reg154));
                      reg294 <= ((($unsigned(reg58) ?
                                  forvar290[(1'h1):(1'h1)] : (~&reg41)) ?
                              $unsigned(reg124[(2'h2):(2'h2)]) : reg84) ?
                          $unsigned({(reg274 - (8'hb7))}) : $unsigned($signed(reg198)));
                    end
                end
              else
                begin
                  if (reg278[(3'h5):(1'h1)])
                    begin
                      reg284 <= ({reg75[(4'ha):(3'h6)]} == $unsigned((&(-reg32))));
                    end
                  else
                    begin
                      reg284 <= (~^$signed(({reg238} > $unsigned(reg151))));
                      reg285 <= $signed(((reg96[(3'h4):(1'h1)] >= (reg224 + reg57)) ?
                          (~$unsigned((8'hb0))) : reg122[(3'h6):(2'h3)]));
                    end
                end
            end
          for (forvar295 = (1'h0); (forvar295 < (1'h0)); forvar295 = (forvar295 + (1'h1)))
            begin
              for (forvar296 = (1'h0); (forvar296 < (2'h3)); forvar296 = (forvar296 + (1'h1)))
                begin
                  if ((reg242[(2'h2):(1'h0)] <<< reg211[(2'h3):(1'h1)]))
                    begin
                      reg297 <= reg278[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg297 <= wire7[(3'h4):(2'h3)];
                      reg298 <= $unsigned(((^reg49[(2'h2):(1'h0)]) || $signed(reg56)));
                    end
                end
            end
          if (reg289[(5'h10):(1'h0)])
            begin
              for (forvar299 = (1'h0); (forvar299 < (1'h1)); forvar299 = (forvar299 + (1'h1)))
                begin
                  for (forvar300 = (1'h0); (forvar300 < (2'h2)); forvar300 = (forvar300 + (1'h1)))
                    begin
                      reg301 <= ((~&(+$unsigned(reg272))) & reg168[(3'h7):(3'h4)]);
                      reg302 <= reg52[(3'h7):(1'h1)];
                      reg303 <= (+$unsigned(((reg207 && (8'h9c)) << (~|reg85))));
                    end
                  for (forvar304 = (1'h0); (forvar304 < (2'h3)); forvar304 = (forvar304 + (1'h1)))
                    begin
                      reg305 <= reg97[(3'h5):(1'h1)];
                    end
                end
              if ({(-{reg16[(2'h2):(1'h1)]})})
                begin
                  if ({$unsigned($unsigned(reg203[(4'hb):(2'h3)]))})
                    begin
                      reg306 <= reg245;
                      reg307 <= reg52[(4'hc):(3'h4)];
                      reg308 <= $unsigned(((8'h9c) < $unsigned(reg258)));
                    end
                  else
                    begin
                      reg306 <= $unsigned(forvar286);
                      reg307 <= ($signed(($signed(reg83) > reg148)) ?
                          reg59 : (!$unsigned({(8'h9c)})));
                    end
                  if ((|$signed({$unsigned(reg247)})))
                    begin
                      reg309 <= (^($signed((reg273 ? reg275 : reg50)) ?
                          reg176 : (reg91 ?
                              $unsigned(reg66) : $unsigned((8'hb1)))));
                      reg310 <= (8'hac);
                    end
                  else
                    begin
                      reg309 <= ((($signed(forvar277) | {reg310}) ?
                          (^(reg96 > reg281)) : (reg19[(3'h4):(3'h4)] ~^ $signed(reg120))) * $signed(reg255[(2'h3):(1'h1)]));
                    end
                  for (forvar311 = (1'h0); (forvar311 < (1'h1)); forvar311 = (forvar311 + (1'h1)))
                    begin
                      reg312 <= $unsigned(((reg262[(3'h6):(1'h0)] || forvar271) == $unsigned((reg42 ^ reg254))));
                      reg313 <= $signed(((8'hb1) + $unsigned(((8'h9f) << reg292))));
                    end
                  for (forvar314 = (1'h0); (forvar314 < (2'h2)); forvar314 = (forvar314 + (1'h1)))
                    begin
                      reg315 <= $signed(((reg214[(4'hc):(3'h4)] + $unsigned(reg234)) ?
                          (((8'ha6) != reg98) ?
                              $unsigned(reg244) : $unsigned(forvar299)) : {(~&reg257)}));
                      reg316 <= {{$signed($unsigned(reg50))}};
                    end
                end
              else
                begin
                  reg306 <= reg78;
                end
            end
          else
            begin
              if ((reg312[(1'h0):(1'h0)] || reg73[(1'h1):(1'h1)]))
                begin
                  for (forvar299 = (1'h0); (forvar299 < (2'h3)); forvar299 = (forvar299 + (1'h1)))
                    begin
                      reg300 <= (reg143[(3'h7):(3'h5)] && reg289);
                      reg301 <= reg274[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  if (reg124[(2'h2):(1'h1)])
                    begin
                      reg299 <= (reg99[(3'h5):(3'h5)] ?
                          $signed(reg46[(3'h6):(3'h6)]) : ((&(reg170 > reg272)) >> {(&reg312)}));
                      reg300 <= reg216;
                    end
                  else
                    begin
                      reg299 <= $signed(reg271);
                      reg300 <= $signed(({reg185[(2'h2):(1'h1)]} - (8'h9d)));
                      reg301 <= ((reg179[(4'h8):(2'h2)] <<< reg65) == $unsigned((reg278[(3'h4):(1'h0)] ~^ (8'hae))));
                    end
                  if ($signed(((!(~^reg142)) <<< ((reg276 ? (8'hb9) : (8'hab)) ?
                      (~|forvar314) : reg205))))
                    begin
                      reg302 <= $unsigned({($unsigned(reg57) ?
                              reg148[(1'h0):(1'h0)] : reg113[(2'h2):(1'h1)])});
                    end
                  else
                    begin
                      reg302 <= reg147[(1'h0):(1'h0)];
                      reg303 <= (^(($signed(reg305) ^~ (reg84 >= reg262)) ?
                          {$signed(reg124)} : $unsigned((~^reg106))));
                    end
                end
              for (forvar304 = (1'h0); (forvar304 < (1'h0)); forvar304 = (forvar304 + (1'h1)))
                begin
                  if (reg285[(4'h9):(3'h4)])
                    begin
                      reg305 <= ($unsigned($signed((reg143 ?
                              (8'hb7) : reg57))) ?
                          ((^((8'hb7) << reg165)) ?
                              (^(reg62 >>> reg259)) : $signed((forvar300 ^~ reg278))) : $unsigned(forvar273[(2'h3):(1'h1)]));
                      reg306 <= (~reg101);
                      reg307 <= reg84;
                      reg308 <= ($signed((8'hb4)) > reg255);
                    end
                  else
                    begin
                      reg305 <= $unsigned($unsigned(reg315));
                      reg306 <= (reg106[(3'h6):(2'h2)] ?
                          ($signed((^~reg106)) ?
                              $unsigned((reg43 ~^ reg257)) : {$signed((8'hac))}) : (-$unsigned((~&reg69))));
                    end
                  reg309 <= (&($signed($unsigned(forvar311)) ?
                      $unsigned((!reg68)) : ((~&reg204) ?
                          (wire265 ? (8'haf) : reg124) : reg159)));
                  for (forvar310 = (1'h0); (forvar310 < (1'h1)); forvar310 = (forvar310 + (1'h1)))
                    begin
                      reg311 <= reg30[(2'h2):(1'h1)];
                      reg312 <= ($unsigned($signed(reg303)) * (~(~{reg252})));
                      reg313 <= $signed(($unsigned($signed(reg216)) ?
                          ({reg154} >= (reg55 != reg48)) : ((reg156 < wire8) ?
                              reg259 : $signed(reg242))));
                    end
                end
              reg314 <= ((&reg255) ?
                  $unsigned({$signed(reg136)}) : (reg117[(2'h2):(1'h1)] + reg182[(3'h7):(2'h2)]));
            end
        end
      if ($unsigned(reg82[(1'h1):(1'h0)]))
        begin
          reg317 <= reg104[(1'h0):(1'h0)];
          for (forvar318 = (1'h0); (forvar318 < (2'h2)); forvar318 = (forvar318 + (1'h1)))
            begin
              reg319 <= $unsigned(($signed($signed(reg309)) + reg222[(3'h4):(2'h3)]));
              for (forvar320 = (1'h0); (forvar320 < (1'h0)); forvar320 = (forvar320 + (1'h1)))
                begin
                  for (forvar321 = (1'h0); (forvar321 < (2'h3)); forvar321 = (forvar321 + (1'h1)))
                    begin
                      reg322 <= {$signed($signed(reg128[(4'hd):(2'h3)]))};
                      reg323 <= $signed(reg64[(2'h2):(1'h1)]);
                      reg324 <= (+((^~wire9) ?
                          (((8'hae) && (8'hb4)) ?
                              reg43 : (|reg272)) : (reg210[(1'h1):(1'h0)] ?
                              reg239 : (^~(8'ha5)))));
                      reg325 <= $unsigned((~(((8'hb3) ?
                          wire266 : (8'ha6)) + reg294[(3'h4):(2'h2)])));
                    end
                  if ((reg122 ?
                      ($unsigned((^~reg49)) ^ ((reg95 ? reg178 : reg284) ?
                          $unsigned(reg239) : (reg95 ?
                              (8'had) : reg287))) : ($signed($unsigned(reg216)) != (8'hb9))))
                    begin
                      reg326 <= ($signed((reg180[(2'h3):(1'h1)] ?
                              (-reg126) : (reg315 ? reg144 : wire6))) ?
                          {reg136} : $unsigned(reg237[(2'h3):(2'h2)]));
                      reg327 <= reg174[(4'hd):(1'h1)];
                    end
                  else
                    begin
                      reg326 <= (^(~^($unsigned((8'hb7)) << (reg319 ?
                          reg200 : reg106))));
                      reg327 <= reg144;
                      reg328 <= (!(^~$unsigned(((8'ha6) ^~ wire11))));
                    end
                  for (forvar329 = (1'h0); (forvar329 < (1'h0)); forvar329 = (forvar329 + (1'h1)))
                    begin
                      reg330 <= reg287;
                      reg331 <= (~|($signed((-reg195)) && ((reg104 ?
                              reg224 : reg298) ?
                          forvar290 : (reg253 & forvar292))));
                      reg332 <= (-(|($unsigned(reg213) ?
                          (reg159 || reg156) : $unsigned(reg249))));
                    end
                  for (forvar333 = (1'h0); (forvar333 < (1'h0)); forvar333 = (forvar333 + (1'h1)))
                    begin
                      reg334 <= (8'hb0);
                    end
                end
            end
          for (forvar335 = (1'h0); (forvar335 < (2'h2)); forvar335 = (forvar335 + (1'h1)))
            begin
              for (forvar336 = (1'h0); (forvar336 < (2'h2)); forvar336 = (forvar336 + (1'h1)))
                begin
                  if ($signed(reg258))
                    begin
                      reg337 <= $unsigned((((reg124 ?
                              reg219 : reg75) ^~ ((8'hb1) ? reg327 : (8'hb8))) ?
                          $unsigned(reg251[(4'h9):(3'h7)]) : $signed({reg84})));
                      reg338 <= (reg173[(4'hd):(2'h2)] ?
                          (!(reg176 <<< (~&reg57))) : reg327[(3'h5):(3'h4)]);
                      reg339 <= reg82;
                      reg340 <= $signed(reg160[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg337 <= {(^~(reg222[(1'h0):(1'h0)] ?
                              {(8'ha0)} : (~&reg340)))};
                    end
                  for (forvar341 = (1'h0); (forvar341 < (1'h1)); forvar341 = (forvar341 + (1'h1)))
                    begin
                      reg342 <= $signed($signed(reg316));
                    end
                end
            end
          if ((+forvar270))
            begin
              for (forvar343 = (1'h0); (forvar343 < (2'h3)); forvar343 = (forvar343 + (1'h1)))
                begin
                  if (({$unsigned(reg178)} << (~|reg58)))
                    begin
                      reg344 <= reg283;
                    end
                  else
                    begin
                      reg344 <= (8'haf);
                      reg345 <= {{((~&reg54) ?
                                  (reg35 ?
                                      reg241 : reg154) : $unsigned(reg158))}};
                      reg346 <= $unsigned(($unsigned($signed(reg27)) << $unsigned((wire267 ?
                          reg49 : reg325))));
                      reg347 <= ($signed($signed(reg292[(3'h6):(3'h4)])) & {reg323[(3'h6):(1'h1)]});
                    end
                  for (forvar348 = (1'h0); (forvar348 < (2'h2)); forvar348 = (forvar348 + (1'h1)))
                    begin
                      reg349 <= (reg143[(2'h3):(1'h0)] ?
                          reg195[(3'h4):(1'h1)] : (~(!(reg337 ?
                              reg156 : reg344))));
                      reg350 <= (reg235[(1'h0):(1'h0)] - reg231);
                    end
                  if ($unsigned(reg136[(3'h5):(3'h4)]))
                    begin
                      reg351 <= (^~($unsigned({reg177}) ?
                          $unsigned(forvar348[(1'h1):(1'h1)]) : ((^reg247) ?
                              (reg163 < reg283) : (~|reg227))));
                      reg352 <= ({($unsigned(forvar333) ?
                              ((8'ha1) << reg126) : (8'ha4))} >= (8'had));
                      reg353 <= {forvar292};
                      reg354 <= $signed($signed(((reg19 ? forvar296 : reg317) ?
                          reg103[(4'h9):(3'h6)] : $signed(wire267))));
                    end
                  else
                    begin
                      reg351 <= (($signed($signed(reg62)) ?
                          (+$unsigned(reg185)) : ($unsigned(reg16) >= reg130)) || $unsigned(reg61));
                      reg352 <= $signed($unsigned($unsigned((reg255 ?
                          reg68 : reg325))));
                      reg353 <= (reg225 >>> (|{(~|reg102)}));
                    end
                  reg355 <= (((forvar336[(1'h1):(1'h0)] ?
                          $signed(reg154) : (~^reg207)) && ((^~reg18) ?
                          (forvar318 ? reg237 : reg319) : (8'hb6))) ?
                      reg97[(1'h0):(1'h0)] : reg40);
                end
            end
          else
            begin
              for (forvar343 = (1'h0); (forvar343 < (2'h2)); forvar343 = (forvar343 + (1'h1)))
                begin
                  if ({$unsigned(reg33)})
                    begin
                      reg344 <= $signed($unsigned(((reg76 ?
                          reg342 : (8'hb5)) + (reg50 ? (8'ha4) : reg148))));
                      reg345 <= ((reg236 + ($signed(reg89) ?
                          $signed(reg288) : (reg94 ?
                              forvar341 : reg315))) ^~ (((-reg49) > (~&reg263)) >> ($signed(reg148) ?
                          wire7 : $signed((8'hb5)))));
                    end
                  else
                    begin
                      reg344 <= {(reg78 >> $signed({reg128}))};
                      reg345 <= {$signed(reg325[(3'h7):(1'h0)])};
                      reg346 <= reg283;
                      reg347 <= reg51[(4'he):(1'h0)];
                    end
                end
              for (forvar348 = (1'h0); (forvar348 < (1'h1)); forvar348 = (forvar348 + (1'h1)))
                begin
                  reg349 <= $signed(((+((8'hb1) ?
                      reg101 : reg307)) + (reg114 ^ reg78)));
                end
              for (forvar350 = (1'h0); (forvar350 < (1'h1)); forvar350 = (forvar350 + (1'h1)))
                begin
                  if (((($unsigned((8'hb2)) | (reg261 ?
                          reg139 : reg317)) <<< $signed($unsigned(reg59))) ?
                      reg351[(1'h0):(1'h0)] : $signed(($unsigned(reg190) * ((8'ha9) ?
                          (8'haf) : reg235)))))
                    begin
                      reg351 <= {(-(-(reg290 > reg281)))};
                      reg352 <= (($unsigned(reg204) ?
                              $unsigned($unsigned(reg235)) : ((reg160 ?
                                      reg54 : forvar343) ?
                                  reg112 : reg186)) ?
                          ($signed((reg68 ?
                              reg303 : reg209)) < reg81) : $unsigned((^(reg212 ?
                              reg136 : reg195))));
                      reg353 <= (({(reg50 ? reg165 : reg22)} ?
                          ($signed(reg214) ?
                              $signed(reg160) : reg104[(4'he):(4'hd)]) : $unsigned((reg331 != reg184))) ~^ $signed({reg217[(3'h4):(1'h0)]}));
                    end
                  else
                    begin
                      reg351 <= {((|reg272[(3'h6):(1'h1)]) * $signed(reg307[(2'h3):(2'h3)]))};
                      reg352 <= (((^~(forvar270 ?
                          reg273 : reg115)) >= reg41[(4'hd):(3'h7)]) * $unsigned(reg99[(3'h5):(1'h0)]));
                      reg353 <= (8'hba);
                    end
                end
              if ((|(~|reg96[(3'h4):(3'h4)])))
                begin
                  for (forvar354 = (1'h0); (forvar354 < (1'h0)); forvar354 = (forvar354 + (1'h1)))
                    begin
                      reg355 <= reg217[(4'hd):(4'hd)];
                    end
                  for (forvar356 = (1'h0); (forvar356 < (1'h0)); forvar356 = (forvar356 + (1'h1)))
                    begin
                      reg357 <= {(~&(~^(reg165 < reg104)))};
                      reg358 <= (({(reg128 ?
                              reg136 : reg191)} <= reg163[(4'hc):(1'h0)]) >>> (~|$unsigned((|wire265))));
                      reg359 <= (((~|(forvar273 ? reg208 : (8'hb2))) ?
                          $unsigned($unsigned(reg131)) : reg64) || reg236);
                      reg360 <= (8'h9d);
                    end
                end
              else
                begin
                  for (forvar354 = (1'h0); (forvar354 < (2'h3)); forvar354 = (forvar354 + (1'h1)))
                    begin
                      reg355 <= (~|reg141[(1'h0):(1'h0)]);
                    end
                end
            end
        end
      else
        begin
          if (($unsigned(reg294[(4'hd):(3'h4)]) * ((reg215 ?
                  ((8'hac) ? reg78 : forvar341) : (reg316 && reg189)) ?
              ((&reg153) || (reg225 ?
                  (8'hb5) : (8'ha5))) : $signed($signed(reg62)))))
            begin
              for (forvar317 = (1'h0); (forvar317 < (2'h3)); forvar317 = (forvar317 + (1'h1)))
                begin
                  for (forvar318 = (1'h0); (forvar318 < (2'h3)); forvar318 = (forvar318 + (1'h1)))
                    begin
                      reg319 <= (reg133[(3'h5):(2'h3)] ?
                          {reg264[(1'h0):(1'h0)]} : (((+forvar335) ?
                                  {reg169} : (reg220 != reg186)) ?
                              {(reg85 & forvar321)} : ((8'hae) >= (^~reg89))));
                      reg320 <= {(~reg83)};
                      reg321 <= $signed((($unsigned(reg322) ?
                              $signed(reg163) : (reg300 ? reg96 : reg67)) ?
                          (|reg350[(2'h2):(2'h2)]) : $unsigned(reg196[(4'ha):(3'h4)])));
                      reg322 <= $signed($unsigned((8'h9e)));
                    end
                end
            end
          else
            begin
              if ($unsigned((reg33 ?
                  $unsigned($unsigned(reg274)) : $signed((reg311 ?
                      reg303 : (8'ha0))))))
                begin
                  for (forvar317 = (1'h0); (forvar317 < (1'h0)); forvar317 = (forvar317 + (1'h1)))
                    begin
                      reg318 <= (reg94 == (8'ha1));
                      reg319 <= (^~reg94);
                      reg320 <= (({$unsigned(reg29)} ?
                              $unsigned((reg52 ?
                                  reg215 : reg253)) : $signed((|reg36))) ?
                          (~((8'ha2) ?
                              (reg323 & (8'hb2)) : (forvar280 ?
                                  reg195 : forvar336))) : reg123);
                      reg321 <= ({$signed((~|reg37))} ?
                          reg278 : {$signed(forvar350)});
                    end
                  if ((^~{reg40[(1'h0):(1'h0)]}))
                    begin
                      reg322 <= reg301[(4'hb):(4'ha)];
                      reg323 <= forvar295[(4'h9):(3'h7)];
                    end
                  else
                    begin
                      reg322 <= reg95;
                      reg323 <= {$signed(($unsigned(wire265) * (8'ha1)))};
                      reg324 <= (^(({reg107} <<< {reg78}) >> reg89));
                    end
                end
              else
                begin
                  for (forvar317 = (1'h0); (forvar317 < (2'h2)); forvar317 = (forvar317 + (1'h1)))
                    begin
                      reg318 <= $signed(reg22);
                      reg319 <= $unsigned(reg308[(2'h3):(1'h0)]);
                      reg320 <= forvar270[(2'h2):(2'h2)];
                    end
                  reg321 <= (reg290[(2'h2):(2'h2)] >>> $unsigned(reg128));
                  if ($signed($unsigned($unsigned((reg128 ?
                      forvar350 : forvar286)))))
                    begin
                      reg322 <= (8'hb8);
                      reg323 <= reg315[(4'ha):(4'h8)];
                      reg324 <= ((^~(+{reg19})) ?
                          (&reg238[(4'h8):(1'h0)]) : (~&(~|(~^reg50))));
                      reg325 <= ($unsigned($signed(reg244[(2'h3):(1'h1)])) ?
                          {((reg315 ?
                                  reg325 : reg152) - {(8'hab)})} : $unsigned((reg262[(3'h6):(1'h0)] ?
                              forvar317 : $signed((8'haa)))));
                    end
                  else
                    begin
                      reg322 <= (&$signed(reg51));
                      reg323 <= reg184[(2'h3):(2'h3)];
                      reg324 <= ({$signed(reg148)} ?
                          ($signed($signed((8'hb2))) && reg344) : $unsigned(((-reg35) & $unsigned((8'hac)))));
                      reg325 <= ((&reg233[(1'h1):(1'h0)]) ?
                          reg326[(1'h1):(1'h1)] : $unsigned((((8'ha1) ~^ (8'ha2)) ?
                              {reg241} : (8'hba))));
                    end
                end
              if ((((forvar270[(2'h3):(1'h1)] ?
                          reg239[(2'h2):(1'h1)] : forvar350[(1'h1):(1'h0)]) ?
                      (8'hb0) : reg30[(1'h1):(1'h1)]) ?
                  $unsigned(($signed(reg217) ?
                      reg134[(1'h0):(1'h0)] : ((8'hb3) - reg272))) : ($signed((^~forvar286)) >>> $unsigned($unsigned(reg196)))))
                begin
                  for (forvar326 = (1'h0); (forvar326 < (1'h1)); forvar326 = (forvar326 + (1'h1)))
                    begin
                      reg327 <= (~&((^forvar295) ?
                          forvar321 : $signed(reg257)));
                      reg328 <= $unsigned($signed(((reg311 ?
                              forvar280 : reg89) ?
                          $unsigned(reg99) : $signed(reg285))));
                      reg329 <= (+((|reg36[(3'h5):(1'h0)]) ~^ {$unsigned(reg241)}));
                      reg330 <= (^~reg99);
                    end
                  reg331 <= ((^reg221) ?
                      $signed(((~&reg181) >= (reg94 ^ reg40))) : $signed((^~$signed(reg36))));
                  if ((((reg23[(1'h0):(1'h0)] & {reg318}) ?
                      reg290 : $signed(reg283)) != {reg224[(4'hc):(3'h4)]}))
                    begin
                      reg332 <= reg121;
                      reg333 <= reg288[(3'h6):(3'h6)];
                      reg334 <= reg325[(4'h9):(3'h4)];
                      reg335 <= (8'haa);
                    end
                  else
                    begin
                      reg332 <= (((~|reg153[(4'hb):(4'hb)]) ?
                          ($signed(reg114) ?
                              $unsigned(reg178) : $unsigned(reg24)) : (~|$unsigned(reg235))) ^~ {(!{reg84})});
                    end
                  if ((~&($signed($unsigned(reg294)) <= (!reg216[(3'h6):(2'h2)]))))
                    begin
                      reg336 <= $unsigned(($unsigned({reg250}) ?
                          $signed(forvar348[(2'h2):(1'h0)]) : (|reg227[(2'h3):(2'h3)])));
                      reg337 <= {$unsigned(reg284[(2'h2):(2'h2)])};
                      reg338 <= (+reg312[(1'h0):(1'h0)]);
                      reg339 <= $unsigned(reg90[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg336 <= (8'haf);
                      reg337 <= reg181[(3'h7):(2'h3)];
                      reg338 <= ($signed($signed($unsigned(reg24))) ?
                          $unsigned($signed(reg55[(3'h5):(2'h3)])) : reg155[(2'h3):(1'h0)]);
                    end
                end
              else
                begin
                  if (reg301[(3'h6):(1'h0)])
                    begin
                      reg326 <= $signed(forvar333[(1'h0):(1'h0)]);
                      reg327 <= {(~|$signed((forvar304 ? reg288 : reg206)))};
                      reg328 <= {(~|reg339[(4'h9):(2'h3)])};
                    end
                  else
                    begin
                      reg326 <= $signed($signed(((&reg20) >> (reg328 ?
                          (8'hb2) : (8'hae)))));
                      reg327 <= $unsigned(reg124);
                      reg328 <= {(!(8'ha8))};
                    end
                end
            end
          for (forvar340 = (1'h0); (forvar340 < (2'h2)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 <= (!$signed($signed(reg236[(4'hb):(3'h6)])));
              reg342 <= (((reg354 < $unsigned(reg178)) ?
                      reg325[(4'ha):(4'h9)] : (reg197 < reg89)) ?
                  $signed($signed($signed(forvar336))) : forvar269[(3'h4):(1'h0)]);
              reg343 <= $signed(forvar295[(4'h8):(3'h5)]);
              for (forvar344 = (1'h0); (forvar344 < (1'h0)); forvar344 = (forvar344 + (1'h1)))
                begin
                  reg345 <= ((!((reg337 ? (8'ha8) : (8'ha7)) ?
                          forvar329[(2'h2):(2'h2)] : (~^reg51))) ?
                      {(reg200[(4'h9):(1'h0)] + $unsigned(reg118))} : reg186);
                  for (forvar346 = (1'h0); (forvar346 < (2'h2)); forvar346 = (forvar346 + (1'h1)))
                    begin
                      reg347 <= reg52;
                      reg348 <= $unsigned(((~^(reg151 ?
                          reg130 : reg36)) ^~ (reg256[(4'h9):(1'h0)] & ((8'hba) & reg327))));
                      reg349 <= $unsigned(reg334);
                      reg350 <= reg276;
                    end
                  reg351 <= $signed($unsigned($signed((reg227 || reg303))));
                end
            end
        end
      for (forvar361 = (1'h0); (forvar361 < (1'h0)); forvar361 = (forvar361 + (1'h1)))
        begin
          reg362 <= reg282[(3'h4):(2'h2)];
          reg363 <= $unsigned(($signed((reg335 ?
              forvar344 : reg245)) << reg164));
          if (forvar320[(4'h9):(4'h8)])
            begin
              if (reg200[(2'h2):(1'h0)])
                begin
                  for (forvar364 = (1'h0); (forvar364 < (2'h3)); forvar364 = (forvar364 + (1'h1)))
                    begin
                      reg365 <= $unsigned(((!(reg332 ? reg351 : reg352)) ?
                          reg283[(2'h2):(1'h0)] : ((~|forvar273) == (reg292 >>> (8'h9d)))));
                    end
                  for (forvar366 = (1'h0); (forvar366 < (1'h1)); forvar366 = (forvar366 + (1'h1)))
                    begin
                      reg367 <= reg365;
                      reg368 <= $unsigned((8'h9e));
                      reg369 <= (reg245[(3'h4):(2'h2)] * $signed($unsigned((reg324 ?
                          wire266 : reg102))));
                    end
                  for (forvar370 = (1'h0); (forvar370 < (2'h3)); forvar370 = (forvar370 + (1'h1)))
                    begin
                      reg371 <= {(8'hb6)};
                      reg372 <= ((($signed(reg355) ?
                                  (&forvar304) : (reg174 ? reg89 : reg342)) ?
                              (~|$unsigned(reg176)) : $unsigned($unsigned(reg231))) ?
                          ($unsigned((|(8'hac))) ?
                              $unsigned($unsigned(reg58)) : (reg262[(1'h1):(1'h0)] <<< {reg84})) : (reg113[(4'he):(4'he)] ?
                              $unsigned({(8'h9d)}) : $signed($signed(reg58))));
                      reg373 <= (8'ha6);
                    end
                end
              else
                begin
                  for (forvar364 = (1'h0); (forvar364 < (1'h1)); forvar364 = (forvar364 + (1'h1)))
                    begin
                      reg365 <= (8'hb4);
                      reg366 <= (reg165 == $signed($unsigned((!reg26))));
                      reg367 <= (reg48[(2'h2):(2'h2)] & $signed($unsigned({reg362})));
                    end
                  if (($signed((|(forvar314 > reg219))) + $unsigned({((8'haf) ?
                          reg237 : reg350)})))
                    begin
                      reg368 <= (reg206[(4'hf):(3'h5)] ?
                          $signed((|reg200[(2'h3):(2'h3)])) : $signed((!(reg22 ^ reg350))));
                      reg369 <= $unsigned(reg32);
                      reg370 <= ((+(reg317 < (~|reg239))) ~^ reg107);
                    end
                  else
                    begin
                      reg368 <= $unsigned({(reg298 ?
                              reg73 : reg289[(5'h10):(1'h1)])});
                      reg369 <= {$signed($unsigned((&reg276)))};
                      reg370 <= {$unsigned({(~|reg209)})};
                    end
                  if ((^((!$unsigned((8'hb7))) ?
                      $signed($signed((8'had))) : reg178)))
                    begin
                      reg371 <= reg152;
                      reg372 <= ((~&reg322) - $signed($signed($unsigned(reg181))));
                      reg373 <= (8'ha7);
                    end
                  else
                    begin
                      reg371 <= $signed((&(~|((8'hae) > forvar277))));
                    end
                end
              reg374 <= ((8'h9e) ?
                  ($signed($unsigned(reg198)) ?
                      ((reg354 << (8'ha0)) & (8'hb8)) : {reg220[(2'h2):(1'h0)]}) : reg222[(3'h7):(2'h3)]);
              for (forvar375 = (1'h0); (forvar375 < (1'h0)); forvar375 = (forvar375 + (1'h1)))
                begin
                  for (forvar376 = (1'h0); (forvar376 < (2'h2)); forvar376 = (forvar376 + (1'h1)))
                    begin
                      reg377 <= $signed((+wire268[(1'h1):(1'h0)]));
                    end
                end
              for (forvar378 = (1'h0); (forvar378 < (1'h1)); forvar378 = (forvar378 + (1'h1)))
                begin
                  if ($unsigned(reg24))
                    begin
                      reg379 <= (~|forvar340);
                      reg380 <= reg139;
                      reg381 <= (reg54 ? reg262[(4'hc):(4'ha)] : (8'hb8));
                      reg382 <= $unsigned($signed((reg290[(1'h0):(1'h0)] ?
                          (+reg315) : ((8'hb0) ? (8'ha8) : reg41))));
                    end
                  else
                    begin
                      reg379 <= ($signed($signed(reg185[(3'h4):(2'h3)])) + (|(-(reg134 ?
                          reg96 : reg345))));
                      reg380 <= reg149;
                    end
                end
            end
          else
            begin
              for (forvar364 = (1'h0); (forvar364 < (1'h1)); forvar364 = (forvar364 + (1'h1)))
                begin
                  for (forvar365 = (1'h0); (forvar365 < (1'h1)); forvar365 = (forvar365 + (1'h1)))
                    begin
                      reg366 <= $unsigned($signed((reg39[(3'h4):(1'h0)] ^~ (&reg341))));
                      reg367 <= (reg341[(2'h3):(2'h2)] || (forvar336[(2'h2):(1'h1)] ?
                          $unsigned({reg223}) : $unsigned((reg100 ?
                              reg24 : reg190))));
                      reg368 <= (-((8'hb4) ^ $unsigned($unsigned((8'hb3)))));
                      reg369 <= reg262[(4'h9):(1'h1)];
                    end
                  if ($unsigned((^~$signed(((8'hae) ? (8'h9e) : (8'hb4))))))
                    begin
                      reg370 <= $signed((((!reg377) <= $unsigned(reg42)) < reg147[(1'h1):(1'h1)]));
                      reg371 <= $unsigned((~reg178[(4'h8):(3'h7)]));
                    end
                  else
                    begin
                      reg370 <= reg65[(1'h1):(1'h1)];
                      reg371 <= reg316[(2'h3):(1'h0)];
                      reg372 <= ((~&{(~&reg294)}) <<< reg158[(4'ha):(1'h0)]);
                      reg373 <= $signed(($signed({reg330}) <= reg85[(3'h6):(1'h0)]));
                    end
                end
              reg374 <= $signed(reg248[(1'h0):(1'h0)]);
              for (forvar375 = (1'h0); (forvar375 < (1'h1)); forvar375 = (forvar375 + (1'h1)))
                begin
                  for (forvar376 = (1'h0); (forvar376 < (2'h3)); forvar376 = (forvar376 + (1'h1)))
                    begin
                      reg377 <= reg78[(1'h0):(1'h0)];
                      reg378 <= reg293[(4'hb):(3'h6)];
                    end
                end
              if (reg143[(1'h1):(1'h0)])
                begin
                  for (forvar379 = (1'h0); (forvar379 < (2'h3)); forvar379 = (forvar379 + (1'h1)))
                    begin
                      reg380 <= $unsigned(reg300[(1'h0):(1'h0)]);
                      reg381 <= (~^(((-reg102) ?
                              (reg35 ?
                                  forvar336 : forvar318) : $signed(forvar270)) ?
                          reg95[(3'h4):(1'h0)] : $signed(reg141)));
                      reg382 <= (reg275[(2'h2):(1'h1)] ? reg71 : (^~(8'hae)));
                      reg383 <= (&(~^{(reg233 ? (8'hb0) : forvar279)}));
                    end
                end
              else
                begin
                  if (((8'h9c) ?
                      reg342[(3'h4):(2'h3)] : $unsigned((-$unsigned((8'hab))))))
                    begin
                      reg379 <= ($signed(reg206) >= $signed(reg154[(2'h2):(2'h2)]));
                      reg380 <= (+reg124);
                      reg381 <= ((-reg57) <= (&$signed((reg120 ~^ reg219))));
                    end
                  else
                    begin
                      reg379 <= (8'hab);
                      reg380 <= $unsigned((&{$unsigned(reg65)}));
                      reg381 <= {$unsigned(forvar321)};
                    end
                end
            end
          reg384 <= $signed(((!{forvar370}) + $unsigned(((8'h9e) & forvar270))));
        end
    end
  module385 #() modinst536 (wire535, clk, reg260, reg68, reg324, reg329);
  always
    @(posedge clk) begin
      reg537 <= (((reg235[(1'h1):(1'h1)] << (reg216 - reg73)) ?
          ($unsigned(reg261) ?
              {(8'haa)} : {reg22}) : $signed(reg180[(2'h2):(2'h2)])) * $unsigned(reg141));
      reg538 <= {reg19[(3'h4):(2'h3)]};
      if ({reg274[(3'h4):(1'h0)]})
        begin
          for (forvar539 = (1'h0); (forvar539 < (2'h3)); forvar539 = (forvar539 + (1'h1)))
            begin
              for (forvar540 = (1'h0); (forvar540 < (2'h3)); forvar540 = (forvar540 + (1'h1)))
                begin
                  reg541 <= $unsigned((((reg122 && reg347) == (reg286 >>> (8'ha6))) ?
                      $signed((reg216 < reg367)) : $signed(reg253)));
                  for (forvar542 = (1'h0); (forvar542 < (1'h1)); forvar542 = (forvar542 + (1'h1)))
                    begin
                      reg543 <= (!$unsigned((8'hb5)));
                      reg544 <= $signed(reg354);
                      reg545 <= {((reg16[(3'h4):(1'h1)] != (reg106 ?
                              reg84 : (8'hb0))) >= reg32[(2'h2):(2'h2)])};
                    end
                  if ((|$unsigned({(reg147 * reg22)})))
                    begin
                      reg546 <= ((!$unsigned((reg181 ? (8'hb7) : reg293))) ?
                          ((+(&(8'hb4))) ?
                              $unsigned((&reg311)) : reg178) : $signed({(-reg330)}));
                      reg547 <= $unsigned((reg276 ?
                          (&{reg258}) : $unsigned($unsigned(reg373))));
                      reg548 <= reg130;
                      reg549 <= ((reg32 | {$unsigned(reg294)}) ?
                          reg90[(3'h4):(2'h3)] : (|((reg193 ?
                                  reg132 : (8'hb8)) ?
                              $signed(reg245) : (8'ha5))));
                    end
                  else
                    begin
                      reg546 <= (reg547[(2'h2):(2'h2)] << (^~$unsigned((reg294 ?
                          reg371 : reg340))));
                    end
                end
            end
          for (forvar550 = (1'h0); (forvar550 < (1'h0)); forvar550 = (forvar550 + (1'h1)))
            begin
              for (forvar551 = (1'h0); (forvar551 < (2'h2)); forvar551 = (forvar551 + (1'h1)))
                begin
                  reg552 <= ((^~{reg48}) ?
                      (~reg67[(1'h1):(1'h0)]) : reg195[(2'h3):(2'h2)]);
                  if ((reg345[(1'h1):(1'h0)] ~^ $signed(reg164)))
                    begin
                      reg553 <= ($unsigned(reg27[(3'h5):(2'h3)]) != (reg323[(3'h4):(1'h1)] + reg293[(4'ha):(3'h6)]));
                      reg554 <= (^(!reg84[(3'h5):(3'h4)]));
                    end
                  else
                    begin
                      reg553 <= ((($unsigned(reg225) << (8'ha9)) ?
                              reg360 : $unsigned(reg19[(3'h5):(1'h1)])) ?
                          (reg182 - (+$signed(reg345))) : (reg209[(1'h1):(1'h1)] ?
                              (reg121[(3'h7):(2'h3)] ?
                                  ((8'haa) ?
                                      reg371 : reg153) : reg320) : $unsigned({reg43})));
                      reg554 <= ($unsigned($unsigned((+reg142))) ?
                          reg233[(1'h0):(1'h0)] : ((reg340[(1'h0):(1'h0)] ?
                                  (reg165 ?
                                      reg73 : (8'ha7)) : $signed(reg212)) ?
                              reg288 : ($signed((8'ha6)) ?
                                  $signed((8'ha1)) : reg16)));
                      reg555 <= (8'hac);
                      reg556 <= $signed(reg348);
                    end
                  reg557 <= {$signed((8'ha7))};
                  reg558 <= reg98[(3'h5):(1'h0)];
                end
              if ($signed(reg242[(1'h1):(1'h1)]))
                begin
                  if ((-((reg41[(3'h6):(1'h0)] ?
                          reg253[(2'h3):(1'h0)] : $signed((8'h9e))) ?
                      $unsigned(reg26[(2'h2):(1'h1)]) : reg77[(1'h1):(1'h1)])))
                    begin
                      reg559 <= wire10;
                      reg560 <= ((reg289[(4'hf):(4'hb)] ?
                          $unsigned($unsigned(reg124)) : $unsigned($signed(reg238))) << $unsigned(reg363[(3'h4):(2'h3)]));
                    end
                  else
                    begin
                      reg559 <= (!({reg152[(4'hc):(3'h5)]} ^ ((reg197 < reg333) ?
                          reg259[(2'h3):(2'h3)] : $signed(reg69))));
                    end
                  if ($signed($signed((~^reg234[(1'h1):(1'h0)]))))
                    begin
                      reg561 <= reg371[(4'hd):(4'hb)];
                      reg562 <= reg537[(4'ha):(2'h3)];
                      reg563 <= $unsigned($signed((reg212 > (~^reg226))));
                      reg564 <= (&reg358[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg561 <= reg109[(4'h8):(2'h2)];
                      reg562 <= $unsigned($unsigned(reg121[(4'h9):(4'h8)]));
                      reg563 <= $unsigned((~&reg307[(3'h4):(2'h2)]));
                    end
                  if ($unsigned($unsigned(reg322)))
                    begin
                      reg565 <= {reg106[(2'h3):(2'h3)]};
                    end
                  else
                    begin
                      reg565 <= (({$signed(reg78)} <= (~^reg315[(1'h1):(1'h0)])) ?
                          (~reg104[(4'hc):(1'h1)]) : reg193);
                      reg566 <= reg213;
                    end
                end
              else
                begin
                  for (forvar559 = (1'h0); (forvar559 < (1'h0)); forvar559 = (forvar559 + (1'h1)))
                    begin
                      reg560 <= (reg70 ?
                          ((reg275 ?
                                  (reg112 ?
                                      reg103 : (8'had)) : $signed(reg370)) ?
                              {reg17} : reg154) : $signed($signed($signed(reg149))));
                      reg561 <= $unsigned($signed((8'hb5)));
                      reg562 <= (^~reg333);
                    end
                  reg563 <= {reg208};
                  for (forvar564 = (1'h0); (forvar564 < (1'h0)); forvar564 = (forvar564 + (1'h1)))
                    begin
                      reg565 <= reg256;
                    end
                  reg566 <= (reg49 <= ($unsigned($unsigned(reg365)) ?
                      reg360 : reg338));
                end
              for (forvar567 = (1'h0); (forvar567 < (1'h0)); forvar567 = (forvar567 + (1'h1)))
                begin
                  if (reg227[(3'h7):(3'h5)])
                    begin
                      reg568 <= $unsigned(reg156[(3'h4):(2'h2)]);
                      reg569 <= (reg239 ^ $signed($signed({reg114})));
                      reg570 <= (+reg254[(4'he):(3'h6)]);
                      reg571 <= (((reg380[(2'h3):(2'h2)] ?
                              (|(8'hab)) : $unsigned(reg245)) <= ((reg299 ?
                              reg569 : reg55) | (reg131 | (8'hb2)))) ?
                          $unsigned($signed((~^reg372))) : ((~^(reg52 ?
                              reg328 : reg272)) == $unsigned(forvar564[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg568 <= $signed(((^$unsigned(reg186)) >>> $unsigned({wire7})));
                    end
                end
              for (forvar572 = (1'h0); (forvar572 < (1'h0)); forvar572 = (forvar572 + (1'h1)))
                begin
                  if ((reg43 ?
                      ({(reg125 ?
                              reg120 : reg558)} && $unsigned(reg314[(1'h0):(1'h0)])) : $unsigned((-$unsigned(reg17)))))
                    begin
                      reg573 <= {(((~(8'hb3)) || reg173[(4'ha):(2'h3)]) ?
                              ((reg332 ? reg552 : (8'hb1)) ?
                                  reg327[(4'hd):(1'h0)] : (reg293 ?
                                      reg141 : reg90)) : $signed((~^reg564)))};
                      reg574 <= $signed(((reg163[(1'h0):(1'h0)] ?
                          (~^reg163) : $unsigned(reg167)) ^~ {$signed(reg91)}));
                      reg575 <= $unsigned($unsigned(reg280));
                    end
                  else
                    begin
                      reg573 <= $signed(reg208[(3'h5):(2'h3)]);
                      reg574 <= reg52;
                      reg575 <= $signed(((~&{reg561}) - (~&{reg104})));
                      reg576 <= (8'hb7);
                    end
                  for (forvar577 = (1'h0); (forvar577 < (2'h3)); forvar577 = (forvar577 + (1'h1)))
                    begin
                      reg578 <= (~^$unsigned(($unsigned((8'hb2)) * (~reg326))));
                      reg579 <= ({(reg552 ? $unsigned(reg346) : {(8'ha6)})} ?
                          {$signed(reg381)} : reg238[(4'hc):(3'h5)]);
                      reg580 <= reg125;
                      reg581 <= ((8'hab) ?
                          {(^~$unsigned((8'had)))} : reg215[(4'h9):(3'h7)]);
                    end
                  for (forvar582 = (1'h0); (forvar582 < (2'h3)); forvar582 = (forvar582 + (1'h1)))
                    begin
                      reg583 <= $signed($signed((^(reg358 <<< reg40))));
                      reg584 <= (~(($signed((8'hb3)) <<< $signed(reg73)) >= ((reg179 ?
                              (8'hb0) : reg359) ?
                          (8'haa) : $signed(reg346))));
                      reg585 <= $unsigned((reg78 ?
                          (((8'ha9) ?
                              reg42 : reg558) > (reg113 <= (8'hb0))) : (~(reg172 ?
                              reg560 : reg300))));
                      reg586 <= ({(!(~|reg83))} ?
                          (^reg299[(3'h5):(1'h0)]) : reg354);
                    end
                  for (forvar587 = (1'h0); (forvar587 < (2'h2)); forvar587 = (forvar587 + (1'h1)))
                    begin
                      reg588 <= $signed({$unsigned($signed(reg40))});
                      reg589 <= ((reg560[(2'h2):(2'h2)] >> ((&reg371) ?
                          (reg69 ^~ reg216) : ((8'h9e) * (8'h9e)))) > {(~|$unsigned(reg30))});
                      reg590 <= $signed((8'ha5));
                      reg591 <= reg590[(3'h7):(2'h2)];
                    end
                end
            end
        end
      else
        begin
          for (forvar539 = (1'h0); (forvar539 < (1'h0)); forvar539 = (forvar539 + (1'h1)))
            begin
              reg540 <= ($signed((~&$unsigned(reg537))) ?
                  (reg300 ?
                      $unsigned($signed(reg537)) : ((~&reg252) ?
                          reg537[(4'h9):(2'h2)] : forvar542)) : (8'haa));
              if (((reg53 <= $unsigned(reg302[(1'h0):(1'h0)])) + (|(~reg139))))
                begin
                  for (forvar541 = (1'h0); (forvar541 < (2'h3)); forvar541 = (forvar541 + (1'h1)))
                    begin
                      reg542 <= $unsigned(reg557[(3'h7):(3'h5)]);
                      reg543 <= $signed(($signed((wire268 ?
                          (8'h9c) : reg147)) <= (~|wire6)));
                      reg544 <= ((({reg51} ^~ (reg308 ?
                              reg379 : reg591)) | (8'hb8)) ?
                          reg54[(3'h5):(1'h1)] : ({$signed(reg578)} ?
                              $unsigned($unsigned((8'h9d))) : $signed($unsigned(reg308))));
                      reg545 <= (($unsigned((reg315 ? reg151 : reg537)) ?
                          (reg112 - (reg20 != reg66)) : {$signed(reg294)}) && (wire11 * reg226));
                    end
                end
              else
                begin
                  reg541 <= $signed((~$unsigned(reg289[(1'h0):(1'h0)])));
                end
              for (forvar546 = (1'h0); (forvar546 < (1'h0)); forvar546 = (forvar546 + (1'h1)))
                begin
                  if (reg561[(4'h9):(2'h2)])
                    begin
                      reg547 <= (reg379[(2'h2):(1'h1)] ?
                          $unsigned(($unsigned(reg31) ?
                              (&reg301) : (reg241 - reg558))) : $unsigned((8'hb1)));
                      reg548 <= wire6;
                    end
                  else
                    begin
                      reg547 <= (&reg170[(4'ha):(3'h4)]);
                      reg548 <= $unsigned(forvar540);
                      reg549 <= (8'ha7);
                    end
                  for (forvar550 = (1'h0); (forvar550 < (2'h2)); forvar550 = (forvar550 + (1'h1)))
                    begin
                      reg551 <= (reg590[(3'h5):(2'h3)] >> $unsigned((((8'hac) ?
                          wire535 : reg231) > reg75)));
                    end
                  if ($signed({$signed($unsigned(reg562))}))
                    begin
                      reg552 <= (8'ha1);
                      reg553 <= $unsigned((((+reg103) ?
                              wire10 : reg83[(3'h4):(2'h3)]) ?
                          $signed((|reg287)) : $unsigned((8'ha1))));
                    end
                  else
                    begin
                      reg552 <= $signed(reg219[(1'h1):(1'h1)]);
                    end
                end
              for (forvar554 = (1'h0); (forvar554 < (1'h0)); forvar554 = (forvar554 + (1'h1)))
                begin
                  if (reg55)
                    begin
                      reg555 <= ((((~|reg357) > reg52) ?
                          $signed($signed(reg248)) : $signed({reg574})) <= reg41);
                      reg556 <= {forvar540[(3'h5):(3'h4)]};
                      reg557 <= $signed($signed((~((8'ha3) ? reg214 : reg22))));
                      reg558 <= (~&reg241);
                    end
                  else
                    begin
                      reg555 <= {reg186[(1'h1):(1'h0)]};
                      reg556 <= (((reg153 && (reg234 ? (8'h9d) : reg29)) ?
                          {(wire266 <= reg580)} : ((reg257 ? reg225 : reg35) ?
                              (reg258 ?
                                  wire8 : reg566) : (~&reg346))) ^ reg313);
                      reg557 <= ((((8'hb1) ?
                              $unsigned(reg277) : reg352) - (!forvar546[(4'h8):(2'h3)])) ?
                          reg203 : ((&reg558) ?
                              $unsigned((8'haa)) : $signed(reg300[(1'h1):(1'h0)])));
                      reg558 <= $unsigned(reg217);
                    end
                  reg559 <= reg272[(4'hc):(3'h5)];
                  reg560 <= $signed((((8'ha7) ?
                      $unsigned((8'hb3)) : (~&(8'ha2))) < reg545[(1'h1):(1'h1)]));
                end
            end
          for (forvar561 = (1'h0); (forvar561 < (1'h0)); forvar561 = (forvar561 + (1'h1)))
            begin
              reg562 <= $unsigned((reg214[(3'h4):(2'h3)] ?
                  ({reg299} != (reg54 + reg260)) : $signed(reg204[(4'he):(3'h6)])));
              reg563 <= (^~$unsigned(((reg72 ? reg112 : (8'haf)) ?
                  $signed(reg275) : (!reg382))));
              for (forvar564 = (1'h0); (forvar564 < (1'h1)); forvar564 = (forvar564 + (1'h1)))
                begin
                  for (forvar565 = (1'h0); (forvar565 < (2'h2)); forvar565 = (forvar565 + (1'h1)))
                    begin
                      reg566 <= reg224[(3'h4):(2'h3)];
                    end
                  if (($unsigned(reg591[(4'h8):(1'h1)]) ?
                      ({reg113} & (reg142 <<< (8'hae))) : (8'hb2)))
                    begin
                      reg567 <= ((^reg141[(1'h1):(1'h0)]) <= ((^~reg170) > forvar561[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg567 <= (reg574[(1'h0):(1'h0)] - (^($signed(reg61) ?
                          reg78[(1'h0):(1'h0)] : (~^reg112))));
                      reg568 <= reg591[(2'h2):(2'h2)];
                      reg569 <= ((|(8'haf)) <<< reg83[(1'h1):(1'h0)]);
                      reg570 <= reg316;
                    end
                  if ($unsigned($unsigned($unsigned(reg252))))
                    begin
                      reg571 <= $unsigned((8'h9e));
                      reg572 <= (|{$unsigned(reg569[(1'h0):(1'h0)])});
                      reg573 <= $unsigned(reg41[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg571 <= ($signed(reg250[(1'h1):(1'h1)]) ?
                          $unsigned(reg590[(4'h8):(3'h6)]) : (reg76[(1'h1):(1'h1)] ?
                              $signed((reg540 ^~ (8'hb1))) : reg95));
                      reg572 <= reg255;
                      reg573 <= $unsigned($unsigned(reg272[(2'h2):(1'h0)]));
                      reg574 <= $signed($signed(reg311));
                    end
                  for (forvar575 = (1'h0); (forvar575 < (2'h2)); forvar575 = (forvar575 + (1'h1)))
                    begin
                      reg576 <= (^((-(reg30 > reg294)) || (&$signed(forvar551))));
                    end
                end
              for (forvar577 = (1'h0); (forvar577 < (2'h3)); forvar577 = (forvar577 + (1'h1)))
                begin
                  if (reg172[(1'h0):(1'h0)])
                    begin
                      reg578 <= {(~|forvar551)};
                    end
                  else
                    begin
                      reg578 <= ({reg324} ?
                          ($signed(reg218) ?
                              reg368 : (&reg568)) : $signed(((reg83 ?
                                  (8'haf) : reg121) ?
                              ((8'ha2) ? reg293 : reg274) : {(8'hab)})));
                      reg579 <= reg212[(4'h9):(2'h2)];
                      reg580 <= (reg50 ? $signed(reg46) : {reg544});
                    end
                  if ((&(reg258[(3'h4):(3'h4)] == reg112)))
                    begin
                      reg581 <= reg236[(4'h8):(3'h7)];
                    end
                  else
                    begin
                      reg581 <= (reg159[(1'h1):(1'h1)] < $unsigned(reg64));
                      reg582 <= reg218[(1'h0):(1'h0)];
                      reg583 <= reg328[(4'ha):(4'h9)];
                    end
                  if (((~&{forvar565[(2'h2):(2'h2)]}) ?
                      $unsigned((reg51 >= (reg103 ~^ reg259))) : reg104[(4'hd):(4'h9)]))
                    begin
                      reg584 <= $signed((reg297 ?
                          reg246 : ({reg368} || $unsigned(wire7))));
                      reg585 <= reg212[(1'h1):(1'h0)];
                      reg586 <= $unsigned(($unsigned((&reg237)) ?
                          $unsigned($unsigned(reg217)) : (~&$unsigned(reg383))));
                      reg587 <= ({reg128} ?
                          $signed(reg337[(1'h1):(1'h1)]) : $unsigned(($signed(reg362) ?
                              {(8'haf)} : ((8'hb3) - reg160))));
                    end
                  else
                    begin
                      reg584 <= reg307[(1'h1):(1'h1)];
                    end
                  for (forvar588 = (1'h0); (forvar588 < (2'h2)); forvar588 = (forvar588 + (1'h1)))
                    begin
                      reg589 <= reg321[(2'h3):(2'h2)];
                      reg590 <= reg82;
                      reg591 <= (8'hae);
                      reg592 <= (~|($signed((reg586 >= reg329)) ?
                          ($unsigned(reg155) * (reg152 ?
                              reg186 : reg589)) : $unsigned((&reg88))));
                    end
                end
            end
        end
      for (forvar593 = (1'h0); (forvar593 < (1'h1)); forvar593 = (forvar593 + (1'h1)))
        begin
          for (forvar594 = (1'h0); (forvar594 < (1'h0)); forvar594 = (forvar594 + (1'h1)))
            begin
              reg595 <= {(reg587 ?
                      ((reg338 << forvar567) ?
                          {reg307} : $unsigned(reg84)) : (reg181 < $signed(forvar541)))};
              for (forvar596 = (1'h0); (forvar596 < (2'h2)); forvar596 = (forvar596 + (1'h1)))
                begin
                  reg597 <= ((({reg299} <= $signed(reg359)) && $unsigned(reg343[(3'h6):(3'h5)])) ?
                      forvar541[(3'h4):(1'h1)] : $signed(((wire265 ?
                          reg36 : reg131) != (reg59 ? (8'hae) : reg340))));
                  for (forvar598 = (1'h0); (forvar598 < (1'h1)); forvar598 = (forvar598 + (1'h1)))
                    begin
                      reg599 <= $unsigned((-(|(^reg592))));
                      reg600 <= $signed(reg219[(1'h0):(1'h0)]);
                    end
                  if ($unsigned({$signed($signed((8'hb6)))}))
                    begin
                      reg601 <= (+$signed((~^$signed(reg45))));
                    end
                  else
                    begin
                      reg601 <= (&reg120[(1'h0):(1'h0)]);
                      reg602 <= (8'hb1);
                      reg603 <= {reg179};
                      reg604 <= $unsigned($unsigned(forvar572));
                    end
                  for (forvar605 = (1'h0); (forvar605 < (2'h3)); forvar605 = (forvar605 + (1'h1)))
                    begin
                      reg606 <= {$unsigned(reg576)};
                      reg607 <= {(reg289 - reg286)};
                      reg608 <= reg65;
                    end
                end
              for (forvar609 = (1'h0); (forvar609 < (2'h3)); forvar609 = (forvar609 + (1'h1)))
                begin
                  for (forvar610 = (1'h0); (forvar610 < (1'h1)); forvar610 = (forvar610 + (1'h1)))
                    begin
                      reg611 <= $signed((~^(wire9[(3'h5):(1'h1)] < (reg46 ?
                          reg365 : reg20))));
                    end
                  for (forvar612 = (1'h0); (forvar612 < (1'h1)); forvar612 = (forvar612 + (1'h1)))
                    begin
                      reg613 <= $unsigned((($signed(reg54) ?
                              (reg95 ? (8'hb2) : reg562) : (~reg604)) ?
                          reg203[(3'h7):(1'h1)] : {(reg263 ?
                                  wire266 : reg301)}));
                    end
                  for (forvar614 = (1'h0); (forvar614 < (2'h3)); forvar614 = (forvar614 + (1'h1)))
                    begin
                      reg615 <= (8'ha0);
                      reg616 <= ((8'ha8) ?
                          (8'hb1) : ($signed({(8'hb8)}) ?
                              (reg139 ?
                                  (~^reg380) : $unsigned(reg224)) : {$signed(reg586)}));
                    end
                end
              if ($signed($signed($signed(reg581[(1'h1):(1'h0)]))))
                begin
                  reg617 <= ($signed(reg16[(3'h4):(1'h1)]) ?
                      ($unsigned(reg556) ?
                          {(reg90 | reg371)} : $signed(reg275[(1'h1):(1'h0)])) : (($signed(reg275) >> $signed(reg69)) ?
                          $signed(reg37) : $unsigned(reg551)));
                  reg618 <= $unsigned($signed((+((8'ha4) ? reg141 : reg181))));
                  if ($unsigned($signed(reg306[(2'h3):(1'h0)])))
                    begin
                      reg619 <= $unsigned($signed((8'hb1)));
                      reg620 <= {(reg559[(2'h3):(2'h2)] < wire265[(3'h5):(3'h5)])};
                      reg621 <= reg134[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg619 <= ((reg167 ^~ $unsigned(wire8[(1'h1):(1'h1)])) <= reg226[(3'h7):(2'h2)]);
                      reg620 <= (reg261 ?
                          {$unsigned(reg231)} : reg107[(3'h4):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar617 = (1'h0); (forvar617 < (2'h3)); forvar617 = (forvar617 + (1'h1)))
                    begin
                      reg618 <= ((8'hac) && $unsigned(forvar582[(2'h2):(1'h0)]));
                    end
                  for (forvar619 = (1'h0); (forvar619 < (1'h0)); forvar619 = (forvar619 + (1'h1)))
                    begin
                      reg620 <= ((-(!reg156)) >= (~^reg313));
                      reg621 <= $unsigned($signed(reg548));
                      reg622 <= ($unsigned(reg131[(4'h8):(1'h1)]) ?
                          $unsigned($signed({(8'ha2)})) : $unsigned(({(8'had)} >>> {reg43})));
                    end
                  for (forvar623 = (1'h0); (forvar623 < (1'h0)); forvar623 = (forvar623 + (1'h1)))
                    begin
                      reg624 <= reg270[(3'h7):(3'h7)];
                      reg625 <= reg83;
                    end
                  reg626 <= reg44[(1'h0):(1'h0)];
                end
            end
        end
    end
  assign wire627 = $signed($unsigned(reg49));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module385  (y, clk, wire389, wire388, wire387, wire386);
  output wire [(32'h642):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire389;
  input wire signed [(5'h10):(1'h0)] wire388;
  input wire [(4'hf):(1'h0)] wire387;
  input wire signed [(2'h3):(1'h0)] wire386;
  wire signed [(2'h2):(1'h0)] wire534;
  wire [(4'he):(1'h0)] wire444;
  wire signed [(3'h4):(1'h0)] wire391;
  wire [(4'hf):(1'h0)] wire390;
  reg signed [(4'h9):(1'h0)] reg510 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg509 = (1'h0);
  reg [(4'hc):(1'h0)] reg504 = (1'h0);
  reg [(4'h9):(1'h0)] reg503 = (1'h0);
  reg [(4'he):(1'h0)] reg500 = (1'h0);
  reg [(5'h10):(1'h0)] reg533 = (1'h0);
  reg [(4'hd):(1'h0)] reg532 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg531 = (1'h0);
  reg [(3'h5):(1'h0)] reg530 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg529 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg528 = (1'h0);
  reg [(4'hc):(1'h0)] reg527 = (1'h0);
  reg [(5'h10):(1'h0)] reg526 = (1'h0);
  reg [(4'he):(1'h0)] reg525 = (1'h0);
  reg [(4'h8):(1'h0)] reg523 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg521 = (1'h0);
  reg [(3'h7):(1'h0)] reg520 = (1'h0);
  reg [(4'ha):(1'h0)] reg519 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg518 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg517 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg516 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg515 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg514 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg513 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg512 = (1'h0);
  reg [(5'h10):(1'h0)] reg511 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg508 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg507 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg506 = (1'h0);
  reg [(3'h6):(1'h0)] reg505 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg502 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg501 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg499 = (1'h0);
  reg signed [(4'he):(1'h0)] reg498 = (1'h0);
  reg [(4'hf):(1'h0)] reg496 = (1'h0);
  reg [(3'h6):(1'h0)] reg495 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg494 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg492 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg487 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg475 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg477 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg474 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg470 = (1'h0);
  reg [(4'he):(1'h0)] reg493 = (1'h0);
  reg [(5'h10):(1'h0)] reg491 = (1'h0);
  reg [(3'h5):(1'h0)] reg490 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg489 = (1'h0);
  reg [(3'h6):(1'h0)] reg488 = (1'h0);
  reg signed [(4'he):(1'h0)] reg486 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg485 = (1'h0);
  reg [(4'h8):(1'h0)] reg484 = (1'h0);
  reg [(4'h9):(1'h0)] reg483 = (1'h0);
  reg [(4'hf):(1'h0)] reg481 = (1'h0);
  reg signed [(4'he):(1'h0)] reg479 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg478 = (1'h0);
  reg [(4'hc):(1'h0)] reg476 = (1'h0);
  reg [(2'h3):(1'h0)] reg473 = (1'h0);
  reg signed [(4'he):(1'h0)] reg472 = (1'h0);
  reg [(5'h10):(1'h0)] reg471 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg469 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg464 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg468 = (1'h0);
  reg [(4'hc):(1'h0)] reg467 = (1'h0);
  reg [(3'h6):(1'h0)] reg466 = (1'h0);
  reg [(4'hf):(1'h0)] reg465 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg463 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg461 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg460 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg459 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg458 = (1'h0);
  reg signed [(4'he):(1'h0)] reg456 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg455 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg454 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg452 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg451 = (1'h0);
  reg [(4'h8):(1'h0)] reg450 = (1'h0);
  reg [(3'h5):(1'h0)] reg446 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg398 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg397 = (1'h0);
  reg [(4'hb):(1'h0)] reg394 = (1'h0);
  reg [(4'h9):(1'h0)] reg392 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg443 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg442 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg441 = (1'h0);
  reg [(3'h4):(1'h0)] reg438 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg437 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg435 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg434 = (1'h0);
  reg [(4'hf):(1'h0)] reg433 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg432 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg431 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg429 = (1'h0);
  reg [(5'h10):(1'h0)] reg428 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg427 = (1'h0);
  reg [(4'hf):(1'h0)] reg426 = (1'h0);
  reg [(3'h4):(1'h0)] reg425 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg423 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg421 = (1'h0);
  reg [(3'h4):(1'h0)] reg420 = (1'h0);
  reg [(4'hc):(1'h0)] reg418 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg417 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg416 = (1'h0);
  reg [(3'h4):(1'h0)] reg415 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg414 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg413 = (1'h0);
  reg [(2'h3):(1'h0)] reg410 = (1'h0);
  reg [(4'ha):(1'h0)] reg402 = (1'h0);
  reg [(3'h5):(1'h0)] reg409 = (1'h0);
  reg [(2'h2):(1'h0)] reg408 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg407 = (1'h0);
  reg [(4'hc):(1'h0)] reg406 = (1'h0);
  reg [(3'h6):(1'h0)] reg405 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg404 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg401 = (1'h0);
  reg [(3'h4):(1'h0)] reg400 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg399 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg396 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar507 = (1'h0);
  reg [(4'hb):(1'h0)] forvar502 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar524 = (1'h0);
  reg [(3'h5):(1'h0)] forvar522 = (1'h0);
  reg [(3'h7):(1'h0)] forvar510 = (1'h0);
  reg [(2'h2):(1'h0)] forvar509 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar504 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar503 = (1'h0);
  reg [(4'hc):(1'h0)] forvar500 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar497 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar493 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar488 = (1'h0);
  reg [(4'hd):(1'h0)] forvar483 = (1'h0);
  reg [(3'h7):(1'h0)] forvar469 = (1'h0);
  reg [(4'h8):(1'h0)] forvar465 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar492 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar487 = (1'h0);
  reg [(3'h6):(1'h0)] forvar482 = (1'h0);
  reg [(2'h2):(1'h0)] forvar480 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar477 = (1'h0);
  reg [(2'h3):(1'h0)] forvar475 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar474 = (1'h0);
  reg [(4'ha):(1'h0)] forvar470 = (1'h0);
  reg [(3'h6):(1'h0)] forvar466 = (1'h0);
  reg [(4'h9):(1'h0)] forvar463 = (1'h0);
  reg [(4'hb):(1'h0)] forvar464 = (1'h0);
  reg [(4'h9):(1'h0)] forvar462 = (1'h0);
  reg [(3'h6):(1'h0)] forvar457 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar449 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar448 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar447 = (1'h0);
  reg [(5'h10):(1'h0)] forvar445 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar403 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar395 = (1'h0);
  reg [(4'h9):(1'h0)] forvar440 = (1'h0);
  reg [(4'he):(1'h0)] forvar439 = (1'h0);
  reg [(3'h6):(1'h0)] forvar436 = (1'h0);
  reg [(4'h8):(1'h0)] forvar430 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar424 = (1'h0);
  reg [(5'h10):(1'h0)] forvar422 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar419 = (1'h0);
  reg [(3'h6):(1'h0)] forvar414 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar412 = (1'h0);
  reg [(4'hd):(1'h0)] forvar411 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar408 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar402 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar398 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar397 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar394 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar393 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar392 = (1'h0);
  assign y = {wire534,
                 wire444,
                 wire391,
                 wire390,
                 reg510,
                 reg509,
                 reg504,
                 reg503,
                 reg500,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 reg523,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 reg512,
                 reg511,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg502,
                 reg501,
                 reg499,
                 reg498,
                 reg496,
                 reg495,
                 reg494,
                 reg492,
                 reg487,
                 reg475,
                 reg477,
                 reg474,
                 reg470,
                 reg493,
                 reg491,
                 reg490,
                 reg489,
                 reg488,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg481,
                 reg479,
                 reg478,
                 reg476,
                 reg473,
                 reg472,
                 reg471,
                 reg469,
                 reg464,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg463,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg446,
                 reg398,
                 reg397,
                 reg394,
                 reg392,
                 reg443,
                 reg442,
                 reg441,
                 reg438,
                 reg437,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 reg425,
                 reg423,
                 reg421,
                 reg420,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg410,
                 reg402,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg401,
                 reg400,
                 reg399,
                 reg396,
                 reg395,
                 forvar507,
                 forvar502,
                 forvar524,
                 forvar522,
                 forvar510,
                 forvar509,
                 forvar504,
                 forvar503,
                 forvar500,
                 forvar497,
                 forvar493,
                 forvar488,
                 forvar483,
                 forvar469,
                 forvar465,
                 forvar492,
                 forvar487,
                 forvar482,
                 forvar480,
                 forvar477,
                 forvar475,
                 forvar474,
                 forvar470,
                 forvar466,
                 forvar463,
                 forvar464,
                 forvar462,
                 forvar457,
                 forvar449,
                 forvar448,
                 forvar447,
                 forvar445,
                 forvar403,
                 forvar395,
                 forvar440,
                 forvar439,
                 forvar436,
                 forvar430,
                 forvar424,
                 forvar422,
                 forvar419,
                 forvar414,
                 forvar412,
                 forvar411,
                 forvar408,
                 forvar402,
                 forvar398,
                 forvar397,
                 forvar394,
                 forvar393,
                 forvar392,
                 (1'h0)};
  assign wire390 = $unsigned(wire386[(2'h2):(1'h1)]);
  assign wire391 = (wire386 ?
                       $signed(($signed(wire387) ?
                           {wire389} : wire386)) : {$unsigned((wire390 <= wire388))});
  always
    @(posedge clk) begin
      if ((($unsigned((wire388 ? wire390 : wire387)) ?
          wire386[(1'h1):(1'h0)] : $signed($unsigned(wire390))) <<< (!$unsigned(wire390))))
        begin
          for (forvar392 = (1'h0); (forvar392 < (1'h1)); forvar392 = (forvar392 + (1'h1)))
            begin
              for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
                begin
                  for (forvar394 = (1'h0); (forvar394 < (1'h0)); forvar394 = (forvar394 + (1'h1)))
                    begin
                      reg395 <= (^~$signed({forvar393[(3'h6):(2'h3)]}));
                      reg396 <= (wire386[(2'h3):(1'h1)] ?
                          $unsigned((8'hba)) : $unsigned($signed($unsigned(reg395))));
                    end
                end
              for (forvar397 = (1'h0); (forvar397 < (2'h3)); forvar397 = (forvar397 + (1'h1)))
                begin
                  for (forvar398 = (1'h0); (forvar398 < (1'h0)); forvar398 = (forvar398 + (1'h1)))
                    begin
                      reg399 <= (((|$signed(wire386)) ^ (8'hac)) > $signed((8'ha7)));
                    end
                  reg400 <= (forvar394 - forvar392[(2'h2):(1'h0)]);
                  reg401 <= ($unsigned((8'ha5)) << wire388);
                end
              if ($unsigned($unsigned($signed((forvar398 ? reg396 : wire387)))))
                begin
                  for (forvar402 = (1'h0); (forvar402 < (2'h3)); forvar402 = (forvar402 + (1'h1)))
                    begin
                      reg403 <= reg400[(3'h4):(1'h1)];
                      reg404 <= $unsigned($signed($unsigned((reg401 >= reg401))));
                      reg405 <= (wire390 ?
                          $unsigned($unsigned(wire390[(4'hd):(1'h1)])) : reg395[(2'h2):(1'h0)]);
                    end
                  if ($signed($signed($signed(reg405))))
                    begin
                      reg406 <= (forvar397 >> reg404[(3'h5):(3'h4)]);
                    end
                  else
                    begin
                      reg406 <= forvar394[(2'h3):(2'h2)];
                      reg407 <= $unsigned($signed(($signed(reg406) == ((8'ha1) ^~ (8'hb6)))));
                      reg408 <= reg406;
                      reg409 <= $signed((forvar397[(3'h4):(2'h3)] ?
                          ((reg395 ^~ forvar397) || $signed(wire390)) : (8'hb1)));
                    end
                end
              else
                begin
                  reg402 <= $signed(reg405);
                  reg403 <= (!((8'h9e) ?
                      (reg403[(1'h1):(1'h0)] ?
                          reg396 : (8'ha8)) : reg409[(1'h1):(1'h0)]));
                  if (($signed($signed((reg403 ? wire386 : wire389))) ?
                      reg402[(2'h2):(2'h2)] : (-$signed(reg403[(2'h3):(2'h2)]))))
                    begin
                      reg404 <= ($signed((-{wire386})) ?
                          ((&(wire388 ^ wire389)) ?
                              forvar397[(3'h4):(1'h0)] : (reg404 ?
                                  ((8'ha7) ? (8'ha2) : (8'hac)) : (forvar393 ?
                                      forvar397 : wire391))) : $unsigned($unsigned(wire388)));
                    end
                  else
                    begin
                      reg404 <= $signed($unsigned($signed((wire389 ?
                          (8'hb0) : reg401))));
                      reg405 <= (~|wire388);
                      reg406 <= ($unsigned($unsigned(reg400)) ?
                          (+(8'ha3)) : ({(wire386 == wire388)} + forvar394[(3'h4):(1'h1)]));
                      reg407 <= reg401;
                    end
                  for (forvar408 = (1'h0); (forvar408 < (2'h2)); forvar408 = (forvar408 + (1'h1)))
                    begin
                      reg409 <= {reg402};
                      reg410 <= (($signed(reg396) >= ($unsigned(wire388) ?
                          $unsigned(reg408) : $unsigned((8'hb3)))) - ((reg401[(3'h5):(2'h2)] ?
                          $signed(reg408) : (reg403 ?
                              forvar392 : forvar393)) != $unsigned($signed(wire390))));
                    end
                end
            end
          for (forvar411 = (1'h0); (forvar411 < (2'h2)); forvar411 = (forvar411 + (1'h1)))
            begin
              if ((reg399 < ({(~^forvar402)} - forvar397[(4'h8):(3'h6)])))
                begin
                  for (forvar412 = (1'h0); (forvar412 < (2'h3)); forvar412 = (forvar412 + (1'h1)))
                    begin
                      reg413 <= $signed($unsigned({$signed(forvar398)}));
                      reg414 <= forvar408[(3'h7):(3'h7)];
                      reg415 <= ((!{{(8'hb6)}}) ?
                          $signed((^~(~&forvar397))) : $signed((~|(-wire391))));
                    end
                  reg416 <= $unsigned(forvar392);
                  reg417 <= $unsigned(reg396[(3'h7):(2'h2)]);
                end
              else
                begin
                  for (forvar412 = (1'h0); (forvar412 < (1'h0)); forvar412 = (forvar412 + (1'h1)))
                    begin
                      reg413 <= {{(8'hae)}};
                    end
                  for (forvar414 = (1'h0); (forvar414 < (1'h1)); forvar414 = (forvar414 + (1'h1)))
                    begin
                      reg415 <= (~(|(8'hb7)));
                      reg416 <= reg402;
                      reg417 <= forvar392;
                      reg418 <= ((^~$signed((~^reg413))) ?
                          (~^{$unsigned(reg395)}) : (^$unsigned(reg400[(2'h3):(2'h2)])));
                    end
                  for (forvar419 = (1'h0); (forvar419 < (1'h1)); forvar419 = (forvar419 + (1'h1)))
                    begin
                      reg420 <= $signed(((^~(wire387 - forvar419)) < ($unsigned(wire386) && $unsigned(wire387))));
                      reg421 <= (+((~&reg414) ?
                          (8'hb0) : $signed(reg396[(3'h7):(3'h4)])));
                    end
                  for (forvar422 = (1'h0); (forvar422 < (1'h1)); forvar422 = (forvar422 + (1'h1)))
                    begin
                      reg423 <= (8'ha4);
                    end
                end
              for (forvar424 = (1'h0); (forvar424 < (2'h3)); forvar424 = (forvar424 + (1'h1)))
                begin
                  reg425 <= ((({(8'hb4)} >> reg410) ?
                          $signed({reg414}) : (reg407[(1'h1):(1'h1)] <= $signed(forvar424))) ?
                      ({(reg401 && wire389)} ?
                          (forvar412[(2'h2):(1'h0)] ?
                              (^~wire386) : reg416[(1'h1):(1'h0)]) : ((!(8'hb9)) <= (reg408 ?
                              (8'hac) : forvar393))) : {(^~(reg395 ?
                              reg418 : (8'ha0)))});
                  if ((~$unsigned((~^(wire390 - forvar422)))))
                    begin
                      reg426 <= $signed($unsigned(($unsigned(reg415) ?
                          $unsigned(forvar424) : wire390)));
                    end
                  else
                    begin
                      reg426 <= ($unsigned({(forvar419 <<< reg407)}) || reg403);
                      reg427 <= $signed($unsigned(({forvar424} ^~ reg420[(2'h2):(1'h1)])));
                      reg428 <= ((reg409 + forvar408) & reg426[(1'h1):(1'h0)]);
                      reg429 <= ($signed($unsigned(forvar393[(1'h0):(1'h0)])) ?
                          reg409 : (forvar393 && reg417));
                    end
                  for (forvar430 = (1'h0); (forvar430 < (1'h1)); forvar430 = (forvar430 + (1'h1)))
                    begin
                      reg431 <= (((~|$unsigned(forvar430)) + reg406[(3'h7):(3'h7)]) == forvar392);
                      reg432 <= $signed(forvar414);
                      reg433 <= $signed((forvar394 ~^ (^~reg413[(1'h1):(1'h0)])));
                    end
                  if (({(8'hb1)} ~^ forvar422))
                    begin
                      reg434 <= reg410;
                      reg435 <= reg425[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg434 <= reg416;
                      reg435 <= $unsigned((~^reg427[(3'h4):(3'h4)]));
                    end
                end
            end
          for (forvar436 = (1'h0); (forvar436 < (2'h3)); forvar436 = (forvar436 + (1'h1)))
            begin
              reg437 <= (forvar402[(4'h8):(3'h5)] ?
                  (8'hb2) : ($unsigned(forvar419[(1'h1):(1'h0)]) ?
                      {reg428[(1'h0):(1'h0)]} : $signed($unsigned(reg400))));
              reg438 <= {(~|$unsigned($unsigned(wire390)))};
              for (forvar439 = (1'h0); (forvar439 < (1'h1)); forvar439 = (forvar439 + (1'h1)))
                begin
                  for (forvar440 = (1'h0); (forvar440 < (1'h1)); forvar440 = (forvar440 + (1'h1)))
                    begin
                      reg441 <= ({reg415[(1'h1):(1'h0)]} ?
                          $signed(reg432) : (8'haa));
                    end
                  reg442 <= forvar394;
                end
              reg443 <= (((((8'hb0) ?
                      forvar414 : forvar440) & $signed(reg399)) > (reg400 ?
                      (forvar419 ? forvar398 : reg408) : reg426)) ?
                  $unsigned((reg403[(1'h0):(1'h0)] | (&(8'hb8)))) : ((reg405[(3'h6):(3'h6)] >= {(8'hab)}) & reg415[(3'h4):(2'h3)]));
            end
        end
      else
        begin
          reg392 <= {(|(|((8'hb2) ? forvar408 : wire387)))};
          for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 <= reg416;
              if (reg437)
                begin
                  for (forvar395 = (1'h0); (forvar395 < (1'h0)); forvar395 = (forvar395 + (1'h1)))
                    begin
                      reg396 <= $signed(reg410[(1'h0):(1'h0)]);
                      reg397 <= reg421[(4'h8):(3'h6)];
                    end
                  for (forvar398 = (1'h0); (forvar398 < (1'h1)); forvar398 = (forvar398 + (1'h1)))
                    begin
                      reg399 <= (^~forvar398);
                      reg400 <= (8'hba);
                    end
                  if ($unsigned(wire390[(4'he):(4'hc)]))
                    begin
                      reg401 <= $unsigned(reg394);
                      reg402 <= (!$signed((~&$unsigned((8'hb1)))));
                    end
                  else
                    begin
                      reg401 <= wire391[(1'h0):(1'h0)];
                      reg402 <= reg392[(3'h5):(2'h3)];
                    end
                  for (forvar403 = (1'h0); (forvar403 < (2'h2)); forvar403 = (forvar403 + (1'h1)))
                    begin
                      reg404 <= ($unsigned(((reg421 ?
                              reg433 : wire391) & $signed((8'ha7)))) ?
                          (((|forvar414) ? wire387 : forvar419) ?
                              (|(forvar440 | reg399)) : $unsigned((&(8'hb4)))) : reg407[(1'h1):(1'h1)]);
                      reg405 <= $signed(((reg394[(1'h1):(1'h1)] && $unsigned(reg432)) > {(wire391 ?
                              (8'ha0) : reg441)}));
                      reg406 <= {$signed($signed(reg423[(4'h8):(3'h6)]))};
                    end
                end
              else
                begin
                  reg395 <= ({((forvar424 + reg421) ^~ $unsigned(reg401))} << (~|(+wire388[(4'hb):(3'h4)])));
                  reg396 <= (^~(8'haa));
                  for (forvar397 = (1'h0); (forvar397 < (2'h2)); forvar397 = (forvar397 + (1'h1)))
                    begin
                      reg398 <= $signed(reg443[(2'h3):(1'h0)]);
                      reg399 <= forvar408[(2'h3):(2'h2)];
                    end
                end
            end
          reg407 <= $signed((~&wire391));
        end
    end
  assign wire444 = (reg406[(3'h4):(2'h3)] ?
                       (reg423[(3'h7):(3'h7)] ?
                           ($unsigned(reg438) ?
                               (reg400 ? reg429 : (8'hb8)) : (reg425 ?
                                   wire388 : reg413)) : $unsigned(((8'haa) ?
                               reg435 : wire386))) : (~&wire388[(1'h1):(1'h1)]));
  always
    @(posedge clk) begin
      for (forvar445 = (1'h0); (forvar445 < (1'h0)); forvar445 = (forvar445 + (1'h1)))
        begin
          reg446 <= $unsigned(reg420[(2'h2):(1'h0)]);
        end
      for (forvar447 = (1'h0); (forvar447 < (2'h3)); forvar447 = (forvar447 + (1'h1)))
        begin
          for (forvar448 = (1'h0); (forvar448 < (1'h1)); forvar448 = (forvar448 + (1'h1)))
            begin
              for (forvar449 = (1'h0); (forvar449 < (2'h2)); forvar449 = (forvar449 + (1'h1)))
                begin
                  if (reg402)
                    begin
                      reg450 <= $signed($signed(reg395[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg450 <= {forvar447[(3'h5):(2'h3)]};
                    end
                end
              if (($unsigned(((reg395 ? reg417 : reg404) ?
                      (reg435 || reg446) : reg410)) ?
                  reg403 : (~^wire444)))
                begin
                  reg451 <= (reg394[(4'h8):(3'h6)] * $unsigned($unsigned(reg402)));
                end
              else
                begin
                  if ((reg443 >> reg434))
                    begin
                      reg451 <= $unsigned((reg427[(3'h5):(3'h4)] + reg405[(3'h5):(1'h0)]));
                      reg452 <= (!wire387[(1'h1):(1'h1)]);
                      reg453 <= {$unsigned(reg426)};
                      reg454 <= (8'h9c);
                    end
                  else
                    begin
                      reg451 <= $unsigned({reg428[(3'h4):(1'h1)]});
                      reg452 <= (~|reg410);
                      reg453 <= reg396[(2'h3):(2'h2)];
                      reg454 <= (~($signed(forvar445) >>> (~&reg441[(1'h1):(1'h1)])));
                    end
                  if ({forvar445})
                    begin
                      reg455 <= reg402[(4'h9):(3'h5)];
                      reg456 <= (reg426[(2'h2):(1'h1)] ?
                          (-$unsigned((reg396 ?
                              reg408 : (8'ha2)))) : ((~|(^~reg427)) ~^ reg418[(3'h6):(1'h1)]));
                    end
                  else
                    begin
                      reg455 <= (8'hae);
                      reg456 <= ($signed((|(reg452 ?
                          (8'ha8) : wire387))) == $signed($unsigned((reg432 <<< reg407))));
                    end
                  for (forvar457 = (1'h0); (forvar457 < (1'h1)); forvar457 = (forvar457 + (1'h1)))
                    begin
                      reg458 <= reg421[(3'h7):(3'h7)];
                      reg459 <= (((|reg423[(2'h2):(1'h1)]) ?
                          (wire388[(5'h10):(4'hd)] ?
                              (reg415 ?
                                  reg420 : reg427) : reg450) : reg410[(2'h3):(1'h1)]) < wire388[(3'h7):(3'h5)]);
                      reg460 <= (((|{(8'h9f)}) > $unsigned((reg399 || reg402))) ?
                          $unsigned($signed((~reg413))) : ($unsigned(reg414) ?
                              {(reg442 | (8'ha1))} : $signed(reg431[(1'h0):(1'h0)])));
                      reg461 <= ((|reg398) ?
                          reg429 : (reg443 * (reg397[(3'h5):(2'h3)] > reg455[(2'h2):(1'h0)])));
                    end
                end
            end
        end
      if ($unsigned(({$unsigned(reg399)} >= reg435[(2'h2):(1'h0)])))
        begin
          for (forvar462 = (1'h0); (forvar462 < (1'h1)); forvar462 = (forvar462 + (1'h1)))
            begin
              if (((~&$signed((wire444 << reg455))) ^~ ($signed(((8'ha5) | forvar449)) ?
                  {$unsigned(reg438)} : (~&reg410))))
                begin
                  reg463 <= {$unsigned((reg459 ^ reg458))};
                  for (forvar464 = (1'h0); (forvar464 < (1'h0)); forvar464 = (forvar464 + (1'h1)))
                    begin
                      reg465 <= forvar448[(1'h1):(1'h1)];
                      reg466 <= (+$signed(wire391[(2'h3):(1'h1)]));
                      reg467 <= reg452;
                      reg468 <= wire390[(3'h6):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar463 = (1'h0); (forvar463 < (1'h1)); forvar463 = (forvar463 + (1'h1)))
                    begin
                      reg464 <= (reg395[(1'h0):(1'h0)] <= forvar457[(2'h3):(2'h3)]);
                      reg465 <= $unsigned(({(~&forvar457)} ?
                          reg452[(1'h0):(1'h0)] : reg425[(2'h3):(2'h3)]));
                    end
                  for (forvar466 = (1'h0); (forvar466 < (2'h3)); forvar466 = (forvar466 + (1'h1)))
                    begin
                      reg467 <= ((reg421[(3'h6):(1'h0)] <<< ((^reg435) <= ((8'hac) ^~ wire391))) | $signed($signed($unsigned(reg438))));
                      reg468 <= forvar448[(1'h0):(1'h0)];
                      reg469 <= reg459;
                    end
                  for (forvar470 = (1'h0); (forvar470 < (2'h3)); forvar470 = (forvar470 + (1'h1)))
                    begin
                      reg471 <= (($signed($unsigned(reg437)) ^~ (reg420[(2'h3):(1'h0)] >> reg405)) < $signed(((reg453 ?
                              reg401 : reg406) ?
                          {reg427} : {reg395})));
                      reg472 <= (^~$signed((reg414 ?
                          ((8'ha3) ? wire389 : reg459) : $signed(reg469))));
                    end
                end
              reg473 <= forvar449;
              for (forvar474 = (1'h0); (forvar474 < (1'h1)); forvar474 = (forvar474 + (1'h1)))
                begin
                  for (forvar475 = (1'h0); (forvar475 < (2'h2)); forvar475 = (forvar475 + (1'h1)))
                    begin
                      reg476 <= reg396;
                    end
                  for (forvar477 = (1'h0); (forvar477 < (2'h2)); forvar477 = (forvar477 + (1'h1)))
                    begin
                      reg478 <= $signed({reg400[(1'h1):(1'h0)]});
                    end
                  reg479 <= $unsigned((reg429 >> ({forvar464} * (+(8'ha6)))));
                  for (forvar480 = (1'h0); (forvar480 < (1'h1)); forvar480 = (forvar480 + (1'h1)))
                    begin
                      reg481 <= ($signed((reg397[(3'h6):(3'h4)] >>> (^reg446))) || reg404[(4'hd):(3'h5)]);
                    end
                end
              for (forvar482 = (1'h0); (forvar482 < (2'h3)); forvar482 = (forvar482 + (1'h1)))
                begin
                  if ((&{$unsigned(reg417)}))
                    begin
                      reg483 <= $signed(reg429[(4'h9):(3'h5)]);
                    end
                  else
                    begin
                      reg483 <= (^~reg450[(3'h4):(3'h4)]);
                      reg484 <= $unsigned({((reg464 ?
                              reg471 : (8'hb7)) + wire390)});
                    end
                  if (forvar449[(3'h6):(1'h0)])
                    begin
                      reg485 <= $signed(($unsigned(((8'hb9) == (8'ha3))) ?
                          $unsigned($unsigned((8'hb5))) : reg392[(4'h8):(3'h5)]));
                      reg486 <= $unsigned($signed((~|{forvar474})));
                    end
                  else
                    begin
                      reg485 <= (8'ha6);
                      reg486 <= (-({(reg431 << reg396)} <<< ((reg437 <<< (8'ha5)) ?
                          reg443[(3'h6):(3'h4)] : ((8'hab) ?
                              (8'hb6) : reg476))));
                    end
                  for (forvar487 = (1'h0); (forvar487 < (2'h2)); forvar487 = (forvar487 + (1'h1)))
                    begin
                      reg488 <= reg425;
                      reg489 <= $unsigned(forvar470[(1'h1):(1'h0)]);
                      reg490 <= reg421[(1'h0):(1'h0)];
                      reg491 <= ($signed($signed((reg433 ? reg403 : (8'ha7)))) ?
                          ((~^$signed(reg415)) > $unsigned((8'ha6))) : $unsigned((forvar482 ^~ reg434[(1'h0):(1'h0)])));
                    end
                  for (forvar492 = (1'h0); (forvar492 < (1'h1)); forvar492 = (forvar492 + (1'h1)))
                    begin
                      reg493 <= $signed(reg467[(4'hb):(4'h9)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar462 = (1'h0); (forvar462 < (1'h0)); forvar462 = (forvar462 + (1'h1)))
            begin
              for (forvar463 = (1'h0); (forvar463 < (1'h1)); forvar463 = (forvar463 + (1'h1)))
                begin
                  reg464 <= $unsigned(reg398);
                  for (forvar465 = (1'h0); (forvar465 < (1'h0)); forvar465 = (forvar465 + (1'h1)))
                    begin
                      reg466 <= (reg460 ?
                          $unsigned($unsigned({forvar480})) : (8'had));
                      reg467 <= reg402;
                      reg468 <= $signed((forvar487 ^ ((reg452 ?
                          reg432 : reg489) & $signed(forvar480))));
                    end
                end
              for (forvar469 = (1'h0); (forvar469 < (2'h3)); forvar469 = (forvar469 + (1'h1)))
                begin
                  if (((~|$unsigned((~|forvar466))) >> $unsigned($unsigned(forvar469[(2'h3):(1'h0)]))))
                    begin
                      reg470 <= $signed(reg402);
                      reg471 <= ((forvar465[(3'h5):(3'h4)] ?
                              $unsigned((~&reg394)) : reg432) ?
                          reg421[(3'h5):(1'h1)] : {(~^reg438)});
                      reg472 <= reg426;
                    end
                  else
                    begin
                      reg470 <= reg392;
                      reg471 <= $unsigned($signed(forvar466));
                    end
                  reg473 <= $signed({(8'hb7)});
                end
              if ($unsigned(reg442))
                begin
                  reg474 <= (reg470 || reg396);
                  for (forvar475 = (1'h0); (forvar475 < (2'h3)); forvar475 = (forvar475 + (1'h1)))
                    begin
                      reg476 <= (reg485[(1'h1):(1'h1)] && $unsigned(((reg423 ?
                          wire391 : reg432) || $signed(reg443))));
                      reg477 <= ((8'ha0) ?
                          $signed(forvar477[(4'h9):(3'h6)]) : ((((8'hb6) != (8'ha7)) * $unsigned(wire390)) ?
                              ($unsigned(reg404) ?
                                  wire390 : (reg483 ?
                                      reg437 : reg395)) : {$signed((8'hb9))}));
                      reg478 <= (8'ha6);
                      reg479 <= $unsigned($signed(((!forvar480) >>> forvar447)));
                    end
                end
              else
                begin
                  for (forvar474 = (1'h0); (forvar474 < (2'h3)); forvar474 = (forvar474 + (1'h1)))
                    begin
                      reg475 <= ({reg461} ?
                          ($unsigned(forvar447[(2'h3):(1'h0)]) && reg491) : ((^~$signed(wire390)) < $unsigned({(8'hb0)})));
                      reg476 <= $signed($signed($unsigned({wire389})));
                      reg477 <= $signed(($signed($signed(reg479)) ?
                          reg489 : (~|(~^(8'ha2)))));
                      reg478 <= (forvar448[(2'h3):(1'h1)] ?
                          forvar470 : (reg425 ?
                              (forvar475[(2'h3):(1'h0)] ?
                                  (reg476 ?
                                      forvar457 : reg485) : reg407[(1'h0):(1'h0)]) : {reg454}));
                    end
                end
            end
          for (forvar480 = (1'h0); (forvar480 < (2'h2)); forvar480 = (forvar480 + (1'h1)))
            begin
              reg481 <= ($unsigned({$signed(reg396)}) ?
                  ($unsigned(reg434) ?
                      forvar463[(4'h9):(3'h4)] : (~reg475)) : ({((8'hac) <= reg446)} ?
                      ($unsigned(reg446) < {reg493}) : $signed((~&reg431))));
              for (forvar482 = (1'h0); (forvar482 < (2'h2)); forvar482 = (forvar482 + (1'h1)))
                begin
                  for (forvar483 = (1'h0); (forvar483 < (1'h0)); forvar483 = (forvar483 + (1'h1)))
                    begin
                      reg484 <= reg416[(4'h8):(1'h0)];
                      reg485 <= (8'ha2);
                      reg486 <= $unsigned(((8'hb0) ?
                          $signed((reg410 ^ reg483)) : forvar449[(3'h6):(1'h1)]));
                      reg487 <= (&($signed(wire389[(3'h7):(3'h4)]) ?
                          $unsigned(((8'hba) || reg409)) : $unsigned(reg470)));
                    end
                  for (forvar488 = (1'h0); (forvar488 < (2'h2)); forvar488 = (forvar488 + (1'h1)))
                    begin
                      reg489 <= (~^(((reg427 != reg446) ?
                              forvar474 : $unsigned(forvar449)) ?
                          ((reg403 ?
                              (8'had) : forvar492) | reg467[(4'h9):(4'h8)]) : (|$signed(reg493))));
                      reg490 <= (!reg427[(3'h4):(1'h0)]);
                      reg491 <= reg431[(4'hf):(3'h7)];
                    end
                end
            end
          reg492 <= (reg394[(2'h2):(1'h0)] | forvar462);
          if ($signed($signed($unsigned($signed(reg407)))))
            begin
              for (forvar493 = (1'h0); (forvar493 < (1'h1)); forvar493 = (forvar493 + (1'h1)))
                begin
                  if (forvar447)
                    begin
                      reg494 <= $signed($unsigned((|{reg438})));
                      reg495 <= (!$signed($signed((reg453 ?
                          (8'ha6) : reg423))));
                      reg496 <= {(~|$unsigned((reg459 ? reg484 : (8'hb6))))};
                    end
                  else
                    begin
                      reg494 <= (((^~$signed(forvar469)) ^ ((reg470 ?
                              reg496 : reg427) < {(8'hb1)})) ?
                          ((8'ha7) || {forvar469[(3'h7):(3'h5)]}) : reg395);
                      reg495 <= {$signed(reg394[(1'h1):(1'h1)])};
                      reg496 <= reg466[(3'h5):(2'h3)];
                    end
                  for (forvar497 = (1'h0); (forvar497 < (1'h0)); forvar497 = (forvar497 + (1'h1)))
                    begin
                      reg498 <= (~&reg454);
                      reg499 <= {(~|((8'ha2) != $unsigned(reg451)))};
                    end
                  for (forvar500 = (1'h0); (forvar500 < (1'h1)); forvar500 = (forvar500 + (1'h1)))
                    begin
                      reg501 <= $unsigned(reg400);
                      reg502 <= forvar464;
                    end
                end
              for (forvar503 = (1'h0); (forvar503 < (1'h0)); forvar503 = (forvar503 + (1'h1)))
                begin
                  for (forvar504 = (1'h0); (forvar504 < (2'h3)); forvar504 = (forvar504 + (1'h1)))
                    begin
                      reg505 <= $signed(forvar463[(3'h4):(2'h2)]);
                      reg506 <= (!reg450[(3'h5):(1'h1)]);
                      reg507 <= (+$signed(((forvar477 ?
                          reg401 : reg395) & (reg485 < reg498))));
                      reg508 <= (wire386 ?
                          $signed((!$unsigned(forvar449))) : reg475);
                    end
                end
              for (forvar509 = (1'h0); (forvar509 < (2'h2)); forvar509 = (forvar509 + (1'h1)))
                begin
                  for (forvar510 = (1'h0); (forvar510 < (2'h3)); forvar510 = (forvar510 + (1'h1)))
                    begin
                      reg511 <= reg409;
                      reg512 <= $signed((((reg392 >= reg486) >= (reg476 | reg438)) < (^(reg428 ?
                          (8'hb4) : reg476))));
                      reg513 <= ($unsigned(reg464) ?
                          $unsigned($signed((8'ha2))) : (($unsigned(reg454) ?
                                  $signed(forvar469) : ((8'hac) ?
                                      reg425 : reg475)) ?
                              (((8'hba) ? reg396 : reg406) + (reg437 ?
                                  reg466 : reg476)) : (&$signed(forvar504))));
                    end
                  if ($signed(reg408[(1'h0):(1'h0)]))
                    begin
                      reg514 <= reg425[(3'h4):(3'h4)];
                      reg515 <= ((~(8'hab)) ?
                          (($signed(reg438) * (reg453 < (8'hb8))) ?
                              (8'had) : ($unsigned(forvar464) ?
                                  reg511[(3'h4):(3'h4)] : $signed(reg464))) : (reg475[(4'h8):(3'h6)] && {$unsigned(reg475)}));
                      reg516 <= reg394[(2'h3):(2'h3)];
                      reg517 <= (8'hb7);
                    end
                  else
                    begin
                      reg514 <= $unsigned(((reg437 ^ (8'ha2)) ?
                          (reg506 <= $signed(reg427)) : ((+(8'h9c)) ?
                              (|reg496) : reg453[(3'h5):(1'h1)])));
                      reg515 <= $signed((8'hb3));
                      reg516 <= forvar493[(4'h8):(3'h7)];
                    end
                  if ((^~reg465[(3'h5):(3'h5)]))
                    begin
                      reg518 <= ($unsigned(reg423[(3'h5):(1'h0)]) ?
                          reg427 : $unsigned((~^(forvar509 > (8'hb6)))));
                      reg519 <= (reg453 ?
                          (reg470[(3'h4):(1'h0)] != $signed({wire386})) : $signed(((reg450 ?
                              forvar477 : reg460) >>> reg471)));
                      reg520 <= reg476[(4'ha):(4'ha)];
                      reg521 <= (&reg437[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg518 <= ($signed(forvar469) < ({reg418[(2'h3):(2'h2)]} ?
                          ($signed(reg429) ?
                              $unsigned(reg433) : (+reg512)) : wire390));
                      reg519 <= $signed(reg498[(4'h9):(3'h4)]);
                    end
                end
              for (forvar522 = (1'h0); (forvar522 < (1'h1)); forvar522 = (forvar522 + (1'h1)))
                begin
                  reg523 <= (reg485 >> $unsigned($signed(reg517)));
                  for (forvar524 = (1'h0); (forvar524 < (1'h0)); forvar524 = (forvar524 + (1'h1)))
                    begin
                      reg525 <= reg475[(3'h5):(2'h2)];
                      reg526 <= (+$signed({reg421}));
                      reg527 <= {$signed((&((8'hb0) ? reg450 : reg434)))};
                      reg528 <= (+(~|($unsigned(reg465) >> (8'ha2))));
                    end
                  if ($unsigned($unsigned((~&$unsigned((8'ha2))))))
                    begin
                      reg529 <= (reg528[(3'h4):(2'h2)] > $signed((+(reg487 ^ reg426))));
                    end
                  else
                    begin
                      reg529 <= ($signed({{reg404}}) ?
                          reg402[(4'h9):(1'h0)] : reg443[(3'h4):(1'h1)]);
                      reg530 <= ($unsigned({(forvar483 ?
                              reg433 : reg453)}) - {reg470[(3'h7):(1'h0)]});
                      reg531 <= $unsigned((reg517[(1'h1):(1'h0)] >= $unsigned(reg490)));
                    end
                  if ($signed((reg415[(1'h1):(1'h1)] ^~ (~^reg395[(3'h4):(1'h0)]))))
                    begin
                      reg532 <= $unsigned((~(~^$unsigned(reg416))));
                    end
                  else
                    begin
                      reg532 <= ((reg467[(4'hc):(4'hb)] >>> {{reg490}}) & (reg475 == (8'h9e)));
                      reg533 <= (~|$unsigned((^~reg427)));
                    end
                end
            end
          else
            begin
              for (forvar493 = (1'h0); (forvar493 < (1'h0)); forvar493 = (forvar493 + (1'h1)))
                begin
                  if ($unsigned($signed(((reg484 != reg479) ?
                      wire386[(1'h0):(1'h0)] : $signed((8'hb6))))))
                    begin
                      reg494 <= {($unsigned((-(8'h9f))) ?
                              $unsigned(reg461) : $unsigned(forvar504[(1'h1):(1'h1)]))};
                    end
                  else
                    begin
                      reg494 <= {(~|{((8'ha7) ? reg432 : reg481)})};
                      reg495 <= reg425[(3'h4):(1'h1)];
                      reg496 <= (((~&(8'hb1)) ?
                          $unsigned($signed(reg494)) : reg416[(2'h2):(1'h1)]) > $signed(reg466));
                    end
                  for (forvar497 = (1'h0); (forvar497 < (1'h1)); forvar497 = (forvar497 + (1'h1)))
                    begin
                      reg498 <= reg512;
                    end
                  if (reg516)
                    begin
                      reg499 <= (~&((reg428 ? forvar503 : $signed(reg450)) ?
                          ((reg484 ^~ reg521) ?
                              (-forvar497) : (reg404 ?
                                  forvar465 : reg499)) : (^~(reg434 ?
                              reg511 : reg421))));
                    end
                  else
                    begin
                      reg499 <= ((reg513[(2'h2):(1'h1)] ?
                          $unsigned($signed(forvar447)) : reg402) >= $signed(reg495[(3'h4):(2'h3)]));
                      reg500 <= (forvar462 ?
                          reg420 : (&((reg520 > reg481) ^ $signed(forvar457))));
                      reg501 <= $signed($unsigned(((reg498 >>> reg476) || (reg464 << reg392))));
                    end
                end
              if ($unsigned($signed(reg434[(1'h1):(1'h0)])))
                begin
                  if (forvar448[(2'h2):(1'h0)])
                    begin
                      reg502 <= $signed(reg435[(4'h9):(1'h1)]);
                      reg503 <= reg475;
                      reg504 <= (reg469 & $signed(forvar449[(4'h8):(3'h5)]));
                      reg505 <= ((((~forvar492) ?
                              (reg463 == reg441) : reg396) != $signed({reg493})) ?
                          reg399 : $unsigned($signed($signed(reg488))));
                    end
                  else
                    begin
                      reg502 <= forvar474[(3'h4):(1'h0)];
                      reg503 <= {(-($unsigned(reg517) ?
                              (&forvar500) : (^~(8'h9f))))};
                      reg504 <= {reg442[(3'h7):(3'h5)]};
                    end
                end
              else
                begin
                  for (forvar502 = (1'h0); (forvar502 < (1'h0)); forvar502 = (forvar502 + (1'h1)))
                    begin
                      reg503 <= {reg514[(3'h7):(1'h0)]};
                      reg504 <= reg461[(2'h3):(1'h0)];
                      reg505 <= reg446[(3'h5):(3'h4)];
                      reg506 <= reg453[(3'h6):(2'h3)];
                    end
                  for (forvar507 = (1'h0); (forvar507 < (1'h1)); forvar507 = (forvar507 + (1'h1)))
                    begin
                      reg508 <= $signed($signed($signed((8'ha6))));
                      reg509 <= $unsigned(reg477[(3'h7):(3'h7)]);
                      reg510 <= $signed((8'hb7));
                      reg511 <= reg486;
                    end
                end
            end
        end
    end
  assign wire534 = ($signed((8'h9e)) ?
                       {(~|reg425[(3'h4):(1'h0)])} : $unsigned((reg461 != (!reg427))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1179
#(parameter param1530 = (((((8'haa) - (8'hba)) <<< ((8'hb9) && (8'h9c))) < ({(8'hb3)} <= {(8'hb2)})) ? ({((8'haa) ? (8'h9f) : (8'ha1))} ? ((8'hb9) ? ((8'hba) ? (8'hb6) : (8'ha1)) : ((8'haa) ? (8'hb7) : (8'h9d))) : ({(8'hb6)} != ((8'ha8) << (8'ha1)))) : (((~&(8'ha0)) ? ((8'ha6) ? (8'hac) : (8'had)) : ((8'haa) ? (8'ha3) : (8'ha6))) | (((8'hb1) ? (8'hae) : (8'hb3)) ? {(8'hab)} : ((8'h9f) ? (8'h9e) : (8'haa))))))
(y, clk, wire1183, wire1182, wire1181, wire1180);
  output wire [(32'h72b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire1183;
  input wire [(4'hc):(1'h0)] wire1182;
  input wire [(3'h7):(1'h0)] wire1181;
  input wire [(4'h8):(1'h0)] wire1180;
  wire signed [(4'h8):(1'h0)] wire1529;
  wire [(4'hb):(1'h0)] wire1528;
  wire signed [(4'ha):(1'h0)] wire1527;
  wire signed [(3'h6):(1'h0)] wire1526;
  wire [(4'hf):(1'h0)] wire1525;
  wire [(5'h10):(1'h0)] wire1472;
  wire signed [(4'hc):(1'h0)] wire1471;
  wire [(4'hc):(1'h0)] wire1375;
  wire [(5'h10):(1'h0)] wire1373;
  wire [(3'h4):(1'h0)] wire1186;
  wire signed [(4'hb):(1'h0)] wire1185;
  wire [(5'h10):(1'h0)] wire1184;
  reg [(4'h8):(1'h0)] reg1516 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1515 = (1'h0);
  reg [(4'hd):(1'h0)] reg1512 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1508 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1503 = (1'h0);
  reg [(4'ha):(1'h0)] reg1502 = (1'h0);
  reg [(4'ha):(1'h0)] reg1475 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1476 = (1'h0);
  reg [(5'h10):(1'h0)] reg1483 = (1'h0);
  reg [(2'h3):(1'h0)] reg1478 = (1'h0);
  reg [(3'h6):(1'h0)] reg1524 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1523 = (1'h0);
  reg [(4'hd):(1'h0)] reg1522 = (1'h0);
  reg [(4'ha):(1'h0)] reg1521 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1519 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1518 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1517 = (1'h0);
  reg [(5'h10):(1'h0)] reg1514 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1513 = (1'h0);
  reg [(3'h5):(1'h0)] reg1511 = (1'h0);
  reg [(4'he):(1'h0)] reg1509 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1507 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1506 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1505 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1504 = (1'h0);
  reg [(2'h2):(1'h0)] reg1500 = (1'h0);
  reg [(4'hb):(1'h0)] reg1499 = (1'h0);
  reg [(3'h7):(1'h0)] reg1498 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1497 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1495 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1494 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1493 = (1'h0);
  reg [(4'hf):(1'h0)] reg1492 = (1'h0);
  reg [(3'h4):(1'h0)] reg1490 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1489 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1488 = (1'h0);
  reg [(4'h8):(1'h0)] reg1487 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1486 = (1'h0);
  reg [(2'h3):(1'h0)] reg1485 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1484 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1482 = (1'h0);
  reg [(2'h3):(1'h0)] reg1481 = (1'h0);
  reg [(4'h8):(1'h0)] reg1480 = (1'h0);
  reg [(3'h4):(1'h0)] reg1479 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1477 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1474 = (1'h0);
  reg [(4'ha):(1'h0)] reg1473 = (1'h0);
  reg [(3'h7):(1'h0)] reg1470 = (1'h0);
  reg [(2'h3):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1468 = (1'h0);
  reg [(2'h2):(1'h0)] reg1467 = (1'h0);
  reg [(4'hd):(1'h0)] reg1466 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1463 = (1'h0);
  reg [(4'ha):(1'h0)] reg1464 = (1'h0);
  reg [(4'ha):(1'h0)] reg1461 = (1'h0);
  reg [(4'hb):(1'h0)] reg1460 = (1'h0);
  reg [(2'h3):(1'h0)] reg1458 = (1'h0);
  reg [(4'hb):(1'h0)] reg1457 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1456 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1455 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1453 = (1'h0);
  reg [(4'hb):(1'h0)] reg1454 = (1'h0);
  reg [(2'h3):(1'h0)] reg1452 = (1'h0);
  reg [(3'h6):(1'h0)] reg1450 = (1'h0);
  reg [(4'h8):(1'h0)] reg1449 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1447 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1446 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1441 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1436 = (1'h0);
  reg [(4'hf):(1'h0)] reg1445 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1444 = (1'h0);
  reg [(4'hc):(1'h0)] reg1443 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1442 = (1'h0);
  reg [(4'hf):(1'h0)] reg1440 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1439 = (1'h0);
  reg [(2'h2):(1'h0)] reg1438 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1437 = (1'h0);
  reg [(4'hd):(1'h0)] reg1434 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1430 = (1'h0);
  reg [(4'he):(1'h0)] reg1433 = (1'h0);
  reg [(4'hf):(1'h0)] reg1432 = (1'h0);
  reg [(5'h10):(1'h0)] reg1431 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1426 = (1'h0);
  reg [(2'h2):(1'h0)] reg1422 = (1'h0);
  reg [(5'h10):(1'h0)] reg1429 = (1'h0);
  reg [(4'ha):(1'h0)] reg1428 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1427 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1425 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1424 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1423 = (1'h0);
  reg [(4'h9):(1'h0)] reg1421 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1420 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1406 = (1'h0);
  reg [(3'h4):(1'h0)] reg1417 = (1'h0);
  reg [(5'h10):(1'h0)] reg1416 = (1'h0);
  reg [(4'hc):(1'h0)] reg1415 = (1'h0);
  reg [(3'h4):(1'h0)] reg1414 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1413 = (1'h0);
  reg [(4'hf):(1'h0)] reg1410 = (1'h0);
  reg [(5'h10):(1'h0)] reg1409 = (1'h0);
  reg [(4'ha):(1'h0)] reg1408 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1407 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1405 = (1'h0);
  reg [(4'he):(1'h0)] reg1404 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1403 = (1'h0);
  reg [(4'hf):(1'h0)] reg1402 = (1'h0);
  reg [(4'h9):(1'h0)] reg1386 = (1'h0);
  reg [(4'hb):(1'h0)] reg1378 = (1'h0);
  reg [(4'he):(1'h0)] reg1401 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1396 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1400 = (1'h0);
  reg [(4'hb):(1'h0)] reg1399 = (1'h0);
  reg [(4'hd):(1'h0)] reg1398 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1397 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1395 = (1'h0);
  reg [(4'hc):(1'h0)] reg1394 = (1'h0);
  reg [(4'he):(1'h0)] reg1393 = (1'h0);
  reg [(2'h2):(1'h0)] reg1392 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1391 = (1'h0);
  reg [(4'he):(1'h0)] reg1390 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1389 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1388 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1387 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1385 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1384 = (1'h0);
  reg [(3'h7):(1'h0)] reg1382 = (1'h0);
  reg [(5'h10):(1'h0)] reg1381 = (1'h0);
  reg [(4'hb):(1'h0)] reg1380 = (1'h0);
  reg [(4'he):(1'h0)] reg1379 = (1'h0);
  reg [(2'h3):(1'h0)] reg1376 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1514 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1506 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1500 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1488 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1487 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1484 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1481 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1520 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1516 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1515 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1512 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1510 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1508 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1503 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1502 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1501 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1496 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1491 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1483 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1478 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1476 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1475 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1465 = (1'h0);
  reg [(4'he):(1'h0)] forvar1461 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1463 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1462 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1459 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1453 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1451 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1448 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1439 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1437 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1441 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1436 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1435 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1430 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1423 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1426 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1422 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1419 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1418 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1412 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1411 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1402 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1406 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1390 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1389 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1385 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1379 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1399 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1391 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1396 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1386 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1383 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1378 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1377 = (1'h0);
  assign y = {wire1529,
                 wire1528,
                 wire1527,
                 wire1526,
                 wire1525,
                 wire1472,
                 wire1471,
                 wire1375,
                 wire1373,
                 wire1186,
                 wire1185,
                 wire1184,
                 reg1516,
                 reg1515,
                 reg1512,
                 reg1508,
                 reg1503,
                 reg1502,
                 reg1475,
                 reg1476,
                 reg1483,
                 reg1478,
                 reg1524,
                 reg1523,
                 reg1522,
                 reg1521,
                 reg1519,
                 reg1518,
                 reg1517,
                 reg1514,
                 reg1513,
                 reg1511,
                 reg1509,
                 reg1507,
                 reg1506,
                 reg1505,
                 reg1504,
                 reg1500,
                 reg1499,
                 reg1498,
                 reg1497,
                 reg1495,
                 reg1494,
                 reg1493,
                 reg1492,
                 reg1490,
                 reg1489,
                 reg1488,
                 reg1487,
                 reg1486,
                 reg1485,
                 reg1484,
                 reg1482,
                 reg1481,
                 reg1480,
                 reg1479,
                 reg1477,
                 reg1474,
                 reg1473,
                 reg1470,
                 reg1469,
                 reg1468,
                 reg1467,
                 reg1466,
                 reg1463,
                 reg1464,
                 reg1461,
                 reg1460,
                 reg1458,
                 reg1457,
                 reg1456,
                 reg1455,
                 reg1453,
                 reg1454,
                 reg1452,
                 reg1450,
                 reg1449,
                 reg1447,
                 reg1446,
                 reg1441,
                 reg1436,
                 reg1445,
                 reg1444,
                 reg1443,
                 reg1442,
                 reg1440,
                 reg1439,
                 reg1438,
                 reg1437,
                 reg1434,
                 reg1430,
                 reg1433,
                 reg1432,
                 reg1431,
                 reg1426,
                 reg1422,
                 reg1429,
                 reg1428,
                 reg1427,
                 reg1425,
                 reg1424,
                 reg1423,
                 reg1421,
                 reg1420,
                 reg1406,
                 reg1417,
                 reg1416,
                 reg1415,
                 reg1414,
                 reg1413,
                 reg1410,
                 reg1409,
                 reg1408,
                 reg1407,
                 reg1405,
                 reg1404,
                 reg1403,
                 reg1402,
                 reg1386,
                 reg1378,
                 reg1401,
                 reg1396,
                 reg1400,
                 reg1399,
                 reg1398,
                 reg1397,
                 reg1395,
                 reg1394,
                 reg1393,
                 reg1392,
                 reg1391,
                 reg1390,
                 reg1389,
                 reg1388,
                 reg1387,
                 reg1385,
                 reg1384,
                 reg1382,
                 reg1381,
                 reg1380,
                 reg1379,
                 reg1376,
                 forvar1514,
                 forvar1506,
                 forvar1500,
                 forvar1488,
                 forvar1487,
                 forvar1484,
                 forvar1481,
                 forvar1520,
                 forvar1516,
                 forvar1515,
                 forvar1512,
                 forvar1510,
                 forvar1508,
                 forvar1503,
                 forvar1502,
                 forvar1501,
                 forvar1496,
                 forvar1491,
                 forvar1483,
                 forvar1478,
                 forvar1476,
                 forvar1475,
                 forvar1465,
                 forvar1461,
                 forvar1463,
                 forvar1462,
                 forvar1459,
                 forvar1453,
                 forvar1451,
                 forvar1448,
                 forvar1439,
                 forvar1437,
                 forvar1441,
                 forvar1436,
                 forvar1435,
                 forvar1430,
                 forvar1423,
                 forvar1426,
                 forvar1422,
                 forvar1419,
                 forvar1418,
                 forvar1412,
                 forvar1411,
                 forvar1402,
                 forvar1406,
                 forvar1390,
                 forvar1389,
                 forvar1385,
                 forvar1379,
                 forvar1399,
                 forvar1391,
                 forvar1396,
                 forvar1386,
                 forvar1383,
                 forvar1378,
                 forvar1377,
                 (1'h0)};
  assign wire1184 = (~(!$unsigned({wire1180})));
  assign wire1185 = (&wire1184);
  assign wire1186 = ($unsigned($signed((|wire1182))) ?
                        wire1181[(3'h5):(1'h1)] : wire1183[(4'ha):(1'h1)]);
  module1187 #() modinst1374 (.wire1189(wire1184), .wire1190(wire1180), .wire1188(wire1185), .clk(clk), .y(wire1373), .wire1191(wire1183));
  assign wire1375 = $unsigned($signed($signed((8'hb3))));
  always
    @(posedge clk) begin
      reg1376 <= wire1186[(2'h2):(1'h0)];
      for (forvar1377 = (1'h0); (forvar1377 < (2'h3)); forvar1377 = (forvar1377 + (1'h1)))
        begin
          if ({($signed((~wire1375)) & {(wire1373 != wire1183)})})
            begin
              for (forvar1378 = (1'h0); (forvar1378 < (1'h1)); forvar1378 = (forvar1378 + (1'h1)))
                begin
                  if (($unsigned(wire1186[(1'h1):(1'h1)]) ?
                      wire1184[(4'he):(3'h5)] : $unsigned($signed((8'hb3)))))
                    begin
                      reg1379 <= $signed({$signed((forvar1377 ?
                              wire1186 : wire1186))});
                      reg1380 <= (reg1379[(2'h3):(2'h2)] ~^ (((forvar1377 ?
                              wire1182 : forvar1378) ^ wire1184) ?
                          wire1180 : (~|(8'hb1))));
                      reg1381 <= forvar1377;
                    end
                  else
                    begin
                      reg1379 <= ((reg1379 == $signed(wire1185[(4'h9):(2'h3)])) ^ (^{((8'ha4) | wire1180)}));
                      reg1380 <= $unsigned(({$unsigned(wire1375)} ?
                          ((wire1183 ?
                              reg1379 : forvar1378) >= wire1183[(4'h8):(4'h8)]) : (wire1373 ?
                              (|wire1181) : reg1380[(1'h0):(1'h0)])));
                      reg1381 <= $signed(((((8'hb1) * wire1184) == reg1379) ?
                          wire1375[(4'hc):(2'h2)] : (|(reg1376 ?
                              wire1181 : reg1381))));
                      reg1382 <= ($signed($signed((wire1186 <<< forvar1377))) && $signed($unsigned((reg1380 && wire1184))));
                    end
                  for (forvar1383 = (1'h0); (forvar1383 < (2'h3)); forvar1383 = (forvar1383 + (1'h1)))
                    begin
                      reg1384 <= $unsigned((~(!(forvar1383 ?
                          wire1186 : (8'haa)))));
                      reg1385 <= reg1384;
                    end
                  for (forvar1386 = (1'h0); (forvar1386 < (2'h2)); forvar1386 = (forvar1386 + (1'h1)))
                    begin
                      reg1387 <= $signed($unsigned(forvar1386));
                      reg1388 <= $unsigned(reg1382);
                      reg1389 <= reg1376[(1'h0):(1'h0)];
                    end
                end
              if ((!reg1381[(1'h1):(1'h1)]))
                begin
                  if ((reg1387[(1'h0):(1'h0)] ?
                      {$unsigned((^forvar1378))} : (8'h9f)))
                    begin
                      reg1390 <= $unsigned(reg1389);
                      reg1391 <= $unsigned(((((8'hba) - wire1185) ?
                              ((8'ha9) ?
                                  (8'hb8) : wire1375) : $signed(wire1180)) ?
                          ($unsigned(forvar1377) ^ $signed(forvar1383)) : $signed((wire1182 >> reg1387))));
                      reg1392 <= {wire1184[(3'h5):(1'h0)]};
                      reg1393 <= $unsigned(wire1184[(4'hb):(1'h1)]);
                    end
                  else
                    begin
                      reg1390 <= {($signed(reg1381[(1'h0):(1'h0)]) ?
                              reg1388[(4'ha):(3'h7)] : reg1382)};
                      reg1391 <= (wire1375 ?
                          (|((wire1185 >= wire1186) - (-reg1381))) : {(reg1381[(4'ha):(4'h9)] ?
                                  ((8'hac) ?
                                      reg1389 : (8'haa)) : $signed((8'hae)))});
                      reg1392 <= forvar1383[(2'h3):(1'h0)];
                    end
                  reg1394 <= $signed((((|reg1381) > (wire1373 ?
                      reg1387 : reg1390)) > $signed(reg1391[(1'h1):(1'h0)])));
                  reg1395 <= (8'hb2);
                  for (forvar1396 = (1'h0); (forvar1396 < (1'h1)); forvar1396 = (forvar1396 + (1'h1)))
                    begin
                      reg1397 <= {$signed(((reg1382 && reg1393) ?
                              reg1388[(3'h4):(1'h1)] : {reg1393}))};
                      reg1398 <= (8'ha8);
                      reg1399 <= $unsigned((8'hac));
                      reg1400 <= $unsigned((~^$signed((reg1390 ?
                          reg1379 : wire1180))));
                    end
                end
              else
                begin
                  reg1390 <= ($signed(reg1381) - $unsigned({{reg1376}}));
                  for (forvar1391 = (1'h0); (forvar1391 < (1'h0)); forvar1391 = (forvar1391 + (1'h1)))
                    begin
                      reg1392 <= wire1182;
                      reg1393 <= (((~|forvar1391[(2'h2):(1'h1)]) ?
                          $signed((reg1385 ~^ reg1390)) : $signed(reg1391)) * reg1400[(3'h5):(1'h1)]);
                      reg1394 <= (8'h9d);
                      reg1395 <= wire1182;
                    end
                  if (((forvar1386 ?
                          $signed((forvar1377 ? reg1388 : reg1392)) : (8'hb8)) ?
                      $unsigned(({(8'haa)} ?
                          (reg1385 << reg1393) : $signed(reg1389))) : reg1380[(4'ha):(2'h2)]))
                    begin
                      reg1396 <= reg1384[(4'ha):(2'h2)];
                      reg1397 <= {(((|forvar1383) + (wire1375 | (8'hab))) ~^ $unsigned(reg1395))};
                      reg1398 <= ($unsigned((+{reg1398})) ?
                          (((wire1185 ^ reg1388) || reg1399) ?
                              $unsigned(reg1384) : {$unsigned(wire1375)}) : (8'ha8));
                    end
                  else
                    begin
                      reg1396 <= (($signed(reg1379[(3'h5):(3'h5)]) ?
                          {$unsigned(reg1392)} : reg1381[(1'h0):(1'h0)]) * $signed({$signed(reg1400)}));
                      reg1397 <= $signed($signed($unsigned(reg1376[(2'h2):(1'h1)])));
                      reg1398 <= $unsigned((8'hb1));
                    end
                  for (forvar1399 = (1'h0); (forvar1399 < (1'h0)); forvar1399 = (forvar1399 + (1'h1)))
                    begin
                      reg1400 <= (!(~$unsigned(wire1182[(4'ha):(4'ha)])));
                      reg1401 <= $unsigned(((^~$unsigned(reg1380)) ?
                          (8'ha7) : ((^~forvar1386) ~^ $unsigned((8'ha7)))));
                    end
                end
            end
          else
            begin
              if (($signed((reg1382[(2'h3):(2'h2)] ?
                      $unsigned(forvar1377) : $signed(reg1395))) ?
                  $unsigned(((wire1186 ^~ reg1387) ?
                      (reg1385 ?
                          forvar1383 : (8'ha8)) : (8'ha6))) : reg1397[(2'h2):(1'h0)]))
                begin
                  reg1378 <= reg1380;
                  for (forvar1379 = (1'h0); (forvar1379 < (1'h1)); forvar1379 = (forvar1379 + (1'h1)))
                    begin
                      reg1380 <= ({(~^(-reg1385))} <= $unsigned($signed(((8'hba) >> (8'hb9)))));
                    end
                  if (((((8'ha7) || $signed(forvar1396)) ?
                          (~|reg1387[(3'h4):(3'h4)]) : {$signed(reg1379)}) ?
                      $signed((+(reg1399 ?
                          forvar1383 : forvar1386))) : (-{$signed(reg1389)})))
                    begin
                      reg1381 <= forvar1396;
                    end
                  else
                    begin
                      reg1381 <= $unsigned((+(8'haa)));
                    end
                  reg1382 <= (^(((forvar1379 ?
                          forvar1396 : forvar1386) ^~ (wire1181 || wire1180)) ?
                      (~&forvar1377[(2'h3):(1'h1)]) : (reg1384[(2'h2):(1'h1)] | $signed(reg1394))));
                end
              else
                begin
                  for (forvar1378 = (1'h0); (forvar1378 < (1'h0)); forvar1378 = (forvar1378 + (1'h1)))
                    begin
                      reg1379 <= $unsigned(({(forvar1391 == reg1400)} - $unsigned($signed(reg1401))));
                      reg1380 <= reg1376[(2'h3):(1'h0)];
                      reg1381 <= reg1389[(2'h3):(2'h3)];
                      reg1382 <= $unsigned((!$unsigned((reg1395 ?
                          reg1381 : reg1399))));
                    end
                  for (forvar1383 = (1'h0); (forvar1383 < (2'h3)); forvar1383 = (forvar1383 + (1'h1)))
                    begin
                      reg1384 <= reg1388;
                    end
                  for (forvar1385 = (1'h0); (forvar1385 < (1'h0)); forvar1385 = (forvar1385 + (1'h1)))
                    begin
                      reg1386 <= $unsigned(((~^$signed(forvar1396)) ?
                          $signed((8'ha7)) : (|(forvar1378 << reg1395))));
                      reg1387 <= reg1397;
                      reg1388 <= $unsigned(($unsigned((^(8'ha0))) ?
                          $unsigned((+reg1398)) : (|wire1183)));
                    end
                end
              for (forvar1389 = (1'h0); (forvar1389 < (2'h3)); forvar1389 = (forvar1389 + (1'h1)))
                begin
                  for (forvar1390 = (1'h0); (forvar1390 < (2'h2)); forvar1390 = (forvar1390 + (1'h1)))
                    begin
                      reg1391 <= $signed((~((^~reg1397) >= reg1393[(4'h9):(3'h6)])));
                      reg1392 <= $unsigned($signed({((8'hab) ^~ forvar1379)}));
                    end
                  if ((&wire1181[(1'h0):(1'h0)]))
                    begin
                      reg1393 <= {$unsigned(((reg1387 || forvar1379) ^ (reg1376 >>> wire1181)))};
                      reg1394 <= (+$signed((&((8'ha0) ?
                          forvar1391 : reg1393))));
                    end
                  else
                    begin
                      reg1393 <= wire1185;
                      reg1394 <= $unsigned(wire1186);
                      reg1395 <= $signed(((^~$unsigned(reg1376)) ^~ reg1399));
                    end
                end
            end
          if ((reg1379[(4'hc):(4'h9)] + $unsigned(($signed(forvar1396) ?
              reg1386[(4'h9):(3'h7)] : (-forvar1391)))))
            begin
              if ({reg1388[(3'h7):(1'h0)]})
                begin
                  if (wire1182)
                    begin
                      reg1402 <= {reg1386[(2'h2):(2'h2)]};
                    end
                  else
                    begin
                      reg1402 <= $signed((reg1396 ?
                          {$signed(reg1390)} : {$signed(wire1180)}));
                      reg1403 <= $unsigned($unsigned(((8'had) ?
                          (forvar1385 ~^ reg1393) : (^reg1381))));
                      reg1404 <= ((forvar1391 && (^reg1384[(2'h3):(1'h1)])) ?
                          (^({reg1380} >> {reg1400})) : ($unsigned($unsigned(reg1382)) ?
                              reg1386 : $unsigned($unsigned(reg1389))));
                      reg1405 <= $unsigned(wire1185);
                    end
                  for (forvar1406 = (1'h0); (forvar1406 < (1'h1)); forvar1406 = (forvar1406 + (1'h1)))
                    begin
                      reg1407 <= $unsigned({reg1381[(5'h10):(4'hc)]});
                    end
                  if ($unsigned($signed(reg1399)))
                    begin
                      reg1408 <= reg1396[(3'h7):(1'h0)];
                      reg1409 <= $unsigned(forvar1383);
                    end
                  else
                    begin
                      reg1408 <= (-wire1185[(3'h4):(2'h3)]);
                      reg1409 <= (+(wire1184[(4'he):(4'hd)] ?
                          ($unsigned(forvar1396) ?
                              (^~reg1397) : reg1376[(2'h3):(1'h0)]) : $signed({forvar1377})));
                      reg1410 <= (~&$unsigned(reg1389[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar1402 = (1'h0); (forvar1402 < (1'h0)); forvar1402 = (forvar1402 + (1'h1)))
                    begin
                      reg1403 <= reg1401[(3'h4):(2'h2)];
                      reg1404 <= $signed({{reg1391[(4'h8):(3'h5)]}});
                      reg1405 <= reg1402;
                    end
                end
              for (forvar1411 = (1'h0); (forvar1411 < (2'h2)); forvar1411 = (forvar1411 + (1'h1)))
                begin
                  for (forvar1412 = (1'h0); (forvar1412 < (2'h3)); forvar1412 = (forvar1412 + (1'h1)))
                    begin
                      reg1413 <= reg1390[(4'h9):(3'h6)];
                    end
                  if (reg1389[(2'h3):(1'h1)])
                    begin
                      reg1414 <= reg1376;
                      reg1415 <= ({forvar1411} ?
                          $unsigned(forvar1390[(2'h2):(1'h1)]) : $signed((|reg1379)));
                    end
                  else
                    begin
                      reg1414 <= (~&(&forvar1379));
                      reg1415 <= wire1183[(3'h5):(2'h3)];
                      reg1416 <= $signed((wire1185[(3'h4):(1'h1)] ?
                          ((^~(8'hba)) - {forvar1399}) : (reg1413[(2'h3):(1'h0)] - (|(8'hba)))));
                    end
                  reg1417 <= ((^$unsigned(forvar1385)) ?
                      (~^$unsigned(forvar1390[(2'h3):(1'h1)])) : (~&(|(|reg1390))));
                end
            end
          else
            begin
              for (forvar1402 = (1'h0); (forvar1402 < (1'h0)); forvar1402 = (forvar1402 + (1'h1)))
                begin
                  if ((!($unsigned((reg1393 ^~ (8'hb1))) >= (^~forvar1383[(1'h0):(1'h0)]))))
                    begin
                      reg1403 <= (({{forvar1377}} ?
                              $unsigned((forvar1402 ?
                                  wire1183 : reg1403)) : $signed(((8'ha6) ?
                                  reg1386 : reg1398))) ?
                          (~|($unsigned(forvar1379) ?
                              ((8'hb4) <= reg1381) : (~^reg1380))) : $unsigned(reg1399));
                      reg1404 <= forvar1386;
                    end
                  else
                    begin
                      reg1403 <= ((($signed(reg1416) ^ (8'ha9)) ?
                              (((8'hae) ?
                                  wire1183 : reg1391) - forvar1383) : reg1394[(4'h8):(2'h3)]) ?
                          $signed((&(reg1413 ?
                              reg1376 : reg1401))) : forvar1377[(2'h2):(1'h1)]);
                      reg1404 <= reg1402[(4'ha):(3'h4)];
                      reg1405 <= $unsigned(reg1376[(1'h0):(1'h0)]);
                      reg1406 <= (reg1380[(4'h9):(3'h4)] || (!$unsigned(forvar1412)));
                    end
                end
            end
          if (reg1384)
            begin
              for (forvar1418 = (1'h0); (forvar1418 < (1'h1)); forvar1418 = (forvar1418 + (1'h1)))
                begin
                  for (forvar1419 = (1'h0); (forvar1419 < (2'h2)); forvar1419 = (forvar1419 + (1'h1)))
                    begin
                      reg1420 <= ((($unsigned(reg1404) ?
                          reg1379[(3'h6):(3'h6)] : (forvar1379 & reg1388)) == $unsigned(reg1390)) >> wire1375);
                      reg1421 <= {$unsigned($signed(reg1388[(4'hb):(1'h1)]))};
                    end
                  for (forvar1422 = (1'h0); (forvar1422 < (2'h3)); forvar1422 = (forvar1422 + (1'h1)))
                    begin
                      reg1423 <= reg1379[(3'h6):(1'h0)];
                      reg1424 <= ($signed((~^reg1389)) ^~ (-(forvar1377 ^~ reg1407)));
                      reg1425 <= ($unsigned($unsigned(reg1417[(2'h3):(1'h0)])) ?
                          (reg1380 || reg1414[(2'h2):(1'h1)]) : ($signed(reg1410[(4'h9):(4'h9)]) & (-$signed(reg1386))));
                    end
                  for (forvar1426 = (1'h0); (forvar1426 < (1'h1)); forvar1426 = (forvar1426 + (1'h1)))
                    begin
                      reg1427 <= {(+forvar1418)};
                      reg1428 <= (+(forvar1391[(3'h7):(3'h7)] ?
                          reg1391[(1'h0):(1'h0)] : $signed($unsigned(forvar1389))));
                      reg1429 <= $signed($signed($unsigned($signed(reg1415))));
                    end
                end
            end
          else
            begin
              for (forvar1418 = (1'h0); (forvar1418 < (1'h1)); forvar1418 = (forvar1418 + (1'h1)))
                begin
                  for (forvar1419 = (1'h0); (forvar1419 < (2'h3)); forvar1419 = (forvar1419 + (1'h1)))
                    begin
                      reg1420 <= (-(8'ha3));
                      reg1421 <= {(($signed(reg1409) ?
                              {reg1423} : reg1395[(4'hf):(4'hf)]) - $signed(forvar1385))};
                      reg1422 <= wire1184;
                    end
                end
              if (((~$unsigned({forvar1378})) ? {reg1404} : $signed((8'hb9))))
                begin
                  for (forvar1423 = (1'h0); (forvar1423 < (2'h3)); forvar1423 = (forvar1423 + (1'h1)))
                    begin
                      reg1424 <= wire1184;
                      reg1425 <= forvar1378;
                    end
                end
              else
                begin
                  for (forvar1423 = (1'h0); (forvar1423 < (1'h1)); forvar1423 = (forvar1423 + (1'h1)))
                    begin
                      reg1424 <= (wire1184 ?
                          (+$unsigned((reg1381 <= wire1373))) : {$signed($unsigned(reg1388))});
                      reg1425 <= wire1185;
                      reg1426 <= (~&wire1185[(4'ha):(3'h6)]);
                    end
                  if (($unsigned($unsigned(forvar1386)) ?
                      ((!(reg1382 ? forvar1422 : forvar1412)) ?
                          $unsigned({reg1425}) : ((forvar1386 ?
                              reg1380 : reg1381) ^~ (reg1407 != wire1180))) : $unsigned($signed($unsigned((8'hab))))))
                    begin
                      reg1427 <= ($signed((+forvar1418[(1'h1):(1'h0)])) >= (reg1381 ?
                          $signed((8'h9d)) : $unsigned(reg1427)));
                      reg1428 <= {$unsigned({$unsigned(wire1373)})};
                      reg1429 <= $unsigned(((|$signed(reg1392)) + $unsigned((^reg1403))));
                    end
                  else
                    begin
                      reg1427 <= (~|$signed({reg1382[(3'h7):(3'h4)]}));
                    end
                end
              if (reg1382)
                begin
                  for (forvar1430 = (1'h0); (forvar1430 < (1'h1)); forvar1430 = (forvar1430 + (1'h1)))
                    begin
                      reg1431 <= (((((8'hae) & forvar1430) ?
                              $unsigned((8'hb9)) : (~&forvar1430)) & (~|(forvar1386 ?
                              reg1423 : reg1398))) ?
                          ((8'ha6) ?
                              ($unsigned(forvar1399) ?
                                  (forvar1383 ?
                                      reg1381 : reg1401) : reg1379) : (~&{(8'hb9)})) : (forvar1377[(1'h0):(1'h0)] & {reg1395[(3'h6):(1'h1)]}));
                      reg1432 <= ({($unsigned(reg1392) <= $signed(reg1413))} ?
                          (wire1185 ?
                              $unsigned(reg1380) : reg1409) : $unsigned((|(~|(8'ha0)))));
                      reg1433 <= $signed($unsigned(($signed((8'ha3)) ?
                          (!reg1404) : ((8'ha9) | forvar1385))));
                    end
                end
              else
                begin
                  if (reg1399[(1'h0):(1'h0)])
                    begin
                      reg1430 <= (reg1379 | (~reg1423[(4'he):(2'h3)]));
                      reg1431 <= $unsigned($signed(wire1375[(3'h7):(1'h0)]));
                    end
                  else
                    begin
                      reg1430 <= wire1180[(3'h6):(3'h6)];
                    end
                end
              reg1434 <= (~&(reg1376 < ($unsigned(forvar1391) ^~ (&reg1392))));
            end
          if ({$unsigned((reg1422[(1'h1):(1'h1)] <<< (reg1381 ?
                  forvar1386 : reg1400)))})
            begin
              for (forvar1435 = (1'h0); (forvar1435 < (1'h0)); forvar1435 = (forvar1435 + (1'h1)))
                begin
                  for (forvar1436 = (1'h0); (forvar1436 < (2'h3)); forvar1436 = (forvar1436 + (1'h1)))
                    begin
                      reg1437 <= ((wire1183[(4'ha):(3'h6)] <= ((reg1397 > reg1420) ^ $signed(reg1387))) * $unsigned($signed($signed(reg1380))));
                      reg1438 <= $unsigned(reg1395[(4'hb):(3'h7)]);
                      reg1439 <= reg1380[(3'h4):(2'h2)];
                      reg1440 <= {{$unsigned($signed(reg1427))}};
                    end
                  for (forvar1441 = (1'h0); (forvar1441 < (1'h0)); forvar1441 = (forvar1441 + (1'h1)))
                    begin
                      reg1442 <= (^~(|($signed(reg1398) ?
                          $unsigned((8'h9d)) : $unsigned(forvar1402))));
                      reg1443 <= $signed($signed((reg1397 >> reg1430[(2'h3):(1'h0)])));
                      reg1444 <= reg1404[(4'ha):(3'h6)];
                    end
                end
              reg1445 <= (reg1394[(3'h5):(1'h1)] <= wire1184[(3'h5):(2'h3)]);
            end
          else
            begin
              if ($unsigned((({reg1386} >> $signed((8'ha3))) ?
                  reg1376 : (~((8'hb3) ? reg1443 : (8'hb9))))))
                begin
                  for (forvar1435 = (1'h0); (forvar1435 < (2'h2)); forvar1435 = (forvar1435 + (1'h1)))
                    begin
                      reg1436 <= {reg1429};
                      reg1437 <= $unsigned((((reg1405 <= reg1401) || $unsigned(forvar1379)) ?
                          ($signed(reg1387) << (forvar1441 ?
                              (8'hab) : forvar1422)) : (~$unsigned((8'hb0)))));
                      reg1438 <= forvar1379;
                    end
                end
              else
                begin
                  for (forvar1435 = (1'h0); (forvar1435 < (1'h1)); forvar1435 = (forvar1435 + (1'h1)))
                    begin
                      reg1436 <= wire1186[(1'h0):(1'h0)];
                    end
                  for (forvar1437 = (1'h0); (forvar1437 < (1'h1)); forvar1437 = (forvar1437 + (1'h1)))
                    begin
                      reg1438 <= wire1181;
                    end
                end
              if ((~^(reg1425[(4'h8):(3'h7)] >>> (8'hb0))))
                begin
                  for (forvar1439 = (1'h0); (forvar1439 < (2'h2)); forvar1439 = (forvar1439 + (1'h1)))
                    begin
                      reg1440 <= {{(forvar1378[(1'h1):(1'h1)] ?
                                  $unsigned(reg1445) : $unsigned(forvar1390))}};
                      reg1441 <= $unsigned($signed(($unsigned(reg1393) ?
                          reg1378[(4'h8):(2'h2)] : forvar1422[(3'h4):(1'h0)])));
                      reg1442 <= $unsigned((|reg1389));
                      reg1443 <= (~^$unsigned($signed({reg1386})));
                    end
                end
              else
                begin
                  for (forvar1439 = (1'h0); (forvar1439 < (1'h1)); forvar1439 = (forvar1439 + (1'h1)))
                    begin
                      reg1440 <= reg1416;
                      reg1441 <= $unsigned((~{$signed(reg1401)}));
                      reg1442 <= forvar1422[(4'h8):(2'h3)];
                      reg1443 <= (((8'had) ?
                          ($unsigned((8'haa)) >>> $unsigned(reg1394)) : ((~reg1379) ?
                              $signed(reg1397) : $unsigned(reg1405))) | ($signed((wire1373 ?
                          (8'hb7) : forvar1391)) + $unsigned((reg1399 ?
                          forvar1402 : reg1405))));
                    end
                  if (($signed(({forvar1419} & reg1436[(2'h2):(2'h2)])) ?
                      ($unsigned((^reg1382)) && reg1405[(3'h7):(1'h0)]) : ({$unsigned(wire1183)} << reg1391[(3'h4):(2'h3)])))
                    begin
                      reg1444 <= $signed($unsigned(($signed(forvar1396) - (~wire1373))));
                      reg1445 <= $signed(((^~forvar1389[(2'h2):(1'h1)]) ?
                          {(reg1413 ^ forvar1437)} : ($signed(forvar1418) ~^ reg1399)));
                      reg1446 <= $unsigned((&(reg1391[(3'h5):(2'h2)] ?
                          $signed((8'ha8)) : wire1375)));
                      reg1447 <= (!reg1387[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg1444 <= $unsigned((!$signed((|reg1440))));
                    end
                  for (forvar1448 = (1'h0); (forvar1448 < (1'h1)); forvar1448 = (forvar1448 + (1'h1)))
                    begin
                      reg1449 <= ((^(^~(wire1183 < reg1437))) ?
                          $signed(forvar1412[(4'h8):(3'h6)]) : $unsigned($unsigned((forvar1391 ?
                              reg1402 : forvar1406))));
                      reg1450 <= forvar1411[(4'ha):(1'h0)];
                    end
                end
              if ({reg1434[(4'hb):(1'h0)]})
                begin
                  for (forvar1451 = (1'h0); (forvar1451 < (2'h2)); forvar1451 = (forvar1451 + (1'h1)))
                    begin
                      reg1452 <= forvar1406[(2'h3):(1'h0)];
                    end
                  for (forvar1453 = (1'h0); (forvar1453 < (1'h0)); forvar1453 = (forvar1453 + (1'h1)))
                    begin
                      reg1454 <= ({((8'haf) + (forvar1453 ?
                              reg1384 : forvar1412))} != ((|(&reg1396)) ?
                          ($unsigned((8'hb2)) ?
                              forvar1418[(1'h0):(1'h0)] : (wire1182 ?
                                  reg1401 : forvar1396)) : {$signed(forvar1378)}));
                    end
                end
              else
                begin
                  for (forvar1451 = (1'h0); (forvar1451 < (1'h1)); forvar1451 = (forvar1451 + (1'h1)))
                    begin
                      reg1452 <= $unsigned($signed($signed((&(8'h9f)))));
                      reg1453 <= reg1425;
                    end
                  if ((((forvar1439 ?
                          (wire1182 ?
                              reg1437 : reg1447) : (&reg1449)) >>> $signed($unsigned(reg1415))) ?
                      ((&(reg1437 ?
                          forvar1436 : reg1427)) <= $signed($signed(reg1409))) : ({reg1442[(3'h6):(1'h1)]} == (!(forvar1437 ?
                          (8'haf) : forvar1391)))))
                    begin
                      reg1454 <= $unsigned($signed((~$unsigned(reg1447))));
                    end
                  else
                    begin
                      reg1454 <= {reg1404};
                      reg1455 <= (~(~|((reg1384 <<< (8'hb4)) ~^ $signed(forvar1441))));
                    end
                  if ((reg1413 ?
                      $unsigned(((reg1382 * reg1387) <<< (8'hb4))) : ((&$unsigned(reg1402)) ^~ $signed((reg1417 ?
                          (8'ha0) : reg1450)))))
                    begin
                      reg1456 <= {(($signed((8'hae)) ?
                              (-reg1425) : $signed(forvar1389)) | ((-forvar1411) ?
                              {reg1441} : $unsigned(reg1426)))};
                      reg1457 <= reg1437;
                    end
                  else
                    begin
                      reg1456 <= $unsigned((|$signed($unsigned(reg1453))));
                      reg1457 <= reg1427[(4'h8):(3'h5)];
                      reg1458 <= {($unsigned((reg1414 ? reg1395 : reg1446)) ?
                              $unsigned(((8'haa) ?
                                  (8'h9c) : reg1394)) : forvar1436)};
                    end
                  for (forvar1459 = (1'h0); (forvar1459 < (1'h1)); forvar1459 = (forvar1459 + (1'h1)))
                    begin
                      reg1460 <= forvar1406[(2'h3):(1'h0)];
                    end
                end
            end
        end
      if (reg1416)
        begin
          reg1461 <= (^reg1434);
        end
      else
        begin
          if ($signed(($unsigned((~forvar1399)) > reg1382[(3'h5):(2'h2)])))
            begin
              reg1461 <= (8'hb4);
              for (forvar1462 = (1'h0); (forvar1462 < (1'h1)); forvar1462 = (forvar1462 + (1'h1)))
                begin
                  for (forvar1463 = (1'h0); (forvar1463 < (2'h2)); forvar1463 = (forvar1463 + (1'h1)))
                    begin
                      reg1464 <= $signed(({reg1397} ?
                          $signed(forvar1406) : ({reg1450} ?
                              (reg1409 * reg1414) : $signed(wire1185))));
                    end
                end
            end
          else
            begin
              for (forvar1461 = (1'h0); (forvar1461 < (1'h0)); forvar1461 = (forvar1461 + (1'h1)))
                begin
                  for (forvar1462 = (1'h0); (forvar1462 < (2'h3)); forvar1462 = (forvar1462 + (1'h1)))
                    begin
                      reg1463 <= $unsigned($unsigned(((8'ha7) ?
                          reg1402 : $unsigned(reg1382))));
                      reg1464 <= {(((reg1396 + wire1375) && (forvar1422 & (8'hb4))) ^ ($unsigned((8'ha2)) != ((8'hb4) ?
                              (8'ha0) : reg1390)))};
                    end
                  for (forvar1465 = (1'h0); (forvar1465 < (1'h1)); forvar1465 = (forvar1465 + (1'h1)))
                    begin
                      reg1466 <= ({reg1434} >> reg1438[(2'h2):(2'h2)]);
                      reg1467 <= ((8'hb8) ?
                          $unsigned(forvar1418[(2'h2):(2'h2)]) : (^((reg1432 ?
                              reg1466 : reg1439) <= (wire1180 ?
                              reg1447 : reg1422))));
                      reg1468 <= ($unsigned(forvar1451[(4'hd):(4'hc)]) | ({(~reg1401)} != $signed(forvar1379)));
                      reg1469 <= {(reg1385[(4'hb):(3'h7)] ?
                              (~&forvar1377) : ((|reg1468) ?
                                  {reg1444} : (|forvar1462)))};
                    end
                  reg1470 <= ({$signed(((8'hb2) > reg1378))} == (reg1404 ?
                      {forvar1423[(3'h7):(1'h0)]} : $unsigned($unsigned(forvar1448))));
                end
            end
        end
    end
  assign wire1471 = ($signed({$signed(wire1375)}) ?
                        (^~reg1409[(4'hb):(2'h2)]) : reg1389[(1'h0):(1'h0)]);
  assign wire1472 = $signed($signed(reg1401[(4'he):(2'h3)]));
  always
    @(posedge clk) begin
      reg1473 <= (reg1456[(3'h5):(2'h2)] | (reg1389 != (wire1471[(2'h3):(1'h0)] ?
          (wire1180 >= reg1434) : reg1416[(4'h9):(3'h6)])));
    end
  always
    @(posedge clk) begin
      reg1474 <= (~^$signed(({reg1423} ?
          $signed(reg1428) : $unsigned(wire1373))));
    end
  always
    @(posedge clk) begin
      if (({reg1396[(3'h6):(1'h0)]} >>> wire1471[(3'h6):(2'h2)]))
        begin
          for (forvar1475 = (1'h0); (forvar1475 < (1'h1)); forvar1475 = (forvar1475 + (1'h1)))
            begin
              for (forvar1476 = (1'h0); (forvar1476 < (2'h2)); forvar1476 = (forvar1476 + (1'h1)))
                begin
                  reg1477 <= $signed(({$unsigned(reg1467)} <= {(reg1430 << reg1450)}));
                  for (forvar1478 = (1'h0); (forvar1478 < (2'h3)); forvar1478 = (forvar1478 + (1'h1)))
                    begin
                      reg1479 <= wire1181;
                      reg1480 <= (reg1461 + (reg1431 ^~ (reg1402[(4'hf):(2'h2)] ?
                          (reg1400 < reg1386) : (reg1461 - reg1441))));
                      reg1481 <= (($signed(reg1477[(1'h0):(1'h0)]) - reg1437) & reg1430[(2'h2):(1'h1)]);
                      reg1482 <= ((reg1431 < (~|(reg1395 <<< reg1381))) ?
                          reg1407[(1'h1):(1'h1)] : $unsigned(($unsigned((8'hb0)) ?
                              ((8'hb8) - (8'hb2)) : reg1447)));
                    end
                end
              if ((($signed(reg1413) ~^ (reg1438[(1'h0):(1'h0)] ?
                  $unsigned(reg1455) : reg1378[(4'hb):(4'h9)])) | wire1375[(1'h0):(1'h0)]))
                begin
                  for (forvar1483 = (1'h0); (forvar1483 < (2'h2)); forvar1483 = (forvar1483 + (1'h1)))
                    begin
                      reg1484 <= $signed({(^$signed(reg1454))});
                      reg1485 <= ((reg1436[(1'h1):(1'h1)] ?
                          {reg1416} : (forvar1483 <= (reg1390 ?
                              reg1382 : reg1457))) || $signed((reg1380 > (^reg1402))));
                    end
                  reg1486 <= reg1481;
                  if (reg1391)
                    begin
                      reg1487 <= reg1404;
                    end
                  else
                    begin
                      reg1487 <= ((reg1469 ?
                              (~(wire1183 ?
                                  reg1479 : wire1373)) : ((reg1434 <= reg1413) ?
                                  (reg1446 ? (8'ha5) : reg1402) : (reg1401 ?
                                      reg1402 : wire1186))) ?
                          (forvar1476 ?
                              ((reg1477 ? reg1385 : reg1397) ?
                                  {reg1454} : reg1463) : ((reg1487 << reg1425) ?
                                  reg1404 : {reg1444})) : ($signed(((8'hb3) ?
                                  reg1425 : reg1482)) ?
                              $signed(reg1422) : $signed($unsigned(wire1183))));
                      reg1488 <= ((reg1470[(2'h2):(1'h0)] ^~ (reg1428[(2'h2):(2'h2)] - reg1405)) ?
                          (((8'hb4) <<< (reg1452 & reg1400)) ?
                              $unsigned($unsigned(reg1430)) : reg1414) : (^~$signed((reg1397 ?
                              reg1415 : (8'hb9)))));
                      reg1489 <= (reg1397[(4'hd):(3'h5)] >> reg1380);
                    end
                end
              else
                begin
                  for (forvar1483 = (1'h0); (forvar1483 < (1'h0)); forvar1483 = (forvar1483 + (1'h1)))
                    begin
                      reg1484 <= (8'hb1);
                      reg1485 <= $unsigned(reg1423);
                      reg1486 <= $unsigned({(^~(&wire1373))});
                    end
                  reg1487 <= reg1402[(3'h5):(1'h0)];
                end
              reg1490 <= forvar1483[(3'h5):(1'h1)];
              for (forvar1491 = (1'h0); (forvar1491 < (1'h0)); forvar1491 = (forvar1491 + (1'h1)))
                begin
                  if (reg1431[(4'hd):(2'h3)])
                    begin
                      reg1492 <= (((8'h9f) && reg1389) ?
                          wire1471[(3'h7):(2'h2)] : (~|reg1433));
                      reg1493 <= $signed(reg1442);
                      reg1494 <= ($unsigned((!$unsigned(reg1427))) && (((wire1181 ?
                              reg1477 : reg1426) - wire1184[(2'h2):(2'h2)]) ?
                          (((8'ha4) ? (8'hb4) : reg1454) >> (wire1375 ?
                              (8'ha9) : reg1397)) : ((~&reg1439) ?
                              ((8'h9d) ?
                                  forvar1476 : wire1375) : reg1427[(3'h7):(3'h6)])));
                    end
                  else
                    begin
                      reg1492 <= reg1463;
                    end
                  reg1495 <= $unsigned((reg1409 ?
                      $signed(reg1438) : ((reg1452 || reg1386) ?
                          (reg1421 ? reg1391 : reg1494) : (&(8'hab)))));
                  for (forvar1496 = (1'h0); (forvar1496 < (1'h1)); forvar1496 = (forvar1496 + (1'h1)))
                    begin
                      reg1497 <= $unsigned(reg1423);
                      reg1498 <= $unsigned(reg1430[(2'h2):(1'h1)]);
                      reg1499 <= {reg1461};
                      reg1500 <= $signed(reg1438[(1'h0):(1'h0)]);
                    end
                end
            end
          for (forvar1501 = (1'h0); (forvar1501 < (2'h3)); forvar1501 = (forvar1501 + (1'h1)))
            begin
              for (forvar1502 = (1'h0); (forvar1502 < (1'h1)); forvar1502 = (forvar1502 + (1'h1)))
                begin
                  for (forvar1503 = (1'h0); (forvar1503 < (2'h2)); forvar1503 = (forvar1503 + (1'h1)))
                    begin
                      reg1504 <= reg1439;
                    end
                  if (reg1480)
                    begin
                      reg1505 <= (!{$signed($signed((8'hb7)))});
                      reg1506 <= $signed((|((-reg1455) ?
                          $unsigned(reg1497) : (~^reg1395))));
                      reg1507 <= $signed(((reg1422[(1'h0):(1'h0)] ?
                              (wire1373 & reg1438) : $unsigned(reg1438)) ?
                          $unsigned($unsigned((8'hba))) : $unsigned($unsigned(reg1427))));
                    end
                  else
                    begin
                      reg1505 <= (~&$unsigned({{reg1461}}));
                      reg1506 <= $signed($signed(reg1477));
                    end
                  for (forvar1508 = (1'h0); (forvar1508 < (1'h1)); forvar1508 = (forvar1508 + (1'h1)))
                    begin
                      reg1509 <= ($signed({reg1420}) ?
                          reg1438[(1'h1):(1'h1)] : (~|($unsigned((8'haa)) ?
                              reg1401 : (forvar1475 & reg1444))));
                    end
                  for (forvar1510 = (1'h0); (forvar1510 < (2'h2)); forvar1510 = (forvar1510 + (1'h1)))
                    begin
                      reg1511 <= (forvar1501 ?
                          (reg1429[(5'h10):(3'h7)] ?
                              (reg1427[(3'h7):(1'h0)] >= reg1490[(3'h4):(2'h3)]) : (~|$unsigned(reg1463))) : (($signed(reg1487) + (reg1396 ?
                                  (8'hac) : reg1407)) ?
                              $unsigned(reg1486) : $signed($unsigned(wire1181))));
                    end
                end
            end
          for (forvar1512 = (1'h0); (forvar1512 < (2'h3)); forvar1512 = (forvar1512 + (1'h1)))
            begin
              reg1513 <= (reg1450[(2'h3):(1'h0)] <= $signed(((~|(8'ha7)) & (wire1182 ?
                  reg1386 : reg1506))));
              reg1514 <= ((~|(8'hb6)) ?
                  (&reg1395) : $signed(((reg1430 ?
                      reg1402 : reg1481) >> (|reg1458))));
              for (forvar1515 = (1'h0); (forvar1515 < (1'h0)); forvar1515 = (forvar1515 + (1'h1)))
                begin
                  for (forvar1516 = (1'h0); (forvar1516 < (1'h1)); forvar1516 = (forvar1516 + (1'h1)))
                    begin
                      reg1517 <= (-reg1423);
                      reg1518 <= (8'h9d);
                      reg1519 <= $signed((reg1453 ?
                          $unsigned($unsigned(forvar1512)) : $signed(reg1406)));
                    end
                  for (forvar1520 = (1'h0); (forvar1520 < (1'h0)); forvar1520 = (forvar1520 + (1'h1)))
                    begin
                      reg1521 <= reg1427;
                      reg1522 <= forvar1510[(1'h0):(1'h0)];
                    end
                end
              reg1523 <= $unsigned($unsigned(({(8'hb8)} == (forvar1496 > reg1430))));
            end
          reg1524 <= ((((reg1456 ? (8'hb0) : (8'h9d)) ?
              (reg1485 ?
                  reg1484 : reg1479) : (reg1433 & reg1505)) >= wire1373) >= reg1403);
        end
      else
        begin
          if ($unsigned((|reg1397)))
            begin
              for (forvar1475 = (1'h0); (forvar1475 < (1'h1)); forvar1475 = (forvar1475 + (1'h1)))
                begin
                  for (forvar1476 = (1'h0); (forvar1476 < (1'h0)); forvar1476 = (forvar1476 + (1'h1)))
                    begin
                      reg1477 <= (^$signed(reg1467));
                      reg1478 <= {(((reg1443 ? reg1406 : reg1447) ?
                                  reg1400[(4'ha):(4'ha)] : (reg1507 * reg1394)) ?
                              ($signed(reg1410) ~^ (reg1417 ?
                                  reg1376 : forvar1491)) : {reg1434[(3'h5):(1'h1)]})};
                      reg1479 <= ((^reg1381) ? reg1398 : (~(~&(+reg1381))));
                      reg1480 <= {reg1436[(1'h0):(1'h0)]};
                    end
                  for (forvar1481 = (1'h0); (forvar1481 < (2'h2)); forvar1481 = (forvar1481 + (1'h1)))
                    begin
                      reg1482 <= reg1473;
                      reg1483 <= $signed($unsigned(($signed(forvar1510) ?
                          $unsigned(reg1509) : reg1453[(4'hd):(4'h9)])));
                      reg1484 <= reg1486[(1'h1):(1'h1)];
                      reg1485 <= wire1373;
                    end
                end
            end
          else
            begin
              if (((|(&reg1522[(3'h7):(3'h5)])) + ((!$signed(forvar1503)) ?
                  (&reg1511[(3'h5):(2'h2)]) : $signed($signed(reg1378)))))
                begin
                  for (forvar1475 = (1'h0); (forvar1475 < (2'h2)); forvar1475 = (forvar1475 + (1'h1)))
                    begin
                      reg1476 <= forvar1508;
                      reg1477 <= (~|reg1463);
                      reg1478 <= (^(reg1401[(3'h5):(3'h4)] <= $signed($unsigned(forvar1483))));
                      reg1479 <= reg1387[(3'h5):(1'h1)];
                    end
                  reg1480 <= reg1416;
                  if (reg1444)
                    begin
                      reg1481 <= $signed((^{$signed(reg1442)}));
                    end
                  else
                    begin
                      reg1481 <= reg1384[(4'ha):(3'h6)];
                      reg1482 <= wire1375;
                      reg1483 <= reg1434[(3'h6):(3'h4)];
                    end
                  for (forvar1484 = (1'h0); (forvar1484 < (2'h2)); forvar1484 = (forvar1484 + (1'h1)))
                    begin
                      reg1485 <= (~^(^~$signed((reg1524 != forvar1516))));
                      reg1486 <= {$signed(reg1519)};
                    end
                end
              else
                begin
                  reg1475 <= wire1184;
                  if (forvar1483)
                    begin
                      reg1476 <= $unsigned(reg1405);
                      reg1477 <= reg1420[(4'hf):(2'h3)];
                    end
                  else
                    begin
                      reg1476 <= reg1437;
                      reg1477 <= $unsigned(((reg1398[(4'ha):(3'h6)] ?
                              (^~reg1487) : reg1468[(4'h9):(3'h6)]) ?
                          $signed((reg1433 ? (8'hac) : reg1429)) : reg1425));
                    end
                end
              for (forvar1487 = (1'h0); (forvar1487 < (2'h2)); forvar1487 = (forvar1487 + (1'h1)))
                begin
                  for (forvar1488 = (1'h0); (forvar1488 < (1'h1)); forvar1488 = (forvar1488 + (1'h1)))
                    begin
                      reg1489 <= {(forvar1502[(4'hd):(4'ha)] ?
                              (~^(reg1488 ?
                                  reg1427 : (8'hb9))) : (reg1500[(2'h2):(1'h0)] ?
                                  (forvar1520 & reg1460) : reg1403[(2'h2):(1'h1)]))};
                      reg1490 <= (($unsigned(reg1394) <<< (8'haa)) ?
                          $signed((~|(reg1388 ~^ reg1470))) : $unsigned($signed((~^wire1184))));
                    end
                  for (forvar1491 = (1'h0); (forvar1491 < (1'h1)); forvar1491 = (forvar1491 + (1'h1)))
                    begin
                      reg1492 <= {{reg1389}};
                      reg1493 <= (~&{reg1461});
                      reg1494 <= ($signed(reg1467[(1'h1):(1'h1)]) ?
                          $unsigned(reg1442[(3'h7):(1'h1)]) : $unsigned(reg1476[(3'h6):(3'h6)]));
                      reg1495 <= (reg1405[(3'h4):(2'h3)] - $unsigned((reg1402[(4'ha):(3'h6)] >> ((8'ha2) ?
                          reg1518 : reg1397))));
                    end
                  for (forvar1496 = (1'h0); (forvar1496 < (1'h0)); forvar1496 = (forvar1496 + (1'h1)))
                    begin
                      reg1497 <= reg1417;
                      reg1498 <= (~^((reg1386[(2'h3):(1'h1)] != (^~reg1394)) ?
                          $unsigned(forvar1488[(4'ha):(3'h6)]) : reg1385));
                    end
                end
              reg1499 <= (forvar1520[(4'h8):(2'h3)] + $unsigned($unsigned({reg1518})));
            end
          for (forvar1500 = (1'h0); (forvar1500 < (1'h0)); forvar1500 = (forvar1500 + (1'h1)))
            begin
              for (forvar1501 = (1'h0); (forvar1501 < (1'h1)); forvar1501 = (forvar1501 + (1'h1)))
                begin
                  reg1502 <= reg1484[(1'h1):(1'h1)];
                  if ($unsigned(forvar1512[(3'h5):(3'h5)]))
                    begin
                      reg1503 <= ((-((reg1414 >= reg1452) ?
                              (reg1506 ^ reg1485) : $unsigned(reg1445))) ?
                          $signed(reg1423[(4'he):(3'h4)]) : reg1479);
                    end
                  else
                    begin
                      reg1503 <= $unsigned($unsigned(reg1499[(3'h4):(2'h3)]));
                      reg1504 <= reg1394[(2'h3):(1'h1)];
                      reg1505 <= {$unsigned({(reg1441 && forvar1520)})};
                    end
                  for (forvar1506 = (1'h0); (forvar1506 < (1'h0)); forvar1506 = (forvar1506 + (1'h1)))
                    begin
                      reg1507 <= (~(-forvar1483[(1'h0):(1'h0)]));
                      reg1508 <= (reg1487[(4'h8):(3'h5)] >>> $unsigned($unsigned((forvar1515 ?
                          forvar1484 : reg1523))));
                      reg1509 <= $unsigned($signed((!(reg1379 ?
                          (8'hba) : reg1498))));
                    end
                end
              for (forvar1510 = (1'h0); (forvar1510 < (1'h1)); forvar1510 = (forvar1510 + (1'h1)))
                begin
                  if (((~^{(reg1445 ?
                          reg1514 : (8'hab))}) >>> reg1518[(1'h0):(1'h0)]))
                    begin
                      reg1511 <= $signed($signed(reg1478));
                      reg1512 <= $signed(reg1466[(4'hc):(4'h9)]);
                    end
                  else
                    begin
                      reg1511 <= reg1473;
                    end
                end
              reg1513 <= $unsigned(($unsigned((wire1471 ? reg1518 : reg1436)) ?
                  wire1184[(1'h1):(1'h0)] : (reg1487 ?
                      (~|reg1478) : $signed(wire1472))));
              if ($unsigned($signed($unsigned($signed(reg1521)))))
                begin
                  for (forvar1514 = (1'h0); (forvar1514 < (1'h1)); forvar1514 = (forvar1514 + (1'h1)))
                    begin
                      reg1515 <= $signed(({reg1466[(4'ha):(3'h4)]} == (forvar1500[(1'h1):(1'h0)] ?
                          reg1390[(3'h4):(3'h4)] : (reg1518 == (8'hae)))));
                      reg1516 <= ($unsigned({$signed(forvar1478)}) ?
                          (($unsigned(reg1483) >> $signed(reg1446)) ?
                              reg1429[(3'h4):(1'h0)] : ($signed((8'hba)) ?
                                  $unsigned(reg1458) : (reg1379 ?
                                      reg1480 : reg1481))) : (8'hb6));
                    end
                end
              else
                begin
                  for (forvar1514 = (1'h0); (forvar1514 < (2'h3)); forvar1514 = (forvar1514 + (1'h1)))
                    begin
                      reg1515 <= (8'hb9);
                    end
                  if ({$signed({(forvar1475 + reg1476)})})
                    begin
                      reg1516 <= (!forvar1506[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1516 <= ({$unsigned($signed(reg1382))} ?
                          wire1185 : $unsigned($unsigned(reg1396)));
                    end
                end
            end
        end
    end
  assign wire1525 = reg1436[(4'h8):(3'h4)];
  assign wire1526 = reg1404;
  assign wire1527 = (-(-((^reg1504) | (wire1185 << reg1509))));
  assign wire1528 = $signed({((~^reg1395) ? reg1432 : reg1512)});
  assign wire1529 = $signed((-(~(reg1499 <<< reg1457))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1187  (y, clk, wire1191, wire1190, wire1189, wire1188);
  output wire [(32'h87a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire1191;
  input wire signed [(3'h5):(1'h0)] wire1190;
  input wire [(4'hf):(1'h0)] wire1189;
  input wire [(4'hb):(1'h0)] wire1188;
  wire [(4'he):(1'h0)] wire1372;
  wire signed [(3'h5):(1'h0)] wire1371;
  wire [(5'h10):(1'h0)] wire1370;
  wire [(3'h5):(1'h0)] wire1250;
  wire [(5'h10):(1'h0)] wire1249;
  wire signed [(4'hb):(1'h0)] wire1248;
  wire [(4'ha):(1'h0)] wire1247;
  wire [(4'hd):(1'h0)] wire1193;
  wire signed [(4'hb):(1'h0)] wire1192;
  reg [(4'hd):(1'h0)] reg1364 = (1'h0);
  reg [(3'h6):(1'h0)] reg1369 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1368 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1367 = (1'h0);
  reg [(4'ha):(1'h0)] reg1366 = (1'h0);
  reg [(4'h8):(1'h0)] reg1365 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1363 = (1'h0);
  reg [(4'h8):(1'h0)] reg1362 = (1'h0);
  reg [(5'h10):(1'h0)] reg1361 = (1'h0);
  reg [(4'he):(1'h0)] reg1360 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1359 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1346 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1343 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1335 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1334 = (1'h0);
  reg [(3'h5):(1'h0)] reg1358 = (1'h0);
  reg [(4'ha):(1'h0)] reg1357 = (1'h0);
  reg [(3'h5):(1'h0)] reg1356 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1355 = (1'h0);
  reg [(4'hb):(1'h0)] reg1353 = (1'h0);
  reg [(4'h9):(1'h0)] reg1352 = (1'h0);
  reg [(4'he):(1'h0)] reg1349 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1348 = (1'h0);
  reg [(4'ha):(1'h0)] reg1347 = (1'h0);
  reg [(4'ha):(1'h0)] reg1345 = (1'h0);
  reg [(4'h9):(1'h0)] reg1344 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1342 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1341 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1340 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1339 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1338 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1337 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1336 = (1'h0);
  reg [(3'h7):(1'h0)] reg1316 = (1'h0);
  reg [(3'h4):(1'h0)] reg1300 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1295 = (1'h0);
  reg [(2'h3):(1'h0)] reg1333 = (1'h0);
  reg [(4'hf):(1'h0)] reg1332 = (1'h0);
  reg [(4'h8):(1'h0)] reg1331 = (1'h0);
  reg [(3'h7):(1'h0)] reg1330 = (1'h0);
  reg [(4'hc):(1'h0)] reg1328 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1326 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1324 = (1'h0);
  reg [(4'ha):(1'h0)] reg1323 = (1'h0);
  reg [(4'hb):(1'h0)] reg1322 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1321 = (1'h0);
  reg [(4'hb):(1'h0)] reg1313 = (1'h0);
  reg [(5'h10):(1'h0)] reg1320 = (1'h0);
  reg [(4'h8):(1'h0)] reg1319 = (1'h0);
  reg [(4'ha):(1'h0)] reg1318 = (1'h0);
  reg [(2'h3):(1'h0)] reg1317 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1315 = (1'h0);
  reg [(3'h5):(1'h0)] reg1314 = (1'h0);
  reg [(4'hd):(1'h0)] reg1304 = (1'h0);
  reg [(4'hd):(1'h0)] reg1312 = (1'h0);
  reg [(4'hd):(1'h0)] reg1311 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1310 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1309 = (1'h0);
  reg [(5'h10):(1'h0)] reg1308 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1307 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1306 = (1'h0);
  reg [(4'hf):(1'h0)] reg1305 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1303 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1302 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1301 = (1'h0);
  reg [(4'hc):(1'h0)] reg1299 = (1'h0);
  reg [(3'h6):(1'h0)] reg1298 = (1'h0);
  reg [(4'hb):(1'h0)] reg1297 = (1'h0);
  reg [(3'h6):(1'h0)] reg1296 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1294 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1293 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1292 = (1'h0);
  reg [(3'h4):(1'h0)] reg1291 = (1'h0);
  reg [(3'h7):(1'h0)] reg1290 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1289 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1287 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1286 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1284 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1283 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1282 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1281 = (1'h0);
  reg [(4'hf):(1'h0)] reg1271 = (1'h0);
  reg [(2'h3):(1'h0)] reg1279 = (1'h0);
  reg [(2'h3):(1'h0)] reg1278 = (1'h0);
  reg [(2'h3):(1'h0)] reg1277 = (1'h0);
  reg [(2'h2):(1'h0)] reg1276 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1267 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1260 = (1'h0);
  reg [(2'h3):(1'h0)] reg1255 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1262 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1275 = (1'h0);
  reg [(4'hf):(1'h0)] reg1274 = (1'h0);
  reg [(4'hb):(1'h0)] reg1273 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1272 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1270 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1269 = (1'h0);
  reg [(3'h7):(1'h0)] reg1268 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1266 = (1'h0);
  reg [(4'h9):(1'h0)] reg1265 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1264 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1263 = (1'h0);
  reg [(4'hf):(1'h0)] reg1251 = (1'h0);
  reg [(5'h10):(1'h0)] reg1261 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1259 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1258 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1257 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1256 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1254 = (1'h0);
  reg [(3'h4):(1'h0)] reg1253 = (1'h0);
  reg [(5'h10):(1'h0)] reg1252 = (1'h0);
  reg [(3'h5):(1'h0)] reg1230 = (1'h0);
  reg [(4'h8):(1'h0)] reg1246 = (1'h0);
  reg [(4'ha):(1'h0)] reg1245 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1244 = (1'h0);
  reg [(2'h3):(1'h0)] reg1243 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1240 = (1'h0);
  reg [(3'h6):(1'h0)] reg1236 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1242 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1241 = (1'h0);
  reg [(3'h5):(1'h0)] reg1239 = (1'h0);
  reg [(4'h8):(1'h0)] reg1238 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1237 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1235 = (1'h0);
  reg [(4'he):(1'h0)] reg1234 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1233 = (1'h0);
  reg [(4'hb):(1'h0)] reg1232 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1231 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1229 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1228 = (1'h0);
  reg [(2'h3):(1'h0)] reg1227 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1226 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1223 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1195 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1216 = (1'h0);
  reg [(4'ha):(1'h0)] reg1207 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1204 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1196 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1194 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1221 = (1'h0);
  reg [(2'h3):(1'h0)] reg1220 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1219 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1218 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1217 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1215 = (1'h0);
  reg [(3'h4):(1'h0)] reg1214 = (1'h0);
  reg [(3'h4):(1'h0)] reg1213 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1212 = (1'h0);
  reg [(3'h6):(1'h0)] reg1211 = (1'h0);
  reg [(4'he):(1'h0)] reg1210 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1209 = (1'h0);
  reg [(4'h9):(1'h0)] reg1208 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1206 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1205 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1203 = (1'h0);
  reg [(3'h4):(1'h0)] reg1202 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1201 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1200 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1199 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1198 = (1'h0);
  reg [(4'h9):(1'h0)] reg1197 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1360 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1363 = (1'h0);
  reg [(4'he):(1'h0)] forvar1364 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1359 = (1'h0);
  reg [(4'he):(1'h0)] forvar1345 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1354 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1351 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1350 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1346 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1343 = (1'h0);
  reg [(4'he):(1'h0)] forvar1335 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1334 = (1'h0);
  reg [(4'he):(1'h0)] forvar1315 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1312 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1308 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1306 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1301 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1296 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1329 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1327 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1325 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1316 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1313 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1307 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1304 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1300 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1295 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1288 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1285 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1283 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1280 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1272 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1266 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1275 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1270 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1265 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1261 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1258 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1256 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1254 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1271 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1267 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1262 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1252 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1260 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1255 = (1'h0);
  reg [(4'he):(1'h0)] forvar1251 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1242 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1237 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1229 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1235 = (1'h0);
  reg [(4'he):(1'h0)] forvar1240 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1236 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1230 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1225 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1224 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1222 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1200 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1214 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1211 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1208 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1205 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1203 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1198 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1216 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1207 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1204 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1196 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1195 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1194 = (1'h0);
  assign y = {wire1372,
                 wire1371,
                 wire1370,
                 wire1250,
                 wire1249,
                 wire1248,
                 wire1247,
                 wire1193,
                 wire1192,
                 reg1364,
                 reg1369,
                 reg1368,
                 reg1367,
                 reg1366,
                 reg1365,
                 reg1363,
                 reg1362,
                 reg1361,
                 reg1360,
                 reg1359,
                 reg1346,
                 reg1343,
                 reg1335,
                 reg1334,
                 reg1358,
                 reg1357,
                 reg1356,
                 reg1355,
                 reg1353,
                 reg1352,
                 reg1349,
                 reg1348,
                 reg1347,
                 reg1345,
                 reg1344,
                 reg1342,
                 reg1341,
                 reg1340,
                 reg1339,
                 reg1338,
                 reg1337,
                 reg1336,
                 reg1316,
                 reg1300,
                 reg1295,
                 reg1333,
                 reg1332,
                 reg1331,
                 reg1330,
                 reg1328,
                 reg1326,
                 reg1324,
                 reg1323,
                 reg1322,
                 reg1321,
                 reg1313,
                 reg1320,
                 reg1319,
                 reg1318,
                 reg1317,
                 reg1315,
                 reg1314,
                 reg1304,
                 reg1312,
                 reg1311,
                 reg1310,
                 reg1309,
                 reg1308,
                 reg1307,
                 reg1306,
                 reg1305,
                 reg1303,
                 reg1302,
                 reg1301,
                 reg1299,
                 reg1298,
                 reg1297,
                 reg1296,
                 reg1294,
                 reg1293,
                 reg1292,
                 reg1291,
                 reg1290,
                 reg1289,
                 reg1287,
                 reg1286,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1281,
                 reg1271,
                 reg1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 reg1267,
                 reg1260,
                 reg1255,
                 reg1262,
                 reg1275,
                 reg1274,
                 reg1273,
                 reg1272,
                 reg1270,
                 reg1269,
                 reg1268,
                 reg1266,
                 reg1265,
                 reg1264,
                 reg1263,
                 reg1251,
                 reg1261,
                 reg1259,
                 reg1258,
                 reg1257,
                 reg1256,
                 reg1254,
                 reg1253,
                 reg1252,
                 reg1230,
                 reg1246,
                 reg1245,
                 reg1244,
                 reg1243,
                 reg1240,
                 reg1236,
                 reg1242,
                 reg1241,
                 reg1239,
                 reg1238,
                 reg1237,
                 reg1235,
                 reg1234,
                 reg1233,
                 reg1232,
                 reg1231,
                 reg1229,
                 reg1228,
                 reg1227,
                 reg1226,
                 reg1223,
                 reg1195,
                 reg1216,
                 reg1207,
                 reg1204,
                 reg1196,
                 reg1194,
                 reg1221,
                 reg1220,
                 reg1219,
                 reg1218,
                 reg1217,
                 reg1215,
                 reg1214,
                 reg1213,
                 reg1212,
                 reg1211,
                 reg1210,
                 reg1209,
                 reg1208,
                 reg1206,
                 reg1205,
                 reg1203,
                 reg1202,
                 reg1201,
                 reg1200,
                 reg1199,
                 reg1198,
                 reg1197,
                 forvar1360,
                 forvar1363,
                 forvar1364,
                 forvar1359,
                 forvar1345,
                 forvar1354,
                 forvar1351,
                 forvar1350,
                 forvar1346,
                 forvar1343,
                 forvar1335,
                 forvar1334,
                 forvar1315,
                 forvar1312,
                 forvar1308,
                 forvar1306,
                 forvar1301,
                 forvar1296,
                 forvar1329,
                 forvar1327,
                 forvar1325,
                 forvar1316,
                 forvar1313,
                 forvar1307,
                 forvar1304,
                 forvar1300,
                 forvar1295,
                 forvar1288,
                 forvar1285,
                 forvar1283,
                 forvar1280,
                 forvar1272,
                 forvar1266,
                 forvar1275,
                 forvar1270,
                 forvar1265,
                 forvar1261,
                 forvar1258,
                 forvar1256,
                 forvar1254,
                 forvar1271,
                 forvar1267,
                 forvar1262,
                 forvar1252,
                 forvar1260,
                 forvar1255,
                 forvar1251,
                 forvar1242,
                 forvar1237,
                 forvar1229,
                 forvar1235,
                 forvar1240,
                 forvar1236,
                 forvar1230,
                 forvar1225,
                 forvar1224,
                 forvar1222,
                 forvar1200,
                 forvar1214,
                 forvar1211,
                 forvar1208,
                 forvar1205,
                 forvar1203,
                 forvar1198,
                 forvar1216,
                 forvar1207,
                 forvar1204,
                 forvar1196,
                 forvar1195,
                 forvar1194,
                 (1'h0)};
  assign wire1192 = {(((wire1189 ? wire1191 : wire1190) ?
                                wire1189 : (wire1190 ? wire1189 : (8'hb6))) ?
                            (wire1189 ?
                                {wire1189} : ((8'hb3) == (8'hb0))) : {$unsigned(wire1191)})};
  assign wire1193 = ((8'hb0) || wire1190[(3'h4):(2'h2)]);
  always
    @(posedge clk) begin
      if (wire1193)
        begin
          for (forvar1194 = (1'h0); (forvar1194 < (2'h2)); forvar1194 = (forvar1194 + (1'h1)))
            begin
              for (forvar1195 = (1'h0); (forvar1195 < (1'h0)); forvar1195 = (forvar1195 + (1'h1)))
                begin
                  for (forvar1196 = (1'h0); (forvar1196 < (1'h0)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 <= $signed(((wire1193[(4'hd):(1'h1)] >>> $unsigned((8'hb0))) * (8'hac)));
                      reg1198 <= $unsigned(wire1193[(4'hb):(4'h8)]);
                      reg1199 <= {forvar1195[(3'h4):(3'h4)]};
                    end
                  if ({{$signed(wire1189[(4'hf):(3'h7)])}})
                    begin
                      reg1200 <= $unsigned((~($unsigned(forvar1195) ?
                          $unsigned(wire1188) : $signed(wire1193))));
                      reg1201 <= $signed({($signed((8'haa)) ?
                              reg1197 : $signed(forvar1195))});
                      reg1202 <= (~|reg1198[(2'h2):(1'h0)]);
                      reg1203 <= forvar1196;
                    end
                  else
                    begin
                      reg1200 <= $unsigned((~|{(wire1193 ?
                              wire1191 : wire1189)}));
                      reg1201 <= {$signed((!(^~forvar1196)))};
                      reg1202 <= ((($signed((8'ha2)) >> $unsigned((8'ha2))) ?
                          $signed({wire1189}) : $unsigned((~^wire1191))) || {(~|forvar1194)});
                      reg1203 <= reg1197;
                    end
                  for (forvar1204 = (1'h0); (forvar1204 < (2'h2)); forvar1204 = (forvar1204 + (1'h1)))
                    begin
                      reg1205 <= ($unsigned((~&$unsigned(forvar1195))) >> (8'ha0));
                      reg1206 <= (-$signed(((~^reg1201) < (reg1201 ?
                          wire1191 : wire1192))));
                    end
                  for (forvar1207 = (1'h0); (forvar1207 < (2'h2)); forvar1207 = (forvar1207 + (1'h1)))
                    begin
                      reg1208 <= ($unsigned($signed((forvar1207 ?
                          reg1205 : wire1188))) >> wire1190[(2'h3):(2'h3)]);
                      reg1209 <= ({reg1208} ?
                          $signed((~^forvar1196[(3'h7):(3'h6)])) : (wire1192 ?
                              $signed(forvar1195) : (reg1203[(4'ha):(3'h7)] + (+wire1188))));
                      reg1210 <= {{((reg1205 != reg1198) ?
                                  {reg1198} : $signed(forvar1204))}};
                    end
                end
              reg1211 <= {$unsigned(((-reg1209) ?
                      (wire1191 << forvar1194) : $signed(reg1201)))};
              if ($signed(reg1208[(3'h7):(3'h4)]))
                begin
                  if (reg1203)
                    begin
                      reg1212 <= (^~{$unsigned({forvar1196})});
                      reg1213 <= reg1203;
                    end
                  else
                    begin
                      reg1212 <= reg1203;
                      reg1213 <= ($signed(({wire1192} * $signed(forvar1195))) || reg1201[(2'h2):(2'h2)]);
                    end
                  reg1214 <= ($unsigned(wire1190) <= {($unsigned(reg1213) ?
                          $signed(reg1212) : (forvar1194 >> forvar1207))});
                end
              else
                begin
                  if (reg1211[(1'h1):(1'h0)])
                    begin
                      reg1212 <= $unsigned(reg1214);
                      reg1213 <= {{(~|(!reg1208))}};
                      reg1214 <= wire1191;
                    end
                  else
                    begin
                      reg1212 <= (+{$unsigned($signed((8'hba)))});
                      reg1213 <= $signed((({(8'hab)} + (|reg1205)) ?
                          (+(+reg1208)) : wire1191[(4'hf):(4'hf)]));
                      reg1214 <= (reg1209[(2'h2):(2'h2)] ?
                          ($signed((8'haa)) * reg1201[(1'h0):(1'h0)]) : $signed(((~(8'hae)) ?
                              wire1188 : (reg1208 ^~ wire1191))));
                      reg1215 <= (((reg1202 ?
                                  reg1211[(2'h3):(1'h1)] : (reg1209 >>> forvar1195)) ?
                              $signed((forvar1194 ?
                                  wire1193 : forvar1207)) : (&((8'ha9) ^ wire1192))) ?
                          reg1199 : wire1190);
                    end
                  for (forvar1216 = (1'h0); (forvar1216 < (2'h2)); forvar1216 = (forvar1216 + (1'h1)))
                    begin
                      reg1217 <= ($signed(reg1203) > $unsigned(((~&wire1189) ?
                          (8'haa) : $signed(reg1202))));
                      reg1218 <= $unsigned($unsigned((reg1203[(4'h9):(3'h5)] * $unsigned(reg1215))));
                      reg1219 <= $signed({reg1200[(4'h9):(2'h3)]});
                      reg1220 <= $signed({({reg1219} ?
                              $signed(reg1203) : $unsigned(forvar1195))});
                    end
                  reg1221 <= ((forvar1194 ?
                          reg1211 : ({reg1219} | $signed(wire1192))) ?
                      reg1214 : forvar1207);
                end
            end
        end
      else
        begin
          reg1194 <= (8'hb5);
          if ((+($signed((forvar1196 ~^ forvar1194)) ?
              $signed(reg1212[(1'h1):(1'h1)]) : (&(+reg1200)))))
            begin
              for (forvar1195 = (1'h0); (forvar1195 < (1'h0)); forvar1195 = (forvar1195 + (1'h1)))
                begin
                  reg1196 <= forvar1207[(3'h5):(2'h2)];
                end
              if (reg1211[(3'h6):(1'h0)])
                begin
                  reg1197 <= reg1220;
                  for (forvar1198 = (1'h0); (forvar1198 < (2'h3)); forvar1198 = (forvar1198 + (1'h1)))
                    begin
                      reg1199 <= $signed($unsigned({$signed((8'ha3))}));
                      reg1200 <= ((!(8'hae)) & (reg1194[(3'h7):(3'h5)] * ((-reg1199) ^~ ((8'hb1) ?
                          reg1210 : reg1200))));
                      reg1201 <= wire1192;
                      reg1202 <= ((forvar1204[(1'h0):(1'h0)] ?
                          $unsigned($signed(reg1198)) : ((!forvar1207) * (reg1217 >>> reg1212))) ~^ (reg1203[(1'h1):(1'h1)] >>> (&(~&wire1191))));
                    end
                  for (forvar1203 = (1'h0); (forvar1203 < (1'h1)); forvar1203 = (forvar1203 + (1'h1)))
                    begin
                      reg1204 <= $unsigned(wire1193[(4'hd):(2'h2)]);
                    end
                  for (forvar1205 = (1'h0); (forvar1205 < (1'h1)); forvar1205 = (forvar1205 + (1'h1)))
                    begin
                      reg1206 <= (^~(~$signed($signed((8'hab)))));
                      reg1207 <= (~^forvar1207[(2'h2):(1'h1)]);
                    end
                end
              else
                begin
                  if (reg1218[(4'hb):(4'ha)])
                    begin
                      reg1197 <= $signed((((reg1203 ?
                              (8'hab) : reg1201) ~^ $signed((8'hae))) ?
                          $signed((wire1190 ?
                              forvar1207 : (8'hb0))) : reg1198));
                      reg1198 <= ($unsigned(reg1203[(4'h9):(3'h5)]) ?
                          forvar1196 : reg1207[(2'h3):(1'h0)]);
                      reg1199 <= forvar1205[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1197 <= (reg1199[(3'h4):(2'h3)] & {$signed((wire1193 <<< (8'ha1)))});
                      reg1198 <= ($unsigned(reg1212) ?
                          {(^~(8'h9f))} : reg1213[(1'h0):(1'h0)]);
                    end
                end
              for (forvar1208 = (1'h0); (forvar1208 < (1'h1)); forvar1208 = (forvar1208 + (1'h1)))
                begin
                  if ((({(reg1199 <= (8'ha1))} <<< reg1203[(3'h4):(1'h0)]) > {$unsigned($unsigned(reg1209))}))
                    begin
                      reg1209 <= (($unsigned(forvar1203) <= (+reg1196)) * ((((8'hb8) <= reg1208) ?
                          reg1218 : $unsigned(reg1194)) != $unsigned((~^reg1196))));
                      reg1210 <= forvar1194[(3'h7):(2'h3)];
                    end
                  else
                    begin
                      reg1209 <= ($unsigned(wire1191[(4'hb):(2'h2)]) ?
                          (((!forvar1204) ?
                                  $unsigned(forvar1205) : ((8'hb9) || reg1219)) ?
                              $unsigned($signed(reg1200)) : ($signed(forvar1195) ?
                                  reg1213 : $signed(forvar1204))) : {(8'ha3)});
                    end
                  for (forvar1211 = (1'h0); (forvar1211 < (1'h0)); forvar1211 = (forvar1211 + (1'h1)))
                    begin
                      reg1212 <= ($signed(((reg1208 <= (8'ha6)) ~^ $unsigned(reg1220))) & ({reg1221[(1'h0):(1'h0)]} <= reg1199[(2'h2):(2'h2)]));
                      reg1213 <= reg1198[(3'h7):(1'h1)];
                    end
                  for (forvar1214 = (1'h0); (forvar1214 < (2'h2)); forvar1214 = (forvar1214 + (1'h1)))
                    begin
                      reg1215 <= (~|(^reg1210));
                      reg1216 <= $unsigned($unsigned((((8'ha6) ?
                              reg1200 : reg1218) ?
                          wire1188 : reg1200)));
                      reg1217 <= {(&$signed(((8'ha3) ? reg1221 : reg1207)))};
                      reg1218 <= (({(|reg1194)} ^~ (8'hb4)) < $unsigned($unsigned((~|reg1212))));
                    end
                end
            end
          else
            begin
              if (forvar1198[(4'hc):(3'h6)])
                begin
                  reg1195 <= wire1189[(3'h6):(3'h5)];
                end
              else
                begin
                  if ({forvar1208[(1'h1):(1'h0)]})
                    begin
                      reg1195 <= forvar1198[(1'h0):(1'h0)];
                      reg1196 <= (wire1188 ~^ ((~(wire1191 ?
                          reg1217 : reg1195)) + ($signed(forvar1204) != $unsigned(wire1191))));
                      reg1197 <= (($signed((reg1217 ?
                              wire1191 : reg1216)) || reg1217) ?
                          (^~(^(reg1213 >> reg1213))) : (((~^wire1191) ?
                              (^~(8'hb4)) : wire1191[(4'hf):(2'h3)]) + (-forvar1195)));
                      reg1198 <= (((wire1191[(3'h4):(1'h0)] ?
                              $unsigned(reg1197) : (reg1215 & reg1195)) <<< reg1221[(2'h3):(1'h1)]) ?
                          $unsigned((+$signed((8'hae)))) : (~&((-reg1217) >> (forvar1196 >> reg1205))));
                    end
                  else
                    begin
                      reg1195 <= forvar1216[(2'h2):(1'h1)];
                      reg1196 <= reg1205;
                    end
                end
              reg1199 <= ($signed($signed($signed(reg1211))) ?
                  $signed({{reg1214}}) : (($signed((8'ha6)) & (~reg1220)) ?
                      $signed((wire1189 ^ forvar1211)) : reg1204));
              for (forvar1200 = (1'h0); (forvar1200 < (1'h0)); forvar1200 = (forvar1200 + (1'h1)))
                begin
                  if (((8'ha2) ?
                      (8'ha9) : $unsigned((forvar1208[(4'h9):(1'h1)] >> (reg1212 || (8'ha9))))))
                    begin
                      reg1201 <= {(^(~|$signed(forvar1200)))};
                      reg1202 <= $signed(($unsigned($unsigned(wire1192)) || ((forvar1205 ?
                          reg1205 : (8'h9f)) ^ forvar1203[(3'h6):(1'h0)])));
                      reg1203 <= ((^~$signed({reg1212})) ?
                          (~forvar1203) : wire1193[(3'h6):(2'h3)]);
                      reg1204 <= {forvar1198};
                    end
                  else
                    begin
                      reg1201 <= (8'haf);
                      reg1202 <= (forvar1198[(4'hd):(4'hd)] ?
                          forvar1196[(1'h1):(1'h0)] : (((reg1218 ?
                                      (8'hb3) : forvar1194) ?
                                  (reg1216 ?
                                      reg1217 : wire1188) : reg1220[(1'h1):(1'h0)]) ?
                              (!$unsigned(reg1205)) : $unsigned(reg1203)));
                      reg1203 <= forvar1200[(2'h3):(1'h0)];
                      reg1204 <= (-($unsigned($unsigned(reg1212)) ?
                          {$unsigned(reg1215)} : {(8'ha6)}));
                    end
                end
              if (((((forvar1216 <<< (8'ha6)) ?
                      ((8'hb8) ? reg1206 : (8'h9f)) : (reg1195 ?
                          forvar1214 : reg1217)) && reg1221[(2'h2):(1'h0)]) ?
                  forvar1211[(2'h2):(2'h2)] : forvar1198[(1'h0):(1'h0)]))
                begin
                  if ($unsigned(reg1202[(1'h0):(1'h0)]))
                    begin
                      reg1205 <= reg1197[(3'h5):(2'h3)];
                      reg1206 <= ((~{$unsigned(reg1219)}) ?
                          $unsigned($unsigned($unsigned(reg1215))) : $unsigned(reg1197));
                    end
                  else
                    begin
                      reg1205 <= (~&$signed((reg1195 ^ reg1214)));
                    end
                  for (forvar1207 = (1'h0); (forvar1207 < (2'h2)); forvar1207 = (forvar1207 + (1'h1)))
                    begin
                      reg1208 <= reg1215;
                      reg1209 <= (~(($signed(forvar1205) <= $signed(reg1205)) ?
                          forvar1205[(4'h9):(2'h3)] : wire1188));
                      reg1210 <= $signed(($signed(reg1221) && ($unsigned(reg1218) != $unsigned(reg1218))));
                    end
                  for (forvar1211 = (1'h0); (forvar1211 < (2'h2)); forvar1211 = (forvar1211 + (1'h1)))
                    begin
                      reg1212 <= reg1213;
                      reg1213 <= (forvar1194 ?
                          ($unsigned((+reg1206)) ?
                              $unsigned($signed((8'hb3))) : reg1211) : forvar1203);
                      reg1214 <= $signed($unsigned(($signed((8'hb7)) ?
                          (reg1210 <<< forvar1198) : (~&(8'hab)))));
                    end
                end
              else
                begin
                  for (forvar1205 = (1'h0); (forvar1205 < (2'h2)); forvar1205 = (forvar1205 + (1'h1)))
                    begin
                      reg1206 <= ($signed(((^forvar1195) ?
                          ((8'hb7) ?
                              forvar1211 : reg1202) : (-forvar1211))) >>> $unsigned(forvar1211[(1'h1):(1'h0)]));
                    end
                  reg1207 <= reg1217[(4'hd):(4'hb)];
                  for (forvar1208 = (1'h0); (forvar1208 < (2'h3)); forvar1208 = (forvar1208 + (1'h1)))
                    begin
                      reg1209 <= (~forvar1208[(3'h7):(3'h7)]);
                      reg1210 <= $unsigned(wire1191);
                    end
                  if (reg1217[(3'h4):(2'h3)])
                    begin
                      reg1211 <= $unsigned($unsigned({reg1212}));
                      reg1212 <= $unsigned($signed((!(reg1217 - wire1193))));
                      reg1213 <= (8'hb1);
                    end
                  else
                    begin
                      reg1211 <= {({wire1188} ?
                              reg1212 : (^~$signed((8'ha9))))};
                      reg1212 <= wire1189;
                    end
                end
            end
        end
      for (forvar1222 = (1'h0); (forvar1222 < (1'h1)); forvar1222 = (forvar1222 + (1'h1)))
        begin
          reg1223 <= (8'ha1);
          if ($signed((reg1195[(4'hc):(4'h8)] ?
              reg1209[(2'h2):(1'h1)] : $signed($signed(wire1190)))))
            begin
              for (forvar1224 = (1'h0); (forvar1224 < (1'h1)); forvar1224 = (forvar1224 + (1'h1)))
                begin
                  for (forvar1225 = (1'h0); (forvar1225 < (1'h1)); forvar1225 = (forvar1225 + (1'h1)))
                    begin
                      reg1226 <= ($signed((8'hb6)) - (|reg1204));
                    end
                  if (reg1198)
                    begin
                      reg1227 <= (($unsigned({(8'hb0)}) != {(forvar1207 ~^ reg1194)}) ?
                          $signed((^(reg1223 ?
                              reg1221 : forvar1211))) : (~^(~|$signed(reg1217))));
                    end
                  else
                    begin
                      reg1227 <= $signed(((reg1220 ?
                          (~|reg1209) : (&reg1226)) - wire1189[(4'hd):(3'h6)]));
                      reg1228 <= $signed({reg1219[(3'h7):(1'h0)]});
                      reg1229 <= reg1201[(3'h6):(3'h6)];
                    end
                  for (forvar1230 = (1'h0); (forvar1230 < (2'h2)); forvar1230 = (forvar1230 + (1'h1)))
                    begin
                      reg1231 <= reg1208;
                      reg1232 <= ($signed((-reg1216)) ?
                          (~&(~&(~|(8'hb2)))) : (~({forvar1214} + (+forvar1203))));
                    end
                  reg1233 <= ($unsigned(forvar1194) ?
                      (8'haf) : (~^(reg1216[(1'h0):(1'h0)] ?
                          reg1216 : (forvar1207 ? forvar1200 : reg1205))));
                end
              reg1234 <= ((|(+(forvar1208 ~^ wire1188))) >= ($signed((reg1198 << (8'ha7))) ?
                  ((reg1205 <= reg1212) > $signed(forvar1225)) : (reg1214 ?
                      forvar1224[(1'h0):(1'h0)] : (forvar1216 ?
                          reg1231 : reg1195))));
              if (forvar1224[(2'h2):(1'h1)])
                begin
                  reg1235 <= (reg1204 ?
                      reg1203[(4'hb):(2'h2)] : $signed(($signed(reg1223) ?
                          ((8'ha0) ? forvar1207 : reg1219) : (8'ha2))));
                  for (forvar1236 = (1'h0); (forvar1236 < (1'h1)); forvar1236 = (forvar1236 + (1'h1)))
                    begin
                      reg1237 <= (reg1227 <= reg1207);
                      reg1238 <= reg1223[(3'h5):(3'h4)];
                      reg1239 <= ($unsigned($unsigned($signed(reg1216))) ~^ $unsigned($unsigned(reg1205)));
                    end
                  for (forvar1240 = (1'h0); (forvar1240 < (2'h3)); forvar1240 = (forvar1240 + (1'h1)))
                    begin
                      reg1241 <= $unsigned(forvar1205[(1'h0):(1'h0)]);
                      reg1242 <= reg1234[(3'h5):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar1235 = (1'h0); (forvar1235 < (2'h3)); forvar1235 = (forvar1235 + (1'h1)))
                    begin
                      reg1236 <= $signed((+$unsigned((~reg1239))));
                    end
                  if ($signed((reg1194[(2'h3):(2'h2)] && {reg1201[(3'h5):(2'h3)]})))
                    begin
                      reg1237 <= $signed(reg1238);
                      reg1238 <= ($unsigned(forvar1225[(1'h0):(1'h0)]) + ($unsigned((forvar1203 >>> reg1227)) ?
                          {$signed((8'hb7))} : ($unsigned(reg1235) >= forvar1236[(3'h7):(2'h3)])));
                      reg1239 <= (^{$unsigned((|forvar1225))});
                      reg1240 <= ((&(~^$unsigned(reg1221))) != (wire1190[(3'h4):(2'h3)] ?
                          reg1197[(3'h4):(2'h3)] : ({reg1239} < ((8'hb2) > forvar1207))));
                    end
                  else
                    begin
                      reg1237 <= ((^(~(reg1212 ?
                          forvar1230 : reg1240))) <= $signed((~&(^~reg1240))));
                    end
                  if (($unsigned(forvar1200[(1'h0):(1'h0)]) ?
                      reg1228 : (reg1218 ?
                          {$signed(reg1221)} : reg1203[(4'hc):(1'h1)])))
                    begin
                      reg1241 <= reg1215[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1241 <= ($signed(forvar1207) ?
                          $unsigned(reg1227) : ((8'haa) ?
                              {reg1208[(4'h9):(2'h3)]} : $unsigned((reg1203 ?
                                  reg1206 : reg1196))));
                      reg1242 <= ($unsigned($unsigned((reg1212 ?
                              reg1211 : reg1218))) ?
                          {{((8'hb8) + reg1218)}} : ((^reg1196) - (((8'h9d) * reg1232) ^ (forvar1225 ~^ (8'ha4)))));
                      reg1243 <= ({(^~forvar1207)} ^ forvar1236);
                    end
                  if ({(~&((forvar1216 ? forvar1235 : reg1231) ?
                          $signed(reg1223) : reg1234[(4'hc):(4'hb)]))})
                    begin
                      reg1244 <= forvar1211;
                      reg1245 <= ((!reg1206[(4'hb):(4'h9)]) ?
                          reg1219[(1'h1):(1'h0)] : (-$signed($unsigned(forvar1204))));
                      reg1246 <= $unsigned(((^~(reg1233 > (8'hb3))) + $signed((~&reg1236))));
                    end
                  else
                    begin
                      reg1244 <= $signed(($unsigned((reg1239 >= forvar1240)) ?
                          reg1203[(1'h0):(1'h0)] : ({reg1226} ?
                              (^reg1194) : reg1214[(1'h0):(1'h0)])));
                    end
                end
            end
          else
            begin
              for (forvar1224 = (1'h0); (forvar1224 < (1'h1)); forvar1224 = (forvar1224 + (1'h1)))
                begin
                  for (forvar1225 = (1'h0); (forvar1225 < (1'h1)); forvar1225 = (forvar1225 + (1'h1)))
                    begin
                      reg1226 <= $signed(reg1242[(3'h6):(3'h5)]);
                      reg1227 <= (~|{(~^reg1217[(4'he):(3'h6)])});
                      reg1228 <= (~($signed((!reg1200)) + ((|reg1208) ?
                          $signed(reg1219) : reg1229)));
                    end
                  for (forvar1229 = (1'h0); (forvar1229 < (1'h0)); forvar1229 = (forvar1229 + (1'h1)))
                    begin
                      reg1230 <= ((($signed(forvar1205) ?
                              (reg1202 >= wire1188) : reg1228) ^ ($unsigned(forvar1240) ^ reg1221)) ?
                          (|forvar1200) : {{$signed(forvar1204)}});
                      reg1231 <= $signed(forvar1216[(3'h7):(1'h1)]);
                      reg1232 <= forvar1236[(3'h5):(1'h1)];
                      reg1233 <= $signed((reg1238 <<< reg1234));
                    end
                end
              reg1234 <= ($unsigned(reg1211) != (wire1188 && $signed(reg1231)));
              if ($unsigned(reg1236))
                begin
                  if (((8'hb7) | (&((reg1232 ?
                      reg1228 : reg1235) == $unsigned(reg1243)))))
                    begin
                      reg1235 <= forvar1198;
                      reg1236 <= forvar1211;
                    end
                  else
                    begin
                      reg1235 <= ($unsigned($signed(((8'hab) ?
                              (8'ha0) : reg1236))) ?
                          reg1212 : (^~$signed((wire1192 ~^ (8'hae)))));
                      reg1236 <= $unsigned((reg1236 ^ {reg1210[(3'h4):(1'h0)]}));
                    end
                  for (forvar1237 = (1'h0); (forvar1237 < (2'h2)); forvar1237 = (forvar1237 + (1'h1)))
                    begin
                      reg1238 <= (|$signed(reg1214[(2'h3):(1'h1)]));
                      reg1239 <= (^~(|$signed((forvar1222 - reg1205))));
                      reg1240 <= $unsigned($unsigned($signed((forvar1235 - reg1212))));
                    end
                  reg1241 <= reg1197[(1'h0):(1'h0)];
                end
              else
                begin
                  for (forvar1235 = (1'h0); (forvar1235 < (1'h0)); forvar1235 = (forvar1235 + (1'h1)))
                    begin
                      reg1236 <= ($unsigned(((forvar1214 ?
                              reg1240 : forvar1225) ?
                          $unsigned((8'hb9)) : {forvar1205})) || forvar1204);
                      reg1237 <= reg1227;
                    end
                  if (reg1199[(3'h5):(3'h5)])
                    begin
                      reg1238 <= reg1227;
                      reg1239 <= (reg1233[(2'h3):(2'h2)] ?
                          (+((forvar1203 <= forvar1205) - $unsigned(reg1235))) : ((-forvar1222) ?
                              $signed($unsigned((8'ha4))) : reg1241[(3'h5):(3'h5)]));
                      reg1240 <= $unsigned(reg1234[(3'h5):(1'h0)]);
                      reg1241 <= (^~(-reg1245));
                    end
                  else
                    begin
                      reg1238 <= (($unsigned((8'ha7)) ?
                          reg1244 : reg1196) >> $unsigned(({reg1244} >> (reg1199 >= (8'had)))));
                      reg1239 <= (($unsigned($signed(reg1231)) > $signed($unsigned(forvar1240))) ?
                          $signed(forvar1230) : $unsigned((wire1192 - (reg1208 != reg1230))));
                    end
                  for (forvar1242 = (1'h0); (forvar1242 < (2'h2)); forvar1242 = (forvar1242 + (1'h1)))
                    begin
                      reg1243 <= (reg1214 + $signed($signed(reg1210[(4'h9):(4'h8)])));
                      reg1244 <= forvar1194;
                      reg1245 <= $signed(reg1223[(3'h5):(3'h4)]);
                    end
                end
            end
        end
    end
  assign wire1247 = wire1191[(3'h5):(2'h2)];
  assign wire1248 = (~&reg1237[(3'h6):(3'h5)]);
  assign wire1249 = ((8'hb9) ?
                        reg1231 : $signed(((reg1208 ? reg1237 : wire1191) ?
                            (&reg1231) : wire1248[(2'h3):(2'h3)])));
  assign wire1250 = (8'ha1);
  always
    @(posedge clk) begin
      if (($unsigned(wire1193[(4'ha):(3'h6)]) ?
          (($signed(reg1239) - (wire1190 < reg1194)) ?
              (-$signed(reg1220)) : reg1231) : ($unsigned(reg1221) ?
              $unsigned({reg1218}) : (|(8'h9e)))))
        begin
          if ((((+(reg1194 | reg1215)) ?
              ((+reg1243) ?
                  $unsigned(reg1194) : reg1228[(3'h5):(2'h2)]) : $unsigned($unsigned(reg1207))) ^~ $signed({(8'hb5)})))
            begin
              if (((~^reg1206) == {wire1189}))
                begin
                  for (forvar1251 = (1'h0); (forvar1251 < (2'h2)); forvar1251 = (forvar1251 + (1'h1)))
                    begin
                      reg1252 <= (+$signed(reg1242[(1'h0):(1'h0)]));
                      reg1253 <= $signed(($signed(reg1242) >= {((8'hb3) ?
                              reg1209 : wire1190)}));
                      reg1254 <= $unsigned((~^reg1211));
                    end
                  for (forvar1255 = (1'h0); (forvar1255 < (2'h3)); forvar1255 = (forvar1255 + (1'h1)))
                    begin
                      reg1256 <= $signed($signed(((reg1218 ?
                          reg1209 : reg1221) + (^~wire1248))));
                      reg1257 <= $unsigned(reg1206);
                      reg1258 <= reg1206;
                      reg1259 <= (^$signed(($unsigned(reg1246) && (^~wire1250))));
                    end
                  for (forvar1260 = (1'h0); (forvar1260 < (1'h0)); forvar1260 = (forvar1260 + (1'h1)))
                    begin
                      reg1261 <= (($signed($unsigned(reg1214)) <<< $signed(reg1257[(1'h1):(1'h1)])) ?
                          $signed(reg1202[(1'h1):(1'h0)]) : $unsigned(reg1230));
                    end
                end
              else
                begin
                  if (((~^{(8'ha7)}) > $signed($signed(reg1223[(3'h5):(1'h0)]))))
                    begin
                      reg1251 <= reg1254[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg1251 <= $signed($unsigned((~^reg1258)));
                    end
                  for (forvar1252 = (1'h0); (forvar1252 < (1'h1)); forvar1252 = (forvar1252 + (1'h1)))
                    begin
                      reg1253 <= reg1211[(3'h6):(2'h3)];
                      reg1254 <= reg1223[(1'h0):(1'h0)];
                    end
                  for (forvar1255 = (1'h0); (forvar1255 < (1'h1)); forvar1255 = (forvar1255 + (1'h1)))
                    begin
                      reg1256 <= $signed({reg1236[(1'h1):(1'h0)]});
                    end
                end
            end
          else
            begin
              reg1251 <= ((~^reg1258[(4'h9):(3'h6)]) ?
                  $signed(($signed(reg1213) == {reg1258})) : ($signed((reg1195 ?
                          (8'h9e) : reg1220)) ?
                      reg1244 : $signed($unsigned(reg1237))));
              for (forvar1252 = (1'h0); (forvar1252 < (1'h0)); forvar1252 = (forvar1252 + (1'h1)))
                begin
                  if ((($unsigned(reg1239) & (reg1206 ?
                      wire1190 : (reg1220 >> (8'haa)))) || reg1257[(1'h0):(1'h0)]))
                    begin
                      reg1253 <= $signed(reg1214[(1'h1):(1'h1)]);
                      reg1254 <= wire1190[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg1253 <= ($unsigned($unsigned($unsigned(reg1226))) ^~ ((reg1199[(1'h0):(1'h0)] < reg1200[(1'h1):(1'h0)]) || ($unsigned(reg1236) ?
                          $signed((8'ha8)) : (reg1212 * wire1193))));
                      reg1254 <= reg1244;
                    end
                end
            end
          if (reg1211[(2'h3):(2'h2)])
            begin
              for (forvar1262 = (1'h0); (forvar1262 < (1'h1)); forvar1262 = (forvar1262 + (1'h1)))
                begin
                  if (($signed(({reg1223} ?
                      (reg1244 & (8'hae)) : (wire1249 < (8'hb8)))) > forvar1262))
                    begin
                      reg1263 <= (^~(^{reg1235}));
                    end
                  else
                    begin
                      reg1263 <= (reg1212 ~^ $unsigned(reg1214[(3'h4):(1'h1)]));
                      reg1264 <= (((~^reg1226) != ($signed(reg1206) * ((8'ha9) <= reg1223))) >= wire1193[(4'hd):(3'h4)]);
                      reg1265 <= wire1250;
                      reg1266 <= reg1228[(1'h1):(1'h0)];
                    end
                  for (forvar1267 = (1'h0); (forvar1267 < (2'h3)); forvar1267 = (forvar1267 + (1'h1)))
                    begin
                      reg1268 <= (reg1257[(1'h1):(1'h1)] ?
                          {(&(8'had))} : $signed($signed(((8'haf) ^ reg1266))));
                      reg1269 <= (wire1189 ?
                          (~|(~$signed(reg1215))) : wire1188[(3'h4):(2'h2)]);
                      reg1270 <= reg1263;
                    end
                end
              if ((^reg1246))
                begin
                  for (forvar1271 = (1'h0); (forvar1271 < (2'h2)); forvar1271 = (forvar1271 + (1'h1)))
                    begin
                      reg1272 <= (~&reg1195[(3'h6):(1'h1)]);
                      reg1273 <= reg1212;
                      reg1274 <= {(~|(8'ha1))};
                      reg1275 <= (reg1228[(3'h4):(3'h4)] ~^ reg1195[(2'h2):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar1271 = (1'h0); (forvar1271 < (2'h2)); forvar1271 = (forvar1271 + (1'h1)))
                    begin
                      reg1272 <= (reg1203 != (8'ha1));
                      reg1273 <= (($signed(reg1252[(3'h7):(3'h4)]) ?
                          (reg1200 ?
                              ((8'hb2) ?
                                  reg1235 : reg1264) : $unsigned(reg1263)) : wire1190) != reg1223[(3'h4):(2'h2)]);
                      reg1274 <= wire1190;
                      reg1275 <= $signed((^~(-(reg1213 ? reg1274 : reg1203))));
                    end
                end
            end
          else
            begin
              reg1262 <= reg1215;
            end
        end
      else
        begin
          if (reg1198[(4'hb):(2'h2)])
            begin
              for (forvar1251 = (1'h0); (forvar1251 < (2'h2)); forvar1251 = (forvar1251 + (1'h1)))
                begin
                  for (forvar1252 = (1'h0); (forvar1252 < (2'h2)); forvar1252 = (forvar1252 + (1'h1)))
                    begin
                      reg1253 <= $signed({((reg1270 ?
                              reg1221 : reg1242) <<< $signed(reg1238))});
                    end
                  for (forvar1254 = (1'h0); (forvar1254 < (2'h3)); forvar1254 = (forvar1254 + (1'h1)))
                    begin
                      reg1255 <= {((~&$unsigned(reg1227)) < reg1220)};
                    end
                  for (forvar1256 = (1'h0); (forvar1256 < (1'h1)); forvar1256 = (forvar1256 + (1'h1)))
                    begin
                      reg1257 <= reg1220[(2'h3):(2'h2)];
                    end
                  for (forvar1258 = (1'h0); (forvar1258 < (1'h1)); forvar1258 = (forvar1258 + (1'h1)))
                    begin
                      reg1259 <= (((reg1229[(2'h2):(1'h0)] ?
                          reg1210 : (-(8'ha4))) <= $unsigned((!wire1192))) ^~ (reg1211 > $unsigned((8'ha1))));
                      reg1260 <= (((reg1219[(4'hb):(1'h0)] < (&reg1265)) ?
                              reg1196[(3'h5):(3'h4)] : reg1215) ?
                          $signed((8'ha9)) : $signed({(reg1201 >>> reg1197)}));
                    end
                end
              for (forvar1261 = (1'h0); (forvar1261 < (2'h2)); forvar1261 = (forvar1261 + (1'h1)))
                begin
                  for (forvar1262 = (1'h0); (forvar1262 < (2'h2)); forvar1262 = (forvar1262 + (1'h1)))
                    begin
                      reg1263 <= reg1243[(1'h1):(1'h1)];
                      reg1264 <= ({$unsigned((reg1239 ?
                              reg1211 : reg1266))} >> (~|reg1253[(3'h4):(1'h1)]));
                    end
                  for (forvar1265 = (1'h0); (forvar1265 < (1'h0)); forvar1265 = (forvar1265 + (1'h1)))
                    begin
                      reg1266 <= $signed(forvar1260);
                      reg1267 <= (|reg1197);
                      reg1268 <= forvar1261;
                    end
                  reg1269 <= wire1192[(2'h3):(2'h3)];
                end
              for (forvar1270 = (1'h0); (forvar1270 < (1'h0)); forvar1270 = (forvar1270 + (1'h1)))
                begin
                  for (forvar1271 = (1'h0); (forvar1271 < (1'h0)); forvar1271 = (forvar1271 + (1'h1)))
                    begin
                      reg1272 <= $signed(($unsigned((^reg1257)) - (^$unsigned(forvar1255))));
                      reg1273 <= ((8'hb6) ~^ $unsigned(reg1200));
                      reg1274 <= $signed($unsigned({{reg1217}}));
                    end
                  for (forvar1275 = (1'h0); (forvar1275 < (1'h0)); forvar1275 = (forvar1275 + (1'h1)))
                    begin
                      reg1276 <= reg1237;
                      reg1277 <= reg1235[(4'hc):(1'h0)];
                      reg1278 <= reg1259;
                      reg1279 <= $unsigned($unsigned((^(wire1247 ?
                          reg1277 : reg1243))));
                    end
                end
            end
          else
            begin
              for (forvar1251 = (1'h0); (forvar1251 < (1'h1)); forvar1251 = (forvar1251 + (1'h1)))
                begin
                  if ((~^reg1272))
                    begin
                      reg1252 <= (|($signed((reg1199 + reg1265)) ?
                          (^~{wire1250}) : ($signed(wire1192) ?
                              (~^reg1272) : $signed(forvar1260))));
                    end
                  else
                    begin
                      reg1252 <= $unsigned(wire1189);
                      reg1253 <= ((8'ha4) || reg1265);
                      reg1254 <= (~reg1251[(4'he):(3'h4)]);
                      reg1255 <= reg1254[(2'h2):(1'h0)];
                    end
                  if (reg1245)
                    begin
                      reg1256 <= $signed((wire1190 ?
                          forvar1252 : (^(reg1240 ? (8'ha2) : reg1240))));
                      reg1257 <= $signed($unsigned(forvar1255));
                    end
                  else
                    begin
                      reg1256 <= $signed((8'hb0));
                      reg1257 <= $signed({(^reg1237)});
                      reg1258 <= (~|(($signed(reg1220) ^ ((8'haf) ?
                              forvar1260 : reg1279)) ?
                          ($unsigned((8'hb1)) ?
                              wire1191[(1'h0):(1'h0)] : (reg1231 | reg1243)) : reg1195));
                    end
                  if (reg1228[(2'h2):(1'h1)])
                    begin
                      reg1259 <= (~$unsigned($unsigned(reg1266)));
                      reg1260 <= reg1219[(4'hb):(3'h6)];
                      reg1261 <= (~$unsigned($unsigned((reg1255 <<< reg1212))));
                    end
                  else
                    begin
                      reg1259 <= wire1193[(4'h9):(4'h9)];
                      reg1260 <= $unsigned((((reg1273 ?
                              (8'hae) : (8'hb9)) ^ reg1210) ?
                          (reg1270 < (~^forvar1252)) : $signed($unsigned(reg1210))));
                    end
                  if (((+($signed(wire1250) ?
                      $signed(reg1276) : $unsigned(reg1231))) == ({$unsigned((8'hb5))} ^~ $unsigned(forvar1265))))
                    begin
                      reg1262 <= $unsigned(({(&reg1215)} >= ((forvar1258 ?
                          forvar1262 : reg1207) > {(8'ha0)})));
                    end
                  else
                    begin
                      reg1262 <= ((reg1218[(4'hc):(4'h9)] <= reg1200[(3'h4):(2'h3)]) ?
                          $signed(((reg1267 + reg1226) ?
                              {reg1242} : reg1200)) : {reg1272});
                      reg1263 <= (~|((forvar1275[(4'ha):(2'h2)] ?
                              (^~forvar1271) : $signed(reg1226)) ?
                          reg1253 : {$signed(forvar1261)}));
                      reg1264 <= {$signed(wire1250[(2'h3):(1'h0)])};
                      reg1265 <= reg1256[(2'h3):(2'h3)];
                    end
                end
              for (forvar1266 = (1'h0); (forvar1266 < (2'h2)); forvar1266 = (forvar1266 + (1'h1)))
                begin
                  for (forvar1267 = (1'h0); (forvar1267 < (1'h0)); forvar1267 = (forvar1267 + (1'h1)))
                    begin
                      reg1268 <= (+(!reg1232[(4'ha):(3'h6)]));
                    end
                  if ($unsigned(({wire1247} - {(^~reg1257)})))
                    begin
                      reg1269 <= (-$signed($signed({reg1219})));
                    end
                  else
                    begin
                      reg1269 <= {reg1259[(1'h0):(1'h0)]};
                      reg1270 <= (($signed({reg1227}) ?
                              ($signed(reg1234) < (-reg1253)) : (~forvar1252)) ?
                          $signed((-$unsigned(reg1245))) : reg1273);
                      reg1271 <= $signed(wire1190[(1'h0):(1'h0)]);
                    end
                  for (forvar1272 = (1'h0); (forvar1272 < (2'h3)); forvar1272 = (forvar1272 + (1'h1)))
                    begin
                      reg1273 <= $unsigned(reg1265[(4'h8):(1'h1)]);
                      reg1274 <= {$unsigned($unsigned((reg1208 ?
                              reg1279 : reg1227)))};
                    end
                  reg1275 <= (forvar1270[(1'h1):(1'h0)] <<< (forvar1260[(3'h7):(3'h5)] << $signed(((8'ha2) != forvar1271))));
                end
            end
        end
      for (forvar1280 = (1'h0); (forvar1280 < (2'h3)); forvar1280 = (forvar1280 + (1'h1)))
        begin
          reg1281 <= (reg1233 ~^ reg1258);
          if ($unsigned($signed((^~((8'hb5) ? (8'h9c) : reg1209)))))
            begin
              reg1282 <= $signed((reg1253[(2'h2):(1'h0)] ^ {reg1238}));
              reg1283 <= $unsigned((((reg1262 >= forvar1255) || (~|reg1281)) ?
                  reg1230[(2'h2):(1'h0)] : wire1189));
            end
          else
            begin
              reg1282 <= reg1233[(2'h2):(1'h1)];
              for (forvar1283 = (1'h0); (forvar1283 < (1'h0)); forvar1283 = (forvar1283 + (1'h1)))
                begin
                  reg1284 <= reg1236[(3'h4):(3'h4)];
                  for (forvar1285 = (1'h0); (forvar1285 < (1'h1)); forvar1285 = (forvar1285 + (1'h1)))
                    begin
                      reg1286 <= wire1190;
                      reg1287 <= $unsigned(reg1235);
                    end
                end
            end
        end
      for (forvar1288 = (1'h0); (forvar1288 < (2'h2)); forvar1288 = (forvar1288 + (1'h1)))
        begin
          if (reg1240)
            begin
              if (forvar1252[(2'h2):(2'h2)])
                begin
                  if (((~((~^reg1245) | forvar1252)) < reg1262[(3'h6):(3'h6)]))
                    begin
                      reg1289 <= $unsigned((!forvar1270));
                    end
                  else
                    begin
                      reg1289 <= ($signed(reg1278[(1'h1):(1'h0)]) | $signed($signed((^(8'hb0)))));
                      reg1290 <= wire1250;
                    end
                  if (forvar1288)
                    begin
                      reg1291 <= $unsigned($signed($unsigned(((8'hac) << reg1246))));
                      reg1292 <= {({reg1209[(1'h1):(1'h0)]} <= (&{reg1210}))};
                    end
                  else
                    begin
                      reg1291 <= ((~^{wire1190[(3'h5):(1'h1)]}) ?
                          $unsigned((8'hb8)) : ((~reg1203) & reg1217));
                      reg1292 <= ((^~($unsigned((8'had)) ?
                          {wire1188} : (+forvar1255))) ^~ $signed(((-(8'h9d)) <<< $signed(reg1198))));
                      reg1293 <= reg1265;
                      reg1294 <= reg1245[(2'h2):(2'h2)];
                    end
                  for (forvar1295 = (1'h0); (forvar1295 < (2'h2)); forvar1295 = (forvar1295 + (1'h1)))
                    begin
                      reg1296 <= {{{(reg1232 ? forvar1267 : (8'had))}}};
                      reg1297 <= reg1214;
                      reg1298 <= $unsigned((+(reg1290 << (~^reg1278))));
                      reg1299 <= $unsigned({$unsigned(((8'ha0) ?
                              reg1264 : reg1263))});
                    end
                  for (forvar1300 = (1'h0); (forvar1300 < (1'h0)); forvar1300 = (forvar1300 + (1'h1)))
                    begin
                      reg1301 <= reg1266;
                      reg1302 <= (reg1274 == reg1284[(3'h6):(2'h2)]);
                      reg1303 <= $unsigned(reg1215);
                    end
                end
              else
                begin
                  if ($signed(reg1215))
                    begin
                      reg1289 <= $unsigned(($unsigned({(8'hb2)}) << (+reg1294)));
                      reg1290 <= {(reg1297 | reg1230[(3'h4):(1'h0)])};
                    end
                  else
                    begin
                      reg1289 <= (reg1198 | (reg1272 ?
                          {{reg1289}} : $signed(reg1201[(3'h6):(1'h0)])));
                      reg1290 <= ({reg1268[(1'h0):(1'h0)]} ?
                          reg1292 : (!{(forvar1300 <= reg1207)}));
                      reg1291 <= (^~reg1198[(4'hd):(3'h4)]);
                    end
                end
              if (reg1208)
                begin
                  for (forvar1304 = (1'h0); (forvar1304 < (2'h3)); forvar1304 = (forvar1304 + (1'h1)))
                    begin
                      reg1305 <= reg1258;
                      reg1306 <= reg1296;
                      reg1307 <= (&(reg1273 > $unsigned(((8'ha0) >>> reg1281))));
                    end
                  if ((8'haa))
                    begin
                      reg1308 <= (($signed((reg1256 <<< (8'ha9))) ?
                              {(reg1303 <<< reg1273)} : ($signed(reg1242) ?
                                  $unsigned((8'hb9)) : $signed(reg1230))) ?
                          $unsigned(reg1263[(4'h8):(2'h2)]) : {$unsigned((forvar1300 <<< reg1297))});
                      reg1309 <= (~^(~(reg1235 > $signed(reg1277))));
                      reg1310 <= reg1195;
                      reg1311 <= ($unsigned($unsigned($unsigned(reg1268))) & ($unsigned((reg1209 ?
                          reg1283 : reg1200)) >= reg1212[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg1308 <= (($signed(((8'h9f) != reg1307)) ?
                              reg1302 : reg1199) ?
                          $unsigned(reg1258) : {reg1269});
                    end
                  reg1312 <= (^$unsigned(((reg1278 != reg1215) | $unsigned(reg1278))));
                end
              else
                begin
                  if (({$signed((reg1220 ? reg1211 : reg1239))} ?
                      (^~reg1220) : $signed(((^~wire1250) <= (wire1190 ?
                          forvar1262 : (8'ha3))))))
                    begin
                      reg1304 <= wire1189[(1'h0):(1'h0)];
                      reg1305 <= ((8'hb7) == $signed((8'ha5)));
                      reg1306 <= $unsigned(forvar1256[(4'ha):(4'h9)]);
                    end
                  else
                    begin
                      reg1304 <= $signed((reg1277 ?
                          $unsigned((reg1197 && reg1270)) : (~&(forvar1285 ?
                              reg1241 : reg1212))));
                    end
                  for (forvar1307 = (1'h0); (forvar1307 < (1'h1)); forvar1307 = (forvar1307 + (1'h1)))
                    begin
                      reg1308 <= $signed((reg1233 ?
                          (^reg1261[(1'h0):(1'h0)]) : (&((8'ha3) || forvar1265))));
                    end
                end
              if ((|(^~{$signed(reg1196)})))
                begin
                  for (forvar1313 = (1'h0); (forvar1313 < (2'h2)); forvar1313 = (forvar1313 + (1'h1)))
                    begin
                      reg1314 <= reg1198[(2'h3):(2'h2)];
                      reg1315 <= {((((8'hab) | reg1263) ?
                                  (&wire1190) : {reg1204}) ?
                              ($unsigned(wire1248) ?
                                  forvar1260[(4'hc):(4'h8)] : {reg1236}) : forvar1307)};
                    end
                  for (forvar1316 = (1'h0); (forvar1316 < (2'h3)); forvar1316 = (forvar1316 + (1'h1)))
                    begin
                      reg1317 <= forvar1262[(3'h4):(3'h4)];
                      reg1318 <= (reg1200 <= (!(~&(wire1192 ?
                          (8'hb3) : reg1204))));
                      reg1319 <= ((((reg1277 ?
                          reg1258 : reg1230) & $signed(forvar1256)) || ($signed((8'hb7)) << $unsigned(reg1210))) ^ wire1189[(4'ha):(4'ha)]);
                      reg1320 <= $unsigned((^~(-$signed(reg1262))));
                    end
                end
              else
                begin
                  if (((reg1312[(1'h1):(1'h0)] ?
                          reg1284[(3'h5):(2'h3)] : ($signed(reg1211) >> (+reg1194))) ?
                      {$unsigned($unsigned(reg1307))} : {($unsigned(forvar1256) <= reg1236)}))
                    begin
                      reg1313 <= $signed(forvar1267);
                      reg1314 <= reg1205;
                    end
                  else
                    begin
                      reg1313 <= reg1242[(2'h2):(1'h0)];
                      reg1314 <= $unsigned($unsigned(reg1254[(2'h2):(2'h2)]));
                      reg1315 <= (forvar1254 ?
                          (+{$signed(reg1200)}) : reg1216[(1'h1):(1'h0)]);
                    end
                end
              if ($unsigned((($signed((8'ha9)) ?
                  reg1283 : ((8'hb9) == forvar1280)) >= ($signed(reg1221) - $signed(reg1258)))))
                begin
                  if (({$unsigned($signed((8'h9d)))} == (|(^(~&reg1232)))))
                    begin
                      reg1321 <= (reg1308 ^~ forvar1285[(3'h5):(2'h3)]);
                      reg1322 <= (reg1319 << (!(~&(reg1214 || reg1206))));
                      reg1323 <= ({($signed(reg1231) ~^ {reg1220})} == $signed($unsigned($signed(forvar1272))));
                      reg1324 <= (reg1261[(3'h6):(2'h2)] ?
                          forvar1316 : (+(+reg1221[(2'h3):(2'h2)])));
                    end
                  else
                    begin
                      reg1321 <= (reg1246 ^ (~^$unsigned($signed((8'hac)))));
                      reg1322 <= $signed($signed($signed((reg1195 ~^ forvar1280))));
                      reg1323 <= $unsigned(((8'ha5) ?
                          (reg1261[(4'hf):(4'he)] >>> $unsigned(reg1293)) : reg1230[(3'h5):(3'h4)]));
                      reg1324 <= (-(-{$signed((8'hb5))}));
                    end
                  for (forvar1325 = (1'h0); (forvar1325 < (2'h3)); forvar1325 = (forvar1325 + (1'h1)))
                    begin
                      reg1326 <= ($signed(reg1313) >= ((+reg1284[(2'h2):(1'h0)]) ?
                          reg1312 : reg1278));
                    end
                  for (forvar1327 = (1'h0); (forvar1327 < (1'h1)); forvar1327 = (forvar1327 + (1'h1)))
                    begin
                      reg1328 <= wire1188;
                    end
                  for (forvar1329 = (1'h0); (forvar1329 < (2'h3)); forvar1329 = (forvar1329 + (1'h1)))
                    begin
                      reg1330 <= reg1307;
                      reg1331 <= ((reg1261 ?
                          (reg1293[(1'h1):(1'h0)] ^~ reg1264) : (reg1273[(3'h7):(1'h0)] & (8'hb0))) <<< ({$unsigned(reg1198)} ?
                          $signed(reg1260[(4'hb):(1'h1)]) : {(reg1258 ?
                                  reg1291 : wire1249)}));
                      reg1332 <= ($signed((~$unsigned(reg1221))) ?
                          $unsigned($unsigned($unsigned((8'hb6)))) : (!reg1205));
                      reg1333 <= reg1276[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  reg1321 <= forvar1275;
                end
            end
          else
            begin
              if (($unsigned($signed(reg1310)) ?
                  $unsigned(((!reg1245) >>> (-reg1270))) : ((~&wire1193) ?
                      {$unsigned(reg1241)} : (-(reg1208 ? reg1305 : reg1312)))))
                begin
                  reg1289 <= (($signed((+(8'hb8))) ?
                      (wire1191[(4'ha):(4'ha)] <= $signed(forvar1270)) : ($unsigned((8'hb3)) ~^ reg1269)) < ((!$unsigned(reg1261)) != $signed((reg1211 ?
                      forvar1261 : (8'hb4)))));
                  reg1290 <= (~$unsigned($signed(((8'ha5) ?
                      reg1194 : reg1270))));
                  if ($unsigned(($unsigned(forvar1266[(2'h3):(2'h2)]) ?
                      ((-reg1312) ?
                          (reg1241 || (8'ha7)) : reg1313[(4'h8):(3'h6)]) : ((^reg1286) + $unsigned(reg1218)))))
                    begin
                      reg1291 <= $unsigned((($unsigned(reg1278) ^ {reg1231}) ?
                          ((forvar1272 & reg1314) << reg1313[(1'h0):(1'h0)]) : (8'h9c)));
                    end
                  else
                    begin
                      reg1291 <= reg1287[(4'he):(3'h6)];
                    end
                  if ({reg1263[(4'he):(3'h7)]})
                    begin
                      reg1292 <= reg1292;
                    end
                  else
                    begin
                      reg1292 <= ($signed(reg1196[(2'h3):(2'h3)]) != $unsigned(reg1245));
                      reg1293 <= (reg1204 ?
                          $unsigned((~(forvar1252 ?
                              (8'ha7) : reg1311))) : ($signed({reg1274}) != wire1188[(1'h1):(1'h0)]));
                      reg1294 <= (8'hb9);
                      reg1295 <= $unsigned(((~((8'hac) ?
                          forvar1285 : reg1230)) && $signed(reg1313)));
                    end
                end
              else
                begin
                  if ((reg1270 >= forvar1272))
                    begin
                      reg1289 <= {wire1191[(4'hf):(2'h3)]};
                    end
                  else
                    begin
                      reg1289 <= reg1304;
                      reg1290 <= $signed((reg1332 > forvar1313));
                    end
                end
              if ((({(-reg1263)} ?
                      $signed((reg1211 | reg1298)) : reg1217[(4'hd):(3'h6)]) ?
                  $signed(($signed(reg1221) ?
                      (reg1270 ? (8'hb1) : reg1217) : reg1219)) : reg1270))
                begin
                  for (forvar1296 = (1'h0); (forvar1296 < (2'h3)); forvar1296 = (forvar1296 + (1'h1)))
                    begin
                      reg1297 <= $unsigned((8'hb9));
                      reg1298 <= (8'hb2);
                      reg1299 <= (reg1272[(2'h3):(2'h2)] >> (~&reg1299[(3'h4):(1'h0)]));
                    end
                  reg1300 <= reg1270;
                  for (forvar1301 = (1'h0); (forvar1301 < (1'h0)); forvar1301 = (forvar1301 + (1'h1)))
                    begin
                      reg1302 <= ((!$signed((8'hb3))) ? reg1194 : forvar1313);
                      reg1303 <= $unsigned($signed(reg1262[(3'h7):(3'h7)]));
                      reg1304 <= (~|(((reg1298 ?
                          reg1195 : reg1221) == $signed(reg1324)) >>> reg1238[(1'h1):(1'h0)]));
                    end
                  reg1305 <= $unsigned(reg1293);
                end
              else
                begin
                  reg1296 <= ((forvar1266 >= $signed($signed((8'hb5)))) ?
                      $signed(($unsigned(reg1197) >> reg1236[(3'h5):(3'h5)])) : reg1259);
                  if ({($unsigned($signed(reg1277)) ?
                          (&reg1198) : (^((8'hb1) >>> reg1317)))})
                    begin
                      reg1297 <= reg1333;
                      reg1298 <= $unsigned((~|$signed($signed(reg1278))));
                      reg1299 <= (^~(~^(~|{reg1302})));
                    end
                  else
                    begin
                      reg1297 <= (forvar1262[(1'h0):(1'h0)] ?
                          $signed(reg1296[(1'h1):(1'h1)]) : (($signed(reg1307) ?
                              reg1220[(2'h2):(1'h1)] : (reg1328 ?
                                  (8'hab) : reg1196)) - {(reg1307 != (8'hae))}));
                      reg1298 <= reg1218[(4'h8):(4'h8)];
                    end
                  reg1300 <= ((^$signed(reg1194[(1'h0):(1'h0)])) << forvar1295);
                end
              for (forvar1306 = (1'h0); (forvar1306 < (2'h2)); forvar1306 = (forvar1306 + (1'h1)))
                begin
                  reg1307 <= $signed({(-$unsigned(reg1294))});
                  for (forvar1308 = (1'h0); (forvar1308 < (1'h0)); forvar1308 = (forvar1308 + (1'h1)))
                    begin
                      reg1309 <= reg1333[(1'h1):(1'h1)];
                      reg1310 <= reg1300[(1'h0):(1'h0)];
                    end
                  reg1311 <= (~&((reg1301 ?
                      (~|reg1243) : $unsigned(reg1231)) * reg1242[(1'h0):(1'h0)]));
                end
              for (forvar1312 = (1'h0); (forvar1312 < (1'h0)); forvar1312 = (forvar1312 + (1'h1)))
                begin
                  if ({reg1201[(2'h3):(1'h1)]})
                    begin
                      reg1313 <= (reg1269 ?
                          $unsigned($signed((~^(8'h9d)))) : reg1310);
                      reg1314 <= $unsigned(reg1322[(3'h5):(3'h5)]);
                    end
                  else
                    begin
                      reg1313 <= ($signed((((8'had) | reg1195) ?
                          (wire1249 ?
                              reg1226 : reg1275) : $unsigned(reg1258))) && reg1310[(2'h3):(1'h1)]);
                    end
                  for (forvar1315 = (1'h0); (forvar1315 < (1'h1)); forvar1315 = (forvar1315 + (1'h1)))
                    begin
                      reg1316 <= (({(reg1283 ?
                              reg1279 : forvar1265)} ^ $unsigned(wire1189[(3'h4):(2'h2)])) == reg1297[(4'h9):(4'h9)]);
                      reg1317 <= {{($signed(reg1261) ?
                                  (forvar1267 < wire1190) : (reg1256 <<< reg1333))}};
                      reg1318 <= $unsigned(((^~(~|reg1313)) ?
                          (reg1315[(4'ha):(3'h5)] ?
                              $unsigned(reg1214) : (^reg1235)) : (~&$signed(forvar1254))));
                      reg1319 <= {(|{$signed((8'haa))})};
                    end
                end
            end
          if (reg1260[(3'h4):(1'h0)])
            begin
              for (forvar1334 = (1'h0); (forvar1334 < (1'h1)); forvar1334 = (forvar1334 + (1'h1)))
                begin
                  for (forvar1335 = (1'h0); (forvar1335 < (2'h2)); forvar1335 = (forvar1335 + (1'h1)))
                    begin
                      reg1336 <= ((($unsigned(reg1319) ?
                          (reg1295 >>> (8'haf)) : (|reg1210)) > (!$signed(reg1313))) < (({reg1245} ~^ (&forvar1254)) ~^ (8'ha8)));
                      reg1337 <= ((reg1336[(3'h5):(3'h5)] ?
                          (reg1196[(1'h1):(1'h0)] >> wire1189) : wire1191[(4'he):(3'h5)]) == (($unsigned(forvar1325) == (wire1189 ?
                              reg1279 : (8'ha3))) ?
                          ($signed(reg1244) ?
                              $unsigned(reg1330) : (forvar1335 ?
                                  reg1235 : reg1232)) : forvar1329));
                      reg1338 <= (({reg1323[(2'h3):(1'h1)]} - reg1260[(2'h2):(1'h0)]) ?
                          ($signed($signed(reg1229)) << $unsigned((reg1203 ?
                              (8'hab) : forvar1308))) : {(forvar1267[(1'h0):(1'h0)] ?
                                  reg1333 : $unsigned(reg1245))});
                    end
                  if (reg1223)
                    begin
                      reg1339 <= (|(reg1326 ?
                          $unsigned(reg1331[(3'h6):(2'h3)]) : (+wire1188[(2'h2):(1'h0)])));
                      reg1340 <= (+$signed(reg1229));
                      reg1341 <= forvar1288[(4'h9):(2'h3)];
                      reg1342 <= forvar1272;
                    end
                  else
                    begin
                      reg1339 <= {$signed(forvar1283[(4'h8):(1'h0)])};
                    end
                  for (forvar1343 = (1'h0); (forvar1343 < (2'h2)); forvar1343 = (forvar1343 + (1'h1)))
                    begin
                      reg1344 <= reg1270[(1'h0):(1'h0)];
                      reg1345 <= $unsigned((reg1307[(3'h4):(2'h2)] ?
                          (~&reg1294[(2'h2):(1'h1)]) : (((8'ha6) ?
                                  (8'hb3) : reg1319) ?
                              $unsigned(reg1338) : reg1281[(2'h2):(1'h1)])));
                    end
                  for (forvar1346 = (1'h0); (forvar1346 < (2'h3)); forvar1346 = (forvar1346 + (1'h1)))
                    begin
                      reg1347 <= {(8'hac)};
                      reg1348 <= ((+{forvar1295[(3'h6):(3'h4)]}) * {((^reg1230) ?
                              $signed(reg1239) : (reg1239 ?
                                  reg1197 : reg1196))});
                      reg1349 <= (($signed((~(8'had))) ?
                              reg1283 : (-(reg1262 - (8'ha3)))) ?
                          $unsigned((~|reg1306[(3'h5):(2'h3)])) : ((|(~^wire1247)) ?
                              ({forvar1270} ?
                                  $unsigned(reg1254) : $unsigned(reg1292)) : $signed((+(8'hab)))));
                    end
                end
              for (forvar1350 = (1'h0); (forvar1350 < (1'h1)); forvar1350 = (forvar1350 + (1'h1)))
                begin
                  for (forvar1351 = (1'h0); (forvar1351 < (1'h0)); forvar1351 = (forvar1351 + (1'h1)))
                    begin
                      reg1352 <= wire1193;
                      reg1353 <= reg1274;
                    end
                  for (forvar1354 = (1'h0); (forvar1354 < (1'h0)); forvar1354 = (forvar1354 + (1'h1)))
                    begin
                      reg1355 <= $unsigned(forvar1325[(1'h1):(1'h0)]);
                      reg1356 <= (reg1202 ?
                          forvar1304[(4'h9):(1'h1)] : (forvar1267 >> forvar1296[(3'h6):(3'h5)]));
                      reg1357 <= $unsigned((8'hb3));
                      reg1358 <= (reg1194[(3'h6):(1'h1)] ?
                          $signed(reg1274[(4'hc):(3'h7)]) : reg1352[(1'h0):(1'h0)]);
                    end
                end
            end
          else
            begin
              if (wire1192[(1'h0):(1'h0)])
                begin
                  if (reg1293[(1'h1):(1'h1)])
                    begin
                      reg1334 <= $signed($unsigned((reg1231[(3'h6):(1'h1)] != $unsigned((8'ha5)))));
                    end
                  else
                    begin
                      reg1334 <= $unsigned(reg1219[(4'hb):(3'h6)]);
                      reg1335 <= {(reg1292 ?
                              (reg1302[(4'h8):(2'h3)] ?
                                  $unsigned(forvar1313) : (reg1322 ?
                                      reg1232 : reg1267)) : $signed((~&reg1251)))};
                      reg1336 <= (~(reg1287[(4'h9):(3'h6)] || (~|reg1306[(2'h2):(1'h1)])));
                    end
                  if (((!(^(forvar1254 == reg1256))) ?
                      (((~&reg1195) ? reg1276[(1'h1):(1'h0)] : (+(8'hb5))) ?
                          $unsigned(forvar1350) : reg1348[(4'hc):(3'h4)]) : wire1193))
                    begin
                      reg1337 <= $unsigned({forvar1334[(3'h5):(1'h0)]});
                      reg1338 <= forvar1327;
                      reg1339 <= $signed(reg1243[(2'h3):(2'h3)]);
                      reg1340 <= ({(^$signed(reg1214))} <<< (+$signed($unsigned(reg1260))));
                    end
                  else
                    begin
                      reg1337 <= forvar1260[(4'hd):(1'h0)];
                      reg1338 <= reg1219;
                    end
                  if (reg1219[(4'ha):(4'h9)])
                    begin
                      reg1341 <= forvar1334[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg1341 <= $unsigned(reg1276[(1'h1):(1'h1)]);
                      reg1342 <= {$signed({(8'ha0)})};
                      reg1343 <= forvar1285;
                      reg1344 <= $signed((((reg1315 ? reg1238 : forvar1283) ?
                          (reg1284 ?
                              forvar1312 : reg1254) : $signed(reg1254)) >> {(reg1208 | reg1337)}));
                    end
                  for (forvar1345 = (1'h0); (forvar1345 < (2'h3)); forvar1345 = (forvar1345 + (1'h1)))
                    begin
                      reg1346 <= ($signed((8'hb5)) ?
                          $signed(({reg1268} ?
                              $unsigned(reg1304) : (^~reg1344))) : $unsigned(((wire1250 == reg1349) ~^ reg1218[(4'h8):(1'h1)])));
                      reg1347 <= reg1199[(3'h7):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar1334 = (1'h0); (forvar1334 < (1'h1)); forvar1334 = (forvar1334 + (1'h1)))
                    begin
                      reg1335 <= (8'hb3);
                      reg1336 <= ({{(reg1267 ? (8'hb7) : reg1348)}} ?
                          ($signed((-reg1263)) ?
                              ((-reg1273) ?
                                  (-reg1204) : (~(8'ha9))) : reg1199) : (reg1357[(3'h6):(2'h3)] ?
                              reg1244 : ($signed(reg1291) < $signed(reg1259))));
                      reg1337 <= ((~^($signed(reg1258) ?
                          (reg1239 >= forvar1295) : $unsigned(forvar1325))) & (forvar1304[(3'h7):(3'h7)] ^~ ((8'ha7) ?
                          (~reg1206) : (reg1206 & forvar1285))));
                    end
                  if ($signed((($signed(reg1245) ?
                          (|reg1338) : (wire1192 && reg1218)) ?
                      (reg1299 ^ $unsigned(forvar1345)) : forvar1267)))
                    begin
                      reg1338 <= $signed((^$signed($signed(reg1287))));
                      reg1339 <= (8'hba);
                      reg1340 <= $signed(forvar1270[(3'h4):(1'h0)]);
                      reg1341 <= $unsigned(forvar1272);
                    end
                  else
                    begin
                      reg1338 <= reg1357;
                    end
                  if (((forvar1254 ?
                          $unsigned(reg1200[(4'h8):(1'h0)]) : $unsigned((reg1312 + reg1317))) ?
                      forvar1301[(3'h4):(2'h3)] : reg1264[(4'hd):(4'hc)]))
                    begin
                      reg1342 <= $unsigned(({reg1315} != reg1267[(4'h8):(2'h3)]));
                    end
                  else
                    begin
                      reg1342 <= reg1237[(1'h1):(1'h1)];
                    end
                  for (forvar1343 = (1'h0); (forvar1343 < (2'h2)); forvar1343 = (forvar1343 + (1'h1)))
                    begin
                      reg1344 <= (($signed($signed(forvar1262)) ?
                          (~&(reg1212 ?
                              (8'ha6) : reg1343)) : reg1228[(3'h5):(3'h4)]) == ($signed((reg1352 ?
                          reg1202 : forvar1312)) ^~ (!{reg1215})));
                    end
                end
              reg1348 <= ((((|reg1207) ?
                      reg1233[(4'h8):(2'h2)] : ((8'ha0) ?
                          (8'ha4) : reg1240)) >>> ((8'h9d) ?
                      reg1233[(3'h6):(3'h5)] : $unsigned(reg1292))) ?
                  reg1213 : ({reg1265[(4'h9):(4'h8)]} ?
                      reg1278 : ((forvar1266 ? forvar1308 : reg1272) ?
                          (forvar1343 <= reg1311) : (8'ha3))));
            end
        end
      if (forvar1255)
        begin
          if (wire1192)
            begin
              if (($signed((reg1206[(1'h0):(1'h0)] && $unsigned(reg1341))) * ($signed({reg1261}) ?
                  (+$signed((8'ha7))) : (forvar1343 || (~&forvar1283)))))
                begin
                  if ((($unsigned((wire1193 > reg1322)) ?
                          ($signed((8'hb1)) ?
                              $unsigned(reg1326) : ((8'ha1) == (8'ha2))) : ((reg1347 <<< wire1190) ^~ forvar1261[(3'h6):(3'h6)])) ?
                      $signed(reg1241) : forvar1262[(2'h3):(1'h1)]))
                    begin
                      reg1359 <= $unsigned(reg1330[(1'h1):(1'h1)]);
                      reg1360 <= $signed((forvar1304 ?
                          $unsigned(reg1324[(3'h4):(3'h4)]) : ((reg1335 >= forvar1258) ?
                              $unsigned(reg1356) : (!reg1206))));
                      reg1361 <= $unsigned({({reg1352} ?
                              $signed(forvar1304) : reg1236)});
                    end
                  else
                    begin
                      reg1359 <= (^$signed(((reg1221 ?
                          reg1296 : (8'h9f)) != {reg1216})));
                    end
                end
              else
                begin
                  reg1359 <= ($signed(($signed(reg1234) <<< (8'h9f))) ?
                      ((reg1233 >>> (~&reg1360)) > reg1360) : (reg1226 ?
                          $unsigned(forvar1296) : $unsigned((reg1214 ~^ forvar1288))));
                  if (wire1190)
                    begin
                      reg1360 <= wire1247;
                      reg1361 <= $signed(reg1251);
                      reg1362 <= reg1353[(4'h9):(3'h6)];
                    end
                  else
                    begin
                      reg1360 <= $unsigned($signed($unsigned($signed(reg1273))));
                      reg1361 <= forvar1295[(1'h0):(1'h0)];
                      reg1362 <= $unsigned((+$unsigned((reg1287 ?
                          reg1197 : forvar1261))));
                    end
                end
            end
          else
            begin
              if ((!$unsigned(reg1306)))
                begin
                  for (forvar1359 = (1'h0); (forvar1359 < (1'h1)); forvar1359 = (forvar1359 + (1'h1)))
                    begin
                      reg1360 <= reg1194;
                      reg1361 <= (reg1287 ?
                          (($unsigned((8'ha1)) + $unsigned(reg1321)) - {(forvar1301 < forvar1256)}) : ($signed((reg1320 && reg1213)) ^ {$signed(forvar1300)}));
                      reg1362 <= $unsigned({(^~wire1189[(1'h0):(1'h0)])});
                      reg1363 <= ((&(8'h9d)) & {(!$unsigned(reg1195))});
                    end
                  for (forvar1364 = (1'h0); (forvar1364 < (2'h3)); forvar1364 = (forvar1364 + (1'h1)))
                    begin
                      reg1365 <= wire1188;
                    end
                  if (forvar1335[(3'h4):(1'h1)])
                    begin
                      reg1366 <= (&{(~^{reg1275})});
                      reg1367 <= (~&$signed($signed((forvar1261 > forvar1258))));
                      reg1368 <= $signed(reg1304[(3'h7):(3'h6)]);
                    end
                  else
                    begin
                      reg1366 <= (~((forvar1329[(3'h6):(3'h6)] ?
                          $unsigned(reg1301) : reg1289) | ((reg1256 ~^ (8'h9d)) << forvar1256[(4'h8):(4'h8)])));
                      reg1367 <= (wire1192 > $unsigned(reg1310));
                      reg1368 <= (!(8'hb7));
                    end
                  reg1369 <= $unsigned($signed($unsigned($unsigned((8'ha2)))));
                end
              else
                begin
                  for (forvar1359 = (1'h0); (forvar1359 < (1'h0)); forvar1359 = (forvar1359 + (1'h1)))
                    begin
                      reg1360 <= $unsigned($unsigned(({reg1236} ?
                          ((8'ha5) ? forvar1346 : forvar1325) : (&reg1331))));
                      reg1361 <= reg1258;
                      reg1362 <= (reg1335 ^~ $signed(forvar1266[(1'h1):(1'h1)]));
                    end
                  for (forvar1363 = (1'h0); (forvar1363 < (2'h2)); forvar1363 = (forvar1363 + (1'h1)))
                    begin
                      reg1364 <= ((reg1292 << reg1305) > $unsigned(reg1202));
                      reg1365 <= $unsigned((^reg1263));
                      reg1366 <= (~^(&forvar1251));
                      reg1367 <= $signed(reg1301[(4'h8):(3'h5)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar1359 = (1'h0); (forvar1359 < (1'h0)); forvar1359 = (forvar1359 + (1'h1)))
            begin
              for (forvar1360 = (1'h0); (forvar1360 < (1'h0)); forvar1360 = (forvar1360 + (1'h1)))
                begin
                  reg1361 <= (reg1197 ?
                      ((((8'ha5) ? reg1322 : (8'ha2)) != ((8'haf) ?
                          wire1192 : reg1287)) >>> $signed(reg1358[(3'h4):(1'h0)])) : (!((reg1342 <<< forvar1262) ?
                          $unsigned(reg1308) : forvar1254)));
                  if ((-forvar1304[(4'h9):(3'h6)]))
                    begin
                      reg1362 <= (^{(reg1236 << (reg1241 ?
                              reg1296 : (8'hb6)))});
                    end
                  else
                    begin
                      reg1362 <= reg1303;
                      reg1363 <= reg1289;
                    end
                  if ($signed(wire1247))
                    begin
                      reg1364 <= {$signed(($unsigned(reg1306) ?
                              $signed(reg1221) : reg1340))};
                      reg1365 <= $signed(forvar1360);
                      reg1366 <= (wire1188 >>> (^~reg1305));
                      reg1367 <= $unsigned($unsigned(reg1367));
                    end
                  else
                    begin
                      reg1364 <= {{$unsigned($unsigned(wire1248))}};
                      reg1365 <= forvar1300;
                      reg1366 <= $signed($unsigned(($signed(reg1299) ?
                          {reg1312} : $signed(reg1245))));
                      reg1367 <= {reg1254};
                    end
                end
            end
          if ({$signed((reg1204[(2'h3):(2'h3)] >> {reg1253}))})
            begin
              reg1368 <= reg1275;
              reg1369 <= (((forvar1308 ?
                      reg1246[(2'h3):(1'h1)] : reg1272[(3'h4):(3'h4)]) ?
                  ((reg1316 ?
                      (8'hb5) : forvar1288) <<< reg1330[(2'h3):(1'h0)]) : forvar1265[(3'h6):(1'h0)]) && (8'hb2));
            end
          else
            begin
              reg1368 <= forvar1345[(3'h6):(3'h6)];
            end
        end
    end
  assign wire1370 = (reg1261 == reg1322[(2'h3):(2'h3)]);
  assign wire1371 = $signed(($signed(wire1191[(4'h9):(1'h1)]) ?
                        (~|$unsigned(reg1268)) : (!((8'ha0) ?
                            (8'hb6) : reg1322))));
  assign wire1372 = reg1321;
endmodule