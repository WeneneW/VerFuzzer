(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'hd7e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire0;
  input wire signed [(4'hf):(1'h0)] wire1;
  input wire signed [(4'hc):(1'h0)] wire2;
  input wire [(4'hd):(1'h0)] wire3;
  input wire [(2'h2):(1'h0)] wire4;
  wire signed [(5'h10):(1'h0)] wire418;
  wire signed [(4'hc):(1'h0)] wire417;
  wire signed [(3'h6):(1'h0)] wire416;
  wire signed [(4'h9):(1'h0)] wire415;
  wire signed [(4'hb):(1'h0)] wire414;
  wire signed [(5'h10):(1'h0)] wire5;
  wire [(3'h6):(1'h0)] wire239;
  wire signed [(2'h2):(1'h0)] wire240;
  wire [(4'hf):(1'h0)] wire301;
  wire signed [(4'hb):(1'h0)] wire302;
  wire signed [(4'h9):(1'h0)] wire412;
  reg [(4'hc):(1'h0)] reg300 = (1'h0);
  reg [(3'h4):(1'h0)] reg299 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg298 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg297 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg296 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg295 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg293 = (1'h0);
  reg [(2'h3):(1'h0)] reg289 = (1'h0);
  reg [(4'ha):(1'h0)] reg282 = (1'h0);
  reg [(4'hf):(1'h0)] reg281 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg277 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg294 = (1'h0);
  reg signed [(4'he):(1'h0)] reg292 = (1'h0);
  reg [(4'hb):(1'h0)] reg291 = (1'h0);
  reg [(2'h3):(1'h0)] reg290 = (1'h0);
  reg [(4'h8):(1'h0)] reg288 = (1'h0);
  reg [(3'h4):(1'h0)] reg287 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg286 = (1'h0);
  reg signed [(4'he):(1'h0)] reg285 = (1'h0);
  reg [(4'ha):(1'h0)] reg284 = (1'h0);
  reg [(4'h8):(1'h0)] reg283 = (1'h0);
  reg [(3'h7):(1'h0)] reg268 = (1'h0);
  reg [(4'h9):(1'h0)] reg263 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg272 = (1'h0);
  reg [(3'h6):(1'h0)] reg267 = (1'h0);
  reg [(4'hb):(1'h0)] reg262 = (1'h0);
  reg [(4'he):(1'h0)] reg280 = (1'h0);
  reg [(3'h6):(1'h0)] reg279 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg278 = (1'h0);
  reg [(2'h2):(1'h0)] reg276 = (1'h0);
  reg [(2'h2):(1'h0)] reg275 = (1'h0);
  reg [(4'h9):(1'h0)] reg274 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg271 = (1'h0);
  reg [(2'h3):(1'h0)] reg270 = (1'h0);
  reg [(4'ha):(1'h0)] reg269 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg266 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg265 = (1'h0);
  reg [(3'h6):(1'h0)] reg264 = (1'h0);
  reg [(4'ha):(1'h0)] reg252 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg250 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg243 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg242 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg261 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg260 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg259 = (1'h0);
  reg [(3'h6):(1'h0)] reg258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg256 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg255 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg253 = (1'h0);
  reg [(4'ha):(1'h0)] reg251 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg248 = (1'h0);
  reg [(4'h8):(1'h0)] reg247 = (1'h0);
  reg [(4'hc):(1'h0)] reg246 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg245 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg244 = (1'h0);
  reg signed [(4'he):(1'h0)] reg241 = (1'h0);
  reg signed [(4'he):(1'h0)] reg229 = (1'h0);
  reg [(4'hd):(1'h0)] reg228 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg238 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg237 = (1'h0);
  reg [(4'he):(1'h0)] reg236 = (1'h0);
  reg signed [(4'he):(1'h0)] reg235 = (1'h0);
  reg [(2'h2):(1'h0)] reg234 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg233 = (1'h0);
  reg [(3'h4):(1'h0)] reg232 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg230 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg227 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg226 = (1'h0);
  reg [(4'h9):(1'h0)] reg225 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg224 = (1'h0);
  reg [(4'hd):(1'h0)] reg223 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg221 = (1'h0);
  reg [(5'h10):(1'h0)] reg222 = (1'h0);
  reg [(3'h4):(1'h0)] reg209 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg219 = (1'h0);
  reg [(5'h10):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg216 = (1'h0);
  reg [(4'ha):(1'h0)] reg215 = (1'h0);
  reg [(4'hd):(1'h0)] reg214 = (1'h0);
  reg [(3'h7):(1'h0)] reg213 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg212 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg211 = (1'h0);
  reg [(4'hb):(1'h0)] reg210 = (1'h0);
  reg [(4'he):(1'h0)] reg208 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg207 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg206 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg204 = (1'h0);
  reg [(2'h2):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg202 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg201 = (1'h0);
  reg [(4'hd):(1'h0)] reg200 = (1'h0);
  reg [(4'he):(1'h0)] reg199 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg198 = (1'h0);
  reg [(4'h8):(1'h0)] reg197 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg195 = (1'h0);
  reg [(4'hb):(1'h0)] reg194 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg193 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg191 = (1'h0);
  reg [(4'hb):(1'h0)] reg188 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg187 = (1'h0);
  reg [(2'h3):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg183 = (1'h0);
  reg [(4'h9):(1'h0)] reg182 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg181 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg178 = (1'h0);
  reg [(4'h9):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg176 = (1'h0);
  reg [(4'hf):(1'h0)] reg174 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg170 = (1'h0);
  reg [(4'he):(1'h0)] reg172 = (1'h0);
  reg [(5'h10):(1'h0)] reg171 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg169 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg167 = (1'h0);
  reg [(3'h7):(1'h0)] reg162 = (1'h0);
  reg [(4'h8):(1'h0)] reg168 = (1'h0);
  reg [(4'ha):(1'h0)] reg166 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg165 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg164 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg163 = (1'h0);
  reg [(4'hb):(1'h0)] reg161 = (1'h0);
  reg [(3'h4):(1'h0)] reg160 = (1'h0);
  reg [(3'h7):(1'h0)] reg159 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg157 = (1'h0);
  reg [(3'h5):(1'h0)] reg156 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg155 = (1'h0);
  reg [(4'he):(1'h0)] reg154 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg153 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg152 = (1'h0);
  reg [(3'h4):(1'h0)] reg151 = (1'h0);
  reg [(3'h5):(1'h0)] reg149 = (1'h0);
  reg [(4'hb):(1'h0)] reg148 = (1'h0);
  reg [(2'h3):(1'h0)] reg147 = (1'h0);
  reg [(4'he):(1'h0)] reg146 = (1'h0);
  reg [(4'h9):(1'h0)] reg135 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg144 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg143 = (1'h0);
  reg [(4'hf):(1'h0)] reg142 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg141 = (1'h0);
  reg [(3'h7):(1'h0)] reg139 = (1'h0);
  reg [(4'hc):(1'h0)] reg138 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg137 = (1'h0);
  reg [(3'h7):(1'h0)] reg136 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg134 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg133 = (1'h0);
  reg [(4'hc):(1'h0)] reg132 = (1'h0);
  reg [(3'h7):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg130 = (1'h0);
  reg [(4'he):(1'h0)] reg129 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg128 = (1'h0);
  reg [(3'h6):(1'h0)] reg127 = (1'h0);
  reg [(4'h9):(1'h0)] reg126 = (1'h0);
  reg [(4'ha):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg124 = (1'h0);
  reg [(2'h3):(1'h0)] reg123 = (1'h0);
  reg [(5'h10):(1'h0)] reg122 = (1'h0);
  reg [(3'h7):(1'h0)] reg121 = (1'h0);
  reg [(3'h5):(1'h0)] reg120 = (1'h0);
  reg [(4'h9):(1'h0)] reg118 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg117 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg116 = (1'h0);
  reg [(4'h9):(1'h0)] reg115 = (1'h0);
  reg [(4'he):(1'h0)] reg102 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg98 = (1'h0);
  reg [(4'hd):(1'h0)] reg111 = (1'h0);
  reg [(4'ha):(1'h0)] reg110 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg109 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg108 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg106 = (1'h0);
  reg [(2'h2):(1'h0)] reg105 = (1'h0);
  reg [(3'h7):(1'h0)] reg104 = (1'h0);
  reg [(4'hd):(1'h0)] reg103 = (1'h0);
  reg [(3'h6):(1'h0)] reg101 = (1'h0);
  reg [(4'he):(1'h0)] reg100 = (1'h0);
  reg [(3'h5):(1'h0)] reg99 = (1'h0);
  reg [(4'ha):(1'h0)] reg97 = (1'h0);
  reg [(4'ha):(1'h0)] reg95 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg94 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg92 = (1'h0);
  reg [(4'he):(1'h0)] reg88 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg76 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg91 = (1'h0);
  reg [(4'hb):(1'h0)] reg90 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg87 = (1'h0);
  reg signed [(4'he):(1'h0)] reg86 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg85 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg83 = (1'h0);
  reg [(4'hc):(1'h0)] reg82 = (1'h0);
  reg [(4'h8):(1'h0)] reg81 = (1'h0);
  reg [(4'h9):(1'h0)] reg80 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg79 = (1'h0);
  reg [(3'h4):(1'h0)] reg78 = (1'h0);
  reg signed [(4'he):(1'h0)] reg75 = (1'h0);
  reg [(3'h7):(1'h0)] reg74 = (1'h0);
  reg [(4'hb):(1'h0)] reg73 = (1'h0);
  reg [(3'h7):(1'h0)] reg72 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg71 = (1'h0);
  reg [(4'ha):(1'h0)] reg70 = (1'h0);
  reg [(4'hb):(1'h0)] reg68 = (1'h0);
  reg [(4'hd):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg66 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg65 = (1'h0);
  reg [(4'ha):(1'h0)] reg64 = (1'h0);
  reg [(4'hd):(1'h0)] reg63 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg60 = (1'h0);
  reg [(5'h10):(1'h0)] reg44 = (1'h0);
  reg [(2'h2):(1'h0)] reg30 = (1'h0);
  reg [(4'ha):(1'h0)] reg27 = (1'h0);
  reg [(3'h7):(1'h0)] reg22 = (1'h0);
  reg [(4'h8):(1'h0)] reg19 = (1'h0);
  reg [(4'hb):(1'h0)] reg16 = (1'h0);
  reg [(4'h9):(1'h0)] reg15 = (1'h0);
  reg [(4'h9):(1'h0)] reg14 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6 = (1'h0);
  reg [(2'h3):(1'h0)] reg61 = (1'h0);
  reg [(4'h9):(1'h0)] reg59 = (1'h0);
  reg [(4'ha):(1'h0)] reg58 = (1'h0);
  reg [(4'ha):(1'h0)] reg57 = (1'h0);
  reg [(4'he):(1'h0)] reg56 = (1'h0);
  reg [(3'h5):(1'h0)] reg55 = (1'h0);
  reg [(4'ha):(1'h0)] reg54 = (1'h0);
  reg [(2'h3):(1'h0)] reg53 = (1'h0);
  reg [(4'he):(1'h0)] reg52 = (1'h0);
  reg [(4'h9):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg48 = (1'h0);
  reg [(3'h6):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg45 = (1'h0);
  reg [(2'h3):(1'h0)] reg42 = (1'h0);
  reg [(4'he):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg39 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg40 = (1'h0);
  reg [(4'ha):(1'h0)] reg38 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg37 = (1'h0);
  reg [(4'h9):(1'h0)] reg36 = (1'h0);
  reg [(3'h6):(1'h0)] reg35 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg34 = (1'h0);
  reg [(3'h4):(1'h0)] reg33 = (1'h0);
  reg [(4'h8):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg31 = (1'h0);
  reg [(4'he):(1'h0)] reg29 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg28 = (1'h0);
  reg [(4'hc):(1'h0)] reg26 = (1'h0);
  reg [(3'h5):(1'h0)] reg25 = (1'h0);
  reg [(3'h4):(1'h0)] reg24 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg23 = (1'h0);
  reg [(3'h4):(1'h0)] reg21 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg20 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg13 = (1'h0);
  reg [(4'h9):(1'h0)] reg12 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg11 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg10 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg9 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg8 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar288 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar287 = (1'h0);
  reg [(5'h10):(1'h0)] forvar283 = (1'h0);
  reg [(3'h5):(1'h0)] forvar279 = (1'h0);
  reg [(3'h7):(1'h0)] forvar293 = (1'h0);
  reg [(3'h4):(1'h0)] forvar289 = (1'h0);
  reg [(4'h9):(1'h0)] forvar282 = (1'h0);
  reg [(4'hf):(1'h0)] forvar281 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar275 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar274 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar270 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar277 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar272 = (1'h0);
  reg [(4'hc):(1'h0)] forvar268 = (1'h0);
  reg [(5'h10):(1'h0)] forvar267 = (1'h0);
  reg [(2'h3):(1'h0)] forvar263 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar262 = (1'h0);
  reg [(4'hc):(1'h0)] forvar241 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar257 = (1'h0);
  reg [(4'hb):(1'h0)] forvar254 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar252 = (1'h0);
  reg [(3'h5):(1'h0)] forvar250 = (1'h0);
  reg [(2'h3):(1'h0)] forvar243 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar242 = (1'h0);
  reg [(4'h9):(1'h0)] forvar224 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar222 = (1'h0);
  reg [(4'hd):(1'h0)] forvar229 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar228 = (1'h0);
  reg [(4'hd):(1'h0)] forvar221 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar220 = (1'h0);
  reg [(4'ha):(1'h0)] forvar211 = (1'h0);
  reg [(4'hf):(1'h0)] forvar208 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar217 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar209 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar205 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar201 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar196 = (1'h0);
  reg [(4'he):(1'h0)] forvar192 = (1'h0);
  reg [(3'h7):(1'h0)] forvar190 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar189 = (1'h0);
  reg [(2'h3):(1'h0)] forvar184 = (1'h0);
  reg [(4'h9):(1'h0)] forvar180 = (1'h0);
  reg [(3'h6):(1'h0)] forvar179 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar175 = (1'h0);
  reg [(4'he):(1'h0)] forvar165 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar170 = (1'h0);
  reg [(4'ha):(1'h0)] forvar166 = (1'h0);
  reg [(2'h2):(1'h0)] forvar163 = (1'h0);
  reg [(3'h5):(1'h0)] forvar159 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar167 = (1'h0);
  reg [(4'hb):(1'h0)] forvar162 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar158 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar150 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar145 = (1'h0);
  reg [(4'hf):(1'h0)] forvar140 = (1'h0);
  reg [(4'ha):(1'h0)] forvar135 = (1'h0);
  reg [(2'h2):(1'h0)] forvar124 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar126 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar119 = (1'h0);
  reg [(3'h4):(1'h0)] forvar114 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar113 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar112 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar107 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar102 = (1'h0);
  reg [(3'h4):(1'h0)] forvar98 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar96 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar83 = (1'h0);
  reg [(3'h6):(1'h0)] forvar75 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar73 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar89 = (1'h0);
  reg [(4'he):(1'h0)] forvar88 = (1'h0);
  reg [(5'h10):(1'h0)] forvar77 = (1'h0);
  reg [(3'h5):(1'h0)] forvar76 = (1'h0);
  reg [(4'ha):(1'h0)] forvar69 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar62 = (1'h0);
  reg [(4'hb):(1'h0)] forvar59 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar57 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar51 = (1'h0);
  reg [(2'h2):(1'h0)] forvar41 = (1'h0);
  reg [(2'h3):(1'h0)] forvar40 = (1'h0);
  reg [(5'h10):(1'h0)] forvar36 = (1'h0);
  reg [(3'h6):(1'h0)] forvar31 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar21 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar9 = (1'h0);
  reg [(4'ha):(1'h0)] forvar11 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar60 = (1'h0);
  reg [(4'hc):(1'h0)] forvar50 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar49 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar46 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar44 = (1'h0);
  reg [(4'hc):(1'h0)] forvar43 = (1'h0);
  reg [(4'hf):(1'h0)] forvar39 = (1'h0);
  reg [(4'h9):(1'h0)] forvar26 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar30 = (1'h0);
  reg [(5'h10):(1'h0)] forvar27 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar22 = (1'h0);
  reg [(3'h5):(1'h0)] forvar19 = (1'h0);
  reg [(4'hd):(1'h0)] forvar18 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar16 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar15 = (1'h0);
  reg [(3'h7):(1'h0)] forvar14 = (1'h0);
  reg [(3'h7):(1'h0)] forvar7 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6 = (1'h0);
  assign y = {wire418,
                 wire417,
                 wire416,
                 wire415,
                 wire414,
                 wire5,
                 wire239,
                 wire240,
                 wire301,
                 wire302,
                 wire412,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg293,
                 reg289,
                 reg282,
                 reg281,
                 reg277,
                 reg294,
                 reg292,
                 reg291,
                 reg290,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg268,
                 reg263,
                 reg272,
                 reg267,
                 reg262,
                 reg280,
                 reg279,
                 reg278,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg271,
                 reg270,
                 reg269,
                 reg266,
                 reg265,
                 reg264,
                 reg252,
                 reg250,
                 reg243,
                 reg242,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg256,
                 reg255,
                 reg253,
                 reg251,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg241,
                 reg229,
                 reg228,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg221,
                 reg222,
                 reg209,
                 reg219,
                 reg218,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg208,
                 reg207,
                 reg206,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg195,
                 reg194,
                 reg193,
                 reg191,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg183,
                 reg182,
                 reg181,
                 reg178,
                 reg177,
                 reg176,
                 reg174,
                 reg173,
                 reg170,
                 reg172,
                 reg171,
                 reg169,
                 reg167,
                 reg162,
                 reg168,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg161,
                 reg160,
                 reg159,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg135,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg102,
                 reg98,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg101,
                 reg100,
                 reg99,
                 reg97,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg88,
                 reg77,
                 reg76,
                 reg91,
                 reg90,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg60,
                 reg44,
                 reg30,
                 reg27,
                 reg22,
                 reg19,
                 reg16,
                 reg15,
                 reg14,
                 reg7,
                 reg6,
                 reg61,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg48,
                 reg47,
                 reg45,
                 reg42,
                 reg41,
                 reg39,
                 reg40,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg29,
                 reg28,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg21,
                 reg20,
                 reg17,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 forvar288,
                 forvar287,
                 forvar283,
                 forvar279,
                 forvar293,
                 forvar289,
                 forvar282,
                 forvar281,
                 forvar275,
                 forvar274,
                 forvar270,
                 forvar277,
                 forvar272,
                 forvar268,
                 forvar267,
                 forvar263,
                 forvar262,
                 forvar241,
                 forvar257,
                 forvar254,
                 forvar252,
                 forvar250,
                 forvar243,
                 forvar242,
                 forvar224,
                 forvar222,
                 forvar229,
                 forvar228,
                 forvar221,
                 forvar220,
                 forvar211,
                 forvar208,
                 forvar217,
                 forvar209,
                 forvar205,
                 forvar201,
                 forvar196,
                 forvar192,
                 forvar190,
                 forvar189,
                 forvar184,
                 forvar180,
                 forvar179,
                 forvar175,
                 forvar165,
                 forvar170,
                 forvar166,
                 forvar163,
                 forvar159,
                 forvar167,
                 forvar162,
                 forvar158,
                 forvar150,
                 forvar145,
                 forvar140,
                 forvar135,
                 forvar124,
                 forvar126,
                 forvar119,
                 forvar114,
                 forvar113,
                 forvar112,
                 forvar107,
                 forvar102,
                 forvar98,
                 forvar96,
                 forvar83,
                 forvar75,
                 forvar73,
                 forvar89,
                 forvar88,
                 forvar77,
                 forvar76,
                 forvar69,
                 forvar62,
                 forvar59,
                 forvar57,
                 forvar51,
                 forvar41,
                 forvar40,
                 forvar36,
                 forvar31,
                 forvar21,
                 forvar9,
                 forvar11,
                 forvar60,
                 forvar50,
                 forvar49,
                 forvar46,
                 forvar44,
                 forvar43,
                 forvar39,
                 forvar26,
                 forvar30,
                 forvar27,
                 forvar22,
                 forvar19,
                 forvar18,
                 forvar16,
                 forvar15,
                 forvar14,
                 forvar7,
                 forvar6,
                 (1'h0)};
  assign wire5 = $signed(wire0);
  always
    @(posedge clk) begin
      if (($signed(($unsigned(wire4) ?
          {wire1} : wire1[(4'hf):(3'h7)])) ^ wire5[(1'h0):(1'h0)]))
        begin
          for (forvar6 = (1'h0); (forvar6 < (2'h3)); forvar6 = (forvar6 + (1'h1)))
            begin
              for (forvar7 = (1'h0); (forvar7 < (2'h2)); forvar7 = (forvar7 + (1'h1)))
                begin
                  if (((((forvar7 ? wire5 : wire2) ?
                              (forvar7 ? wire1 : forvar7) : (wire0 ?
                                  forvar6 : forvar7)) ?
                          $unsigned($signed(wire3)) : $unsigned((forvar7 ?
                              wire1 : forvar7))) ?
                      wire1 : ((^{wire3}) ?
                          $signed((&wire3)) : wire0[(3'h4):(3'h4)])))
                    begin
                      reg8 <= (8'hb2);
                      reg9 <= wire0;
                      reg10 <= forvar6;
                    end
                  else
                    begin
                      reg8 <= {(reg9 ?
                              (-(^~forvar7)) : $signed($unsigned(reg10)))};
                      reg9 <= $unsigned($signed((~&(wire5 ? wire4 : wire1))));
                      reg10 <= wire5;
                      reg11 <= $signed($unsigned(($signed((8'ha5)) ~^ $signed((8'hb7)))));
                    end
                  reg12 <= $signed($signed($unsigned(forvar6)));
                end
              reg13 <= forvar6;
            end
          for (forvar14 = (1'h0); (forvar14 < (2'h3)); forvar14 = (forvar14 + (1'h1)))
            begin
              for (forvar15 = (1'h0); (forvar15 < (2'h3)); forvar15 = (forvar15 + (1'h1)))
                begin
                  for (forvar16 = (1'h0); (forvar16 < (1'h0)); forvar16 = (forvar16 + (1'h1)))
                    begin
                      reg17 <= (+forvar6);
                    end
                end
              for (forvar18 = (1'h0); (forvar18 < (1'h1)); forvar18 = (forvar18 + (1'h1)))
                begin
                  for (forvar19 = (1'h0); (forvar19 < (2'h2)); forvar19 = (forvar19 + (1'h1)))
                    begin
                      reg20 <= ((forvar14 * (~|$signed((8'hb0)))) <<< $unsigned({$unsigned(forvar6)}));
                    end
                  if (((wire0 ? (~|(8'hb7)) : forvar6[(4'ha):(2'h3)]) ?
                      ((-(reg11 >>> reg10)) ^~ ((forvar14 ?
                          wire0 : (8'ha9)) - $unsigned(forvar7))) : ((^~{(8'hae)}) >>> $signed(reg17))))
                    begin
                      reg21 <= ((forvar14 ?
                          ((reg11 > forvar16) | reg8[(1'h0):(1'h0)]) : ((reg11 ?
                              reg12 : wire5) <= (^~(8'ha0)))) >>> reg10);
                    end
                  else
                    begin
                      reg21 <= (({reg20} | reg8) ?
                          forvar18 : $signed($unsigned((wire2 ?
                              forvar16 : (8'hac)))));
                    end
                  for (forvar22 = (1'h0); (forvar22 < (1'h1)); forvar22 = (forvar22 + (1'h1)))
                    begin
                      reg23 <= reg9[(3'h4):(2'h3)];
                      reg24 <= ($unsigned((+{forvar19})) > (8'haa));
                      reg25 <= reg11;
                    end
                end
            end
          if ((^~{(wire1 || (~|reg10))}))
            begin
              reg26 <= (reg21[(2'h3):(2'h2)] ?
                  forvar7[(1'h0):(1'h0)] : ({reg17[(1'h0):(1'h0)]} ?
                      {wire0} : $signed($signed(reg8))));
              for (forvar27 = (1'h0); (forvar27 < (2'h3)); forvar27 = (forvar27 + (1'h1)))
                begin
                  if (forvar6[(2'h2):(1'h0)])
                    begin
                      reg28 <= ($unsigned((-{reg9})) <= $unsigned((((8'hb8) ?
                          wire5 : (8'hb6)) & $unsigned(wire1))));
                      reg29 <= reg24;
                    end
                  else
                    begin
                      reg28 <= $signed((~((8'ha4) ?
                          (reg8 & reg21) : (-forvar14))));
                      reg29 <= reg24;
                    end
                end
              for (forvar30 = (1'h0); (forvar30 < (1'h1)); forvar30 = (forvar30 + (1'h1)))
                begin
                  if ($unsigned($unsigned(reg10[(1'h0):(1'h0)])))
                    begin
                      reg31 <= $signed(forvar15[(3'h4):(2'h3)]);
                      reg32 <= forvar27;
                    end
                  else
                    begin
                      reg31 <= ($signed(($unsigned(reg21) + (wire3 ?
                          forvar14 : (8'hb0)))) * $unsigned($unsigned({reg10})));
                    end
                  if ((!(8'ha1)))
                    begin
                      reg33 <= (reg13[(3'h6):(2'h3)] ^ forvar27[(3'h5):(2'h2)]);
                      reg34 <= wire0[(4'h9):(1'h1)];
                      reg35 <= $unsigned($signed(((-reg21) < $unsigned(forvar22))));
                      reg36 <= wire2[(4'h8):(1'h1)];
                    end
                  else
                    begin
                      reg33 <= reg35[(3'h4):(1'h1)];
                      reg34 <= wire0[(1'h1):(1'h1)];
                      reg35 <= ((-{(reg35 ?
                              reg31 : (8'hb9))}) + ({reg31} & $signed((reg21 ?
                          forvar22 : wire4))));
                    end
                end
              reg37 <= $signed((forvar19[(1'h0):(1'h0)] - ((|reg9) + $unsigned(reg28))));
            end
          else
            begin
              for (forvar26 = (1'h0); (forvar26 < (2'h2)); forvar26 = (forvar26 + (1'h1)))
                begin
                  for (forvar27 = (1'h0); (forvar27 < (1'h1)); forvar27 = (forvar27 + (1'h1)))
                    begin
                      reg28 <= $signed($unsigned(forvar14[(3'h5):(2'h3)]));
                      reg29 <= forvar6;
                    end
                  for (forvar30 = (1'h0); (forvar30 < (1'h1)); forvar30 = (forvar30 + (1'h1)))
                    begin
                      reg31 <= $signed((+((^~reg33) ?
                          ((8'hb6) * reg10) : reg10)));
                    end
                  if (($signed($unsigned((reg21 ?
                      reg21 : (8'ha1)))) && wire2[(4'h9):(4'h8)]))
                    begin
                      reg32 <= reg20[(4'hc):(4'h8)];
                    end
                  else
                    begin
                      reg32 <= (forvar30[(3'h5):(3'h5)] ?
                          $unsigned(forvar7[(3'h5):(3'h4)]) : (~^($signed(forvar16) <<< wire0)));
                      reg33 <= $unsigned({reg24[(2'h3):(1'h1)]});
                      reg34 <= (~^wire2[(2'h2):(2'h2)]);
                    end
                  if ({(8'hb9)})
                    begin
                      reg35 <= (~&((~(reg36 ?
                          (8'hba) : reg12)) <= $signed($unsigned(reg12))));
                      reg36 <= (^~forvar22[(4'hc):(4'hb)]);
                      reg37 <= forvar30[(5'h10):(4'hd)];
                      reg38 <= wire3;
                    end
                  else
                    begin
                      reg35 <= $signed(reg17);
                      reg36 <= ($signed(($unsigned(forvar16) != (forvar26 <<< (8'hac)))) ?
                          ((reg37 ^~ (reg25 ?
                              reg8 : reg11)) && (forvar7 >= reg35)) : $unsigned(({reg34} ?
                              (forvar30 ? forvar26 : reg37) : (forvar6 ?
                                  forvar18 : forvar18))));
                      reg37 <= {$signed((reg24 << (reg11 ? forvar22 : reg8)))};
                    end
                end
              if ({reg34})
                begin
                  for (forvar39 = (1'h0); (forvar39 < (2'h3)); forvar39 = (forvar39 + (1'h1)))
                    begin
                      reg40 <= $signed((reg32[(3'h7):(3'h7)] ?
                          wire0 : $unsigned((reg33 ? (8'h9e) : reg37))));
                    end
                end
              else
                begin
                  if ((~forvar27[(2'h3):(1'h1)]))
                    begin
                      reg39 <= ($signed((wire2[(1'h0):(1'h0)] >= wire3[(4'hb):(4'ha)])) || (forvar19[(2'h3):(1'h1)] ?
                          $unsigned($signed(reg36)) : $signed(((8'hb7) >> reg10))));
                      reg40 <= ({((wire5 + forvar18) ?
                              reg36[(2'h3):(2'h3)] : {forvar14})} + ((|reg31[(5'h10):(5'h10)]) ?
                          {$signed(forvar30)} : ({reg8} ?
                              (&reg36) : (-forvar39))));
                      reg41 <= (~&$signed($unsigned($signed(forvar16))));
                      reg42 <= $unsigned($signed((8'ha9)));
                    end
                  else
                    begin
                      reg39 <= ($signed({(+forvar16)}) || (reg38[(3'h4):(1'h1)] != ({reg26} * $signed(forvar16))));
                      reg40 <= reg24;
                    end
                end
            end
          for (forvar43 = (1'h0); (forvar43 < (1'h0)); forvar43 = (forvar43 + (1'h1)))
            begin
              for (forvar44 = (1'h0); (forvar44 < (1'h0)); forvar44 = (forvar44 + (1'h1)))
                begin
                  reg45 <= reg23[(3'h6):(3'h6)];
                  for (forvar46 = (1'h0); (forvar46 < (1'h1)); forvar46 = (forvar46 + (1'h1)))
                    begin
                      reg47 <= reg12;
                      reg48 <= ((reg9 ? reg26[(1'h0):(1'h0)] : {{forvar30}}) ?
                          $signed((^~(forvar46 ?
                              reg38 : reg38))) : $signed(reg34[(4'h8):(2'h2)]));
                    end
                end
              for (forvar49 = (1'h0); (forvar49 < (2'h2)); forvar49 = (forvar49 + (1'h1)))
                begin
                  for (forvar50 = (1'h0); (forvar50 < (2'h3)); forvar50 = (forvar50 + (1'h1)))
                    begin
                      reg51 <= ((+forvar18[(3'h6):(1'h0)]) & (-reg31));
                      reg52 <= (^({reg35} >>> reg9));
                      reg53 <= forvar6[(4'ha):(3'h5)];
                      reg54 <= (-wire4);
                    end
                  reg55 <= ($signed(reg29[(3'h4):(3'h4)]) | reg33[(2'h2):(1'h0)]);
                  if ((~^((8'ha9) | (^(+(8'h9f))))))
                    begin
                      reg56 <= (^$signed($unsigned((8'hb1))));
                      reg57 <= (^reg29[(4'h8):(1'h0)]);
                      reg58 <= reg57[(4'h9):(4'h9)];
                      reg59 <= ((8'hb2) <<< $signed({reg36}));
                    end
                  else
                    begin
                      reg56 <= wire0;
                      reg57 <= reg37;
                      reg58 <= (reg33 ? $unsigned(reg39) : (8'h9d));
                      reg59 <= reg54[(4'h8):(3'h7)];
                    end
                  for (forvar60 = (1'h0); (forvar60 < (2'h3)); forvar60 = (forvar60 + (1'h1)))
                    begin
                      reg61 <= wire0[(4'hd):(4'h9)];
                    end
                end
            end
        end
      else
        begin
          if ((-reg40[(3'h5):(2'h2)]))
            begin
              reg6 <= $unsigned((($signed(wire1) ? reg31 : reg56) ?
                  {(8'h9e)} : wire3[(4'h9):(2'h2)]));
            end
          else
            begin
              if (((forvar6[(2'h3):(1'h1)] ?
                      $unsigned((8'hb5)) : ($unsigned(reg9) ?
                          $signed(wire4) : {wire0})) ?
                  (~&(reg41[(4'h8):(3'h4)] * (&reg40))) : {(8'ha8)}))
                begin
                  if (($unsigned(forvar27) <= (^($unsigned(forvar60) < $signed((8'ha6))))))
                    begin
                      reg6 <= $signed({reg25});
                    end
                  else
                    begin
                      reg6 <= $unsigned(($signed(forvar14[(3'h4):(2'h2)]) || wire4[(1'h0):(1'h0)]));
                      reg7 <= reg6;
                    end
                  if ($signed(forvar50))
                    begin
                      reg8 <= $signed((+reg40[(4'ha):(4'h9)]));
                      reg9 <= reg45[(3'h4):(1'h1)];
                      reg10 <= ((&(+reg40)) < reg47[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg8 <= reg35;
                      reg9 <= wire3;
                      reg10 <= (reg6[(4'h9):(1'h1)] ^~ reg11[(1'h1):(1'h0)]);
                    end
                  for (forvar11 = (1'h0); (forvar11 < (1'h1)); forvar11 = (forvar11 + (1'h1)))
                    begin
                      reg12 <= $signed(({forvar15} >= ({reg25} ?
                          $signed(reg37) : {reg38})));
                    end
                  if (wire2)
                    begin
                      reg13 <= reg24[(1'h0):(1'h0)];
                      reg14 <= reg11;
                      reg15 <= (&reg37);
                    end
                  else
                    begin
                      reg13 <= (((+(reg23 == reg54)) ?
                          ($unsigned(forvar7) >> $unsigned(forvar27)) : {$unsigned((8'ha0))}) >>> $unsigned((~|$signed(reg52))));
                      reg14 <= forvar60[(3'h7):(1'h0)];
                      reg15 <= $unsigned($signed((^~$unsigned(reg6))));
                      reg16 <= $unsigned({wire0});
                    end
                end
              else
                begin
                  if (((~&(8'haf)) & reg11))
                    begin
                      reg6 <= reg42;
                      reg7 <= reg8;
                      reg8 <= (forvar11[(1'h0):(1'h0)] ?
                          ((forvar50[(2'h3):(1'h1)] ?
                                  reg54 : (reg25 ? (8'hb1) : reg11)) ?
                              $signed($unsigned(reg36)) : ($unsigned(reg20) * (8'hab))) : {$unsigned(reg56[(1'h0):(1'h0)])});
                    end
                  else
                    begin
                      reg6 <= forvar7;
                      reg7 <= $unsigned(forvar18[(1'h1):(1'h0)]);
                      reg8 <= $signed($signed(forvar22));
                    end
                  for (forvar9 = (1'h0); (forvar9 < (1'h0)); forvar9 = (forvar9 + (1'h1)))
                    begin
                      reg10 <= ((reg34[(2'h3):(1'h0)] ?
                              forvar44 : (|$unsigned(forvar15))) ?
                          (((~|reg17) ?
                              (reg38 ?
                                  forvar19 : (8'hb9)) : forvar15) && {(~^(8'ha1))}) : forvar19);
                      reg11 <= $signed($unsigned($signed($unsigned(reg59))));
                      reg12 <= (-(^$signed(reg55[(2'h3):(2'h2)])));
                      reg13 <= $signed(($unsigned(reg53) ?
                          {((8'ha3) ? reg53 : reg33)} : (-(reg45 ?
                              forvar46 : forvar44))));
                    end
                  if ((reg47[(1'h0):(1'h0)] ?
                      (^(~^$unsigned((8'hb2)))) : forvar9))
                    begin
                      reg14 <= ((forvar60 ?
                              (reg47[(3'h6):(3'h6)] ?
                                  reg41 : $signed(reg9)) : ((reg34 ^ reg51) >= reg6[(4'hd):(4'hb)])) ?
                          wire1 : (~&{$signed(reg36)}));
                      reg15 <= {(((reg26 >> forvar50) ~^ (~(8'h9c))) ?
                              (forvar50 & {reg55}) : reg11)};
                      reg16 <= (!forvar11[(4'ha):(4'h9)]);
                      reg17 <= reg15;
                    end
                  else
                    begin
                      reg14 <= $signed((8'hb2));
                      reg15 <= $unsigned((($unsigned(reg11) ?
                          (reg38 <<< forvar43) : {reg57}) ^~ forvar27));
                      reg16 <= $unsigned((8'ha8));
                      reg17 <= ({reg12} != reg8);
                    end
                end
              for (forvar18 = (1'h0); (forvar18 < (1'h0)); forvar18 = (forvar18 + (1'h1)))
                begin
                  if (reg54[(1'h0):(1'h0)])
                    begin
                      reg19 <= wire0;
                    end
                  else
                    begin
                      reg19 <= (+$signed((~|((8'hb5) * (8'hb2)))));
                    end
                  reg20 <= ($signed(((reg25 ^~ reg9) || ((8'hb2) ?
                      forvar50 : reg58))) ^~ (~&(forvar43[(4'ha):(1'h1)] | $signed(wire5))));
                  for (forvar21 = (1'h0); (forvar21 < (2'h3)); forvar21 = (forvar21 + (1'h1)))
                    begin
                      reg22 <= (((forvar9 ?
                              $signed((8'haa)) : $unsigned(reg38)) ?
                          forvar50[(2'h3):(1'h0)] : forvar14) + $signed(({forvar18} ?
                          $signed(forvar46) : reg6[(4'ha):(3'h5)])));
                    end
                  if (reg17)
                    begin
                      reg23 <= (!reg25);
                    end
                  else
                    begin
                      reg23 <= (($unsigned((reg15 ? reg31 : reg41)) ?
                              ((8'hb5) | {reg40}) : reg59[(3'h7):(3'h4)]) ?
                          $unsigned(reg22) : $unsigned((reg14[(3'h7):(3'h6)] ?
                              {reg6} : forvar11)));
                      reg24 <= reg37[(3'h6):(1'h0)];
                      reg25 <= reg26[(4'hc):(4'ha)];
                      reg26 <= {reg56[(4'hb):(3'h5)]};
                    end
                end
              if ($signed((wire1 < reg41)))
                begin
                  if ({(-((reg45 ? reg45 : forvar46) ?
                          (|reg26) : $unsigned(reg12)))})
                    begin
                      reg27 <= $signed(({reg7} ? reg12[(2'h3):(1'h0)] : reg12));
                      reg28 <= {reg61[(2'h2):(2'h2)]};
                      reg29 <= $signed((reg39 ?
                          $unsigned((forvar44 ?
                              (8'hb6) : (8'ha7))) : {reg53[(1'h1):(1'h1)]}));
                    end
                  else
                    begin
                      reg27 <= ((|(+{forvar21})) ?
                          (forvar46[(4'h9):(2'h2)] ?
                              reg33[(2'h2):(1'h1)] : $unsigned($signed((8'had)))) : {(reg28 < $signed(reg24))});
                    end
                  if ((reg34[(1'h1):(1'h1)] << (({wire0} & $unsigned(reg22)) ?
                      $unsigned((reg48 ? reg48 : reg37)) : (8'hab))))
                    begin
                      reg30 <= {$unsigned((|(&reg42)))};
                    end
                  else
                    begin
                      reg30 <= (~$signed(reg26[(3'h6):(3'h4)]));
                    end
                  for (forvar31 = (1'h0); (forvar31 < (2'h3)); forvar31 = (forvar31 + (1'h1)))
                    begin
                      reg32 <= forvar26;
                      reg33 <= $unsigned(((8'hab) ?
                          (reg55[(1'h0):(1'h0)] ?
                              $signed(reg59) : (^reg35)) : reg21[(1'h1):(1'h0)]));
                      reg34 <= (reg27[(3'h6):(1'h0)] >>> $unsigned((-forvar49)));
                      reg35 <= ($unsigned((~{reg13})) ?
                          ({$signed(reg30)} ^~ {((8'hab) != reg39)}) : $unsigned({reg42[(1'h1):(1'h1)]}));
                    end
                  for (forvar36 = (1'h0); (forvar36 < (2'h3)); forvar36 = (forvar36 + (1'h1)))
                    begin
                      reg37 <= $signed($unsigned(forvar39[(4'hb):(3'h4)]));
                      reg38 <= (8'ha6);
                      reg39 <= $signed(reg42[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar27 = (1'h0); (forvar27 < (1'h0)); forvar27 = (forvar27 + (1'h1)))
                    begin
                      reg28 <= ($signed(reg59[(2'h3):(2'h3)]) ?
                          ({(wire3 ? reg22 : wire4)} ?
                              reg36[(3'h7):(1'h1)] : $unsigned((8'hb2))) : (($signed(forvar21) & ((8'hb7) || wire0)) >> reg59));
                      reg29 <= $unsigned(((reg53 ? reg8 : {(8'hab)}) ?
                          (forvar44[(3'h7):(1'h1)] ~^ ((8'hab) ?
                              reg21 : forvar39)) : (~^(^forvar31))));
                    end
                  for (forvar30 = (1'h0); (forvar30 < (1'h0)); forvar30 = (forvar30 + (1'h1)))
                    begin
                      reg31 <= $signed(($unsigned(((8'hb6) == (8'ha6))) ?
                          (8'ha8) : $unsigned((reg33 ? reg7 : forvar6))));
                      reg32 <= reg30;
                      reg33 <= {($signed($signed(reg52)) ?
                              (reg10 ^ (forvar46 ? reg54 : reg36)) : (8'ha8))};
                      reg34 <= (~reg10[(2'h3):(2'h2)]);
                    end
                  reg35 <= (((forvar7 || {reg9}) || ($signed((8'ha3)) | reg27)) ?
                      (({(8'hac)} >>> forvar7) ?
                          ((wire1 ?
                              forvar16 : forvar11) ^~ reg10) : (^~(^wire2))) : reg21);
                end
              for (forvar40 = (1'h0); (forvar40 < (2'h2)); forvar40 = (forvar40 + (1'h1)))
                begin
                  for (forvar41 = (1'h0); (forvar41 < (2'h2)); forvar41 = (forvar41 + (1'h1)))
                    begin
                      reg42 <= (-$signed(((~^reg45) < $unsigned((8'ha1)))));
                    end
                  for (forvar43 = (1'h0); (forvar43 < (2'h2)); forvar43 = (forvar43 + (1'h1)))
                    begin
                      reg44 <= (+reg30[(1'h0):(1'h0)]);
                      reg45 <= (($unsigned(reg21[(2'h2):(2'h2)]) ?
                          ($unsigned(forvar22) ?
                              (reg56 ?
                                  (8'had) : (8'h9c)) : $signed(reg27)) : reg41[(2'h2):(1'h0)]) >>> (~$signed(reg21[(1'h1):(1'h1)])));
                    end
                  for (forvar46 = (1'h0); (forvar46 < (1'h1)); forvar46 = (forvar46 + (1'h1)))
                    begin
                      reg47 <= (~&forvar43);
                    end
                  reg48 <= $signed($signed(reg54));
                end
            end
          for (forvar49 = (1'h0); (forvar49 < (1'h1)); forvar49 = (forvar49 + (1'h1)))
            begin
              for (forvar50 = (1'h0); (forvar50 < (2'h2)); forvar50 = (forvar50 + (1'h1)))
                begin
                  for (forvar51 = (1'h0); (forvar51 < (2'h3)); forvar51 = (forvar51 + (1'h1)))
                    begin
                      reg52 <= reg51[(3'h5):(1'h1)];
                      reg53 <= ((((~|(8'h9f)) ?
                                  $unsigned(wire1) : ((8'hb3) ?
                                      reg38 : reg44)) ?
                              forvar15 : (wire1[(2'h2):(2'h2)] ?
                                  $signed(reg34) : (reg23 ?
                                      forvar46 : forvar22))) ?
                          forvar41 : reg24);
                      reg54 <= reg61[(1'h0):(1'h0)];
                      reg55 <= (+$signed(($signed(forvar7) * (~|reg19))));
                    end
                  reg56 <= (^~$unsigned(($signed((8'ha5)) ^ $signed(forvar36))));
                end
              for (forvar57 = (1'h0); (forvar57 < (2'h2)); forvar57 = (forvar57 + (1'h1)))
                begin
                  reg58 <= $unsigned((^reg57[(4'h8):(1'h1)]));
                  for (forvar59 = (1'h0); (forvar59 < (1'h0)); forvar59 = (forvar59 + (1'h1)))
                    begin
                      reg60 <= (+reg33);
                      reg61 <= (^~(((reg7 ? forvar6 : reg48) ?
                          $unsigned((8'haa)) : $unsigned(forvar44)) < $unsigned(reg25[(2'h2):(2'h2)])));
                    end
                  for (forvar62 = (1'h0); (forvar62 < (1'h1)); forvar62 = (forvar62 + (1'h1)))
                    begin
                      reg63 <= forvar59;
                      reg64 <= (forvar9[(3'h7):(3'h4)] - (&$signed($signed(reg40))));
                      reg65 <= reg26;
                    end
                  if ($signed(wire5[(1'h1):(1'h1)]))
                    begin
                      reg66 <= $unsigned((8'ha6));
                      reg67 <= $signed((-($signed(reg24) & (reg31 ?
                          reg6 : reg66))));
                      reg68 <= $signed($unsigned($unsigned(wire5[(4'h8):(3'h4)])));
                    end
                  else
                    begin
                      reg66 <= ((|forvar7) & $signed($signed((forvar6 - (8'ha1)))));
                      reg67 <= wire4;
                      reg68 <= (-$signed(forvar21[(3'h7):(2'h2)]));
                    end
                end
            end
          if ((reg54[(4'h9):(3'h4)] ?
              $unsigned($signed($unsigned(reg47))) : $unsigned((reg52 > $unsigned(reg11)))))
            begin
              for (forvar69 = (1'h0); (forvar69 < (2'h2)); forvar69 = (forvar69 + (1'h1)))
                begin
                  reg70 <= forvar57;
                  if ((reg7[(4'he):(4'hd)] < $signed({(forvar31 * reg15)})))
                    begin
                      reg71 <= $unsigned((~&(^~(reg52 ^ reg11))));
                      reg72 <= (+(reg29 ?
                          (forvar41[(1'h0):(1'h0)] ~^ (reg44 <<< forvar9)) : {((8'hb5) ?
                                  reg13 : reg29)}));
                    end
                  else
                    begin
                      reg71 <= (($unsigned($unsigned(forvar62)) * forvar46) ?
                          $unsigned(((reg68 ?
                              reg35 : reg53) > (~^reg44))) : (~((~(8'ha9)) ?
                              (reg17 ? forvar19 : reg61) : (&forvar19))));
                    end
                  if ($signed(((forvar59 & (reg6 != (8'hb6))) >> forvar31[(1'h0):(1'h0)])))
                    begin
                      reg73 <= $signed($signed((!(~|(8'hb4)))));
                      reg74 <= {(($unsigned(reg59) ?
                                  (~&reg55) : (forvar43 ? forvar18 : reg37)) ?
                              (+$signed(reg21)) : $signed((reg68 ?
                                  reg13 : reg25)))};
                      reg75 <= (~^$unsigned((^~$signed(forvar51))));
                    end
                  else
                    begin
                      reg73 <= ((^({reg73} ?
                              (~|reg15) : (reg53 ? reg52 : forvar21))) ?
                          $unsigned(reg60[(4'h9):(3'h5)]) : reg17);
                      reg74 <= (reg65[(3'h4):(2'h3)] != reg12);
                      reg75 <= (~|$signed((&{(8'h9d)})));
                    end
                end
              for (forvar76 = (1'h0); (forvar76 < (2'h3)); forvar76 = (forvar76 + (1'h1)))
                begin
                  for (forvar77 = (1'h0); (forvar77 < (1'h0)); forvar77 = (forvar77 + (1'h1)))
                    begin
                      reg78 <= $signed($signed((|(8'ha0))));
                      reg79 <= {(reg63[(4'h8):(2'h3)] ?
                              (reg74[(3'h5):(2'h2)] >>> {(8'ha1)}) : (reg15[(1'h0):(1'h0)] - forvar18[(4'h8):(3'h7)]))};
                      reg80 <= (wire4 ?
                          reg41 : (($unsigned((8'ha1)) && $unsigned(reg40)) > (^forvar39)));
                    end
                  if (((((forvar49 ? (8'h9d) : forvar15) ?
                          reg10 : (~&forvar39)) > (~&$unsigned(reg11))) ?
                      $signed($signed(forvar51[(4'h9):(3'h7)])) : $signed($signed(reg26))))
                    begin
                      reg81 <= (reg59[(1'h0):(1'h0)] ?
                          ((|$signed(reg9)) ?
                              {reg30} : {$unsigned(reg45)}) : forvar41[(2'h2):(2'h2)]);
                      reg82 <= (~^reg79[(1'h1):(1'h1)]);
                      reg83 <= reg59[(4'h9):(4'h8)];
                      reg84 <= ((reg42 ?
                          reg9[(4'h9):(4'h8)] : reg83) <<< (reg20[(2'h3):(2'h2)] ?
                          ((reg70 ?
                              reg71 : reg47) + (8'hb7)) : ($unsigned(forvar60) ?
                              $unsigned(reg71) : (~&forvar62))));
                    end
                  else
                    begin
                      reg81 <= $signed(($unsigned((reg83 <= forvar14)) < (reg70[(3'h7):(1'h0)] ?
                          $signed(reg8) : $unsigned(forvar59))));
                      reg82 <= forvar31[(3'h5):(2'h2)];
                    end
                  if ($signed(reg26))
                    begin
                      reg85 <= $signed((8'h9e));
                    end
                  else
                    begin
                      reg85 <= $unsigned($signed(({(8'ha9)} + forvar41)));
                      reg86 <= {$unsigned((reg40[(1'h1):(1'h1)] * (~&forvar39)))};
                      reg87 <= {(&((reg81 && reg60) >= forvar77))};
                    end
                end
              for (forvar88 = (1'h0); (forvar88 < (2'h2)); forvar88 = (forvar88 + (1'h1)))
                begin
                  for (forvar89 = (1'h0); (forvar89 < (1'h0)); forvar89 = (forvar89 + (1'h1)))
                    begin
                      reg90 <= forvar19;
                      reg91 <= $signed(forvar51[(4'hd):(3'h4)]);
                    end
                end
            end
          else
            begin
              for (forvar69 = (1'h0); (forvar69 < (2'h3)); forvar69 = (forvar69 + (1'h1)))
                begin
                  if (reg73[(3'h4):(1'h0)])
                    begin
                      reg70 <= (!$signed(((~reg33) ?
                          (reg84 * (8'h9d)) : $unsigned(forvar39))));
                    end
                  else
                    begin
                      reg70 <= (&$unsigned(reg35));
                      reg71 <= {forvar18[(4'ha):(4'h9)]};
                      reg72 <= $unsigned($unsigned(forvar51[(2'h2):(1'h1)]));
                    end
                  for (forvar73 = (1'h0); (forvar73 < (2'h3)); forvar73 = (forvar73 + (1'h1)))
                    begin
                      reg74 <= $unsigned($unsigned(($unsigned(reg67) >> $signed(reg13))));
                    end
                end
              if ($signed((forvar89[(3'h7):(2'h2)] ?
                  ((reg66 ^ (8'hac)) * $unsigned(reg57)) : ($unsigned(reg59) != reg87[(4'hd):(4'hb)]))))
                begin
                  for (forvar75 = (1'h0); (forvar75 < (1'h0)); forvar75 = (forvar75 + (1'h1)))
                    begin
                      reg76 <= (~$signed($unsigned((^~forvar75))));
                      reg77 <= $unsigned(((~&((8'ha6) ? reg24 : wire4)) ?
                          $signed({reg65}) : $unsigned((&(8'h9e)))));
                      reg78 <= ((((reg91 ? reg79 : reg29) < (forvar50 ?
                                  reg33 : reg61)) ?
                              reg35 : forvar19) ?
                          {($signed(reg30) ?
                                  (reg53 == forvar49) : ((8'hba) ?
                                      (8'ha3) : reg85))} : (-reg87[(4'h9):(2'h2)]));
                    end
                  if (reg44)
                    begin
                      reg79 <= (($unsigned({reg78}) ?
                          $unsigned(((8'hac) >= reg59)) : (^~(-reg28))) == (~|reg86));
                      reg80 <= reg36[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg79 <= reg23[(2'h2):(2'h2)];
                      reg80 <= ((($unsigned(forvar36) ?
                              (+(8'ha2)) : $signed(forvar76)) ?
                          $signed({forvar26}) : reg36) >> ($unsigned((reg38 | forvar43)) ?
                          $unsigned(forvar36[(4'h9):(4'h9)]) : reg32[(2'h2):(1'h0)]));
                      reg81 <= ($unsigned(((reg75 << reg47) - $unsigned(reg90))) + reg39);
                      reg82 <= wire3;
                    end
                  for (forvar83 = (1'h0); (forvar83 < (2'h2)); forvar83 = (forvar83 + (1'h1)))
                    begin
                      reg84 <= ($unsigned($unsigned(wire5)) ?
                          ((forvar60[(3'h7):(3'h5)] ?
                              reg71[(1'h0):(1'h0)] : reg76) != (8'hb9)) : (8'hb5));
                      reg85 <= $unsigned(reg77[(1'h1):(1'h0)]);
                      reg86 <= $signed({{(reg85 ? reg40 : reg40)}});
                      reg87 <= $signed((&$signed($unsigned(forvar40))));
                    end
                  reg88 <= reg78;
                end
              else
                begin
                  for (forvar75 = (1'h0); (forvar75 < (1'h0)); forvar75 = (forvar75 + (1'h1)))
                    begin
                      reg76 <= $unsigned(reg42);
                      reg77 <= ((((reg14 || (8'hb5)) ?
                          reg76 : $unsigned(forvar73)) * ((~&reg7) ~^ reg65)) ^~ ($signed((reg77 >>> (8'h9d))) * $signed((forvar62 > forvar19))));
                      reg78 <= forvar30[(4'h8):(3'h5)];
                      reg79 <= ((~|reg90) > (8'hae));
                    end
                end
              for (forvar89 = (1'h0); (forvar89 < (1'h0)); forvar89 = (forvar89 + (1'h1)))
                begin
                  reg90 <= reg39;
                  if (((forvar62[(3'h5):(3'h4)] ?
                      reg21 : $signed($signed((8'had)))) >>> $unsigned({(reg23 ?
                          reg10 : forvar59)})))
                    begin
                      reg91 <= {(reg35[(2'h3):(2'h3)] || (reg55 | reg44))};
                    end
                  else
                    begin
                      reg91 <= (8'hb7);
                    end
                  if ((^~$signed((forvar69 ? $signed(forvar43) : (8'hb1)))))
                    begin
                      reg92 <= (~&(&forvar26));
                      reg93 <= reg15[(3'h5):(2'h3)];
                      reg94 <= $unsigned($signed(((reg22 < forvar49) - $signed((8'hac)))));
                      reg95 <= {reg53};
                    end
                  else
                    begin
                      reg92 <= (8'hb5);
                    end
                end
            end
          for (forvar96 = (1'h0); (forvar96 < (1'h1)); forvar96 = (forvar96 + (1'h1)))
            begin
              reg97 <= forvar89[(1'h1):(1'h0)];
              if ($signed(((!(forvar39 == (8'hb8))) > $signed($signed(reg55)))))
                begin
                  for (forvar98 = (1'h0); (forvar98 < (2'h2)); forvar98 = (forvar98 + (1'h1)))
                    begin
                      reg99 <= $signed(((((8'hb6) ?
                          reg83 : reg44) ^ reg57[(3'h6):(3'h4)]) | reg52[(4'h8):(2'h2)]));
                      reg100 <= ($unsigned($unsigned((~reg84))) ?
                          reg76 : (($unsigned(reg74) ^ (!forvar16)) ?
                              $signed(reg85[(3'h6):(3'h6)]) : ((+forvar26) != forvar62)));
                      reg101 <= reg23;
                    end
                  for (forvar102 = (1'h0); (forvar102 < (1'h0)); forvar102 = (forvar102 + (1'h1)))
                    begin
                      reg103 <= (&(~$signed(reg63)));
                      reg104 <= $unsigned(($signed((forvar30 ^ (8'haf))) >> ((reg19 ?
                          forvar39 : reg16) == (forvar77 ? reg47 : reg40))));
                      reg105 <= ({($signed(reg7) < reg81[(4'h8):(2'h3)])} ?
                          reg64[(1'h1):(1'h1)] : (~^reg87[(4'h9):(1'h1)]));
                      reg106 <= reg86;
                    end
                  for (forvar107 = (1'h0); (forvar107 < (2'h3)); forvar107 = (forvar107 + (1'h1)))
                    begin
                      reg108 <= (~&reg77);
                      reg109 <= {$signed($signed(forvar51[(4'hc):(3'h6)]))};
                      reg110 <= {reg23[(2'h3):(1'h1)]};
                      reg111 <= (8'h9e);
                    end
                end
              else
                begin
                  reg98 <= $signed((&forvar9));
                  if (($unsigned($unsigned((reg38 ? reg13 : reg66))) ?
                      ((~|$signed((8'h9e))) ?
                          reg20[(4'ha):(4'h9)] : $signed(reg58)) : (reg73[(2'h3):(2'h3)] ?
                          reg88 : ((forvar50 > forvar44) == (&reg87)))))
                    begin
                      reg99 <= (reg85[(2'h2):(1'h1)] ?
                          (reg80 > forvar69[(1'h0):(1'h0)]) : (reg47 == ((reg54 ?
                                  (8'hb6) : reg57) ?
                              reg22 : (reg19 ? reg44 : reg35))));
                      reg100 <= reg13;
                      reg101 <= ($signed((forvar41[(1'h0):(1'h0)] >>> (reg38 ^ forvar77))) ?
                          $unsigned(reg73[(3'h4):(1'h1)]) : $signed(forvar69));
                      reg102 <= ((forvar41[(2'h2):(1'h0)] ?
                          reg38 : $signed(reg88[(4'hb):(1'h1)])) > ($signed((reg37 >>> wire4)) ?
                          $unsigned($signed(reg55)) : $unsigned((forvar77 ?
                              reg16 : forvar39))));
                    end
                  else
                    begin
                      reg99 <= (~^(~^((^~reg93) ?
                          $signed(wire3) : $signed(reg105))));
                      reg100 <= reg63;
                      reg101 <= $signed($unsigned(forvar77));
                      reg102 <= ($unsigned(forvar21) | reg111[(2'h2):(2'h2)]);
                    end
                  if ($unsigned($unsigned(reg98)))
                    begin
                      reg103 <= {{$unsigned(reg80[(3'h5):(3'h5)])}};
                      reg104 <= $unsigned(forvar77[(4'he):(4'ha)]);
                      reg105 <= $signed(forvar77[(1'h0):(1'h0)]);
                      reg106 <= {($signed((reg30 ?
                              reg75 : reg79)) == reg71[(1'h1):(1'h1)])};
                    end
                  else
                    begin
                      reg103 <= (~$unsigned(forvar51[(3'h4):(1'h1)]));
                      reg104 <= $signed((^~(&reg32[(3'h4):(2'h3)])));
                      reg105 <= $unsigned({$unsigned((reg71 ? reg63 : reg11))});
                    end
                end
            end
        end
      for (forvar112 = (1'h0); (forvar112 < (1'h0)); forvar112 = (forvar112 + (1'h1)))
        begin
          for (forvar113 = (1'h0); (forvar113 < (1'h1)); forvar113 = (forvar113 + (1'h1)))
            begin
              for (forvar114 = (1'h0); (forvar114 < (1'h0)); forvar114 = (forvar114 + (1'h1)))
                begin
                  if ((8'hb2))
                    begin
                      reg115 <= (~|(&reg77));
                      reg116 <= $unsigned(reg9);
                      reg117 <= $unsigned(($signed($unsigned(reg59)) == reg86));
                      reg118 <= $signed(forvar73);
                    end
                  else
                    begin
                      reg115 <= (^~$unsigned((+reg41[(4'h9):(3'h5)])));
                      reg116 <= (reg98 ? reg40 : $signed((+{reg103})));
                      reg117 <= (forvar41 ?
                          (forvar15[(1'h0):(1'h0)] >>> reg97[(4'ha):(3'h6)]) : reg104[(3'h6):(2'h3)]);
                      reg118 <= reg44;
                    end
                  for (forvar119 = (1'h0); (forvar119 < (2'h3)); forvar119 = (forvar119 + (1'h1)))
                    begin
                      reg120 <= (|$signed((^~$signed(reg15))));
                      reg121 <= reg53;
                      reg122 <= forvar60[(3'h6):(3'h6)];
                      reg123 <= (wire5[(4'h9):(4'h9)] >>> $unsigned(reg53));
                    end
                end
            end
          if ($signed($signed(reg6)))
            begin
              if (((!$signed(forvar119)) >> $signed($signed((~&(8'hb4))))))
                begin
                  reg124 <= ((forvar113 ?
                      $unsigned(forvar113[(4'hb):(4'h9)]) : $signed(reg73[(2'h3):(1'h1)])) < (|forvar113));
                  if ((&(+((-reg74) ? (forvar27 == reg84) : (^(8'ha5))))))
                    begin
                      reg125 <= $signed((+forvar51[(3'h5):(2'h3)]));
                      reg126 <= forvar7[(3'h7):(3'h4)];
                      reg127 <= reg117[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg125 <= (&$unsigned(($signed(forvar31) > (reg67 ?
                          reg32 : forvar26))));
                      reg126 <= (($signed(forvar19[(2'h2):(2'h2)]) >= {(~|(8'hba))}) + ({(forvar113 < reg54)} < ($unsigned(reg15) ?
                          $unsigned(reg15) : $unsigned(forvar46))));
                    end
                end
              else
                begin
                  if ((({$unsigned(reg111)} ?
                          (8'h9f) : $unsigned(reg73[(1'h1):(1'h1)])) ?
                      reg56 : ((forvar15[(1'h1):(1'h0)] & (-reg115)) ?
                          forvar50 : forvar31)))
                    begin
                      reg124 <= $signed((forvar113 ?
                          $unsigned({reg109}) : (^$unsigned(reg109))));
                      reg125 <= reg42[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg124 <= $unsigned((~^reg105));
                    end
                  for (forvar126 = (1'h0); (forvar126 < (2'h2)); forvar126 = (forvar126 + (1'h1)))
                    begin
                      reg127 <= $unsigned(reg55[(3'h4):(3'h4)]);
                      reg128 <= reg11[(4'h8):(1'h0)];
                      reg129 <= $unsigned((~|reg84[(2'h3):(2'h2)]));
                    end
                end
            end
          else
            begin
              for (forvar124 = (1'h0); (forvar124 < (2'h2)); forvar124 = (forvar124 + (1'h1)))
                begin
                  reg125 <= $signed((((reg92 ^~ reg74) <<< $signed(reg35)) ^~ (reg125[(3'h7):(3'h6)] ?
                      (+forvar60) : (wire4 ? forvar57 : reg14))));
                  for (forvar126 = (1'h0); (forvar126 < (1'h0)); forvar126 = (forvar126 + (1'h1)))
                    begin
                      reg127 <= $signed({((reg61 ? reg121 : forvar15) ?
                              ((8'ha5) | reg21) : $signed((8'hab)))});
                    end
                  reg128 <= {reg87};
                  if ((!$signed({(wire0 ? forvar36 : reg68)})))
                    begin
                      reg129 <= $unsigned((|reg36[(3'h7):(2'h3)]));
                      reg130 <= $signed(reg22[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg129 <= ((~^forvar27[(4'ha):(2'h3)]) ?
                          {$unsigned($signed((8'hb4)))} : forvar39);
                      reg130 <= reg8[(3'h7):(1'h1)];
                    end
                end
              if (($unsigned((|(&reg123))) ^ forvar43))
                begin
                  if ($signed(((~|forvar62[(1'h0):(1'h0)]) ?
                      (~|(^reg123)) : $signed(reg31[(3'h7):(3'h6)]))))
                    begin
                      reg131 <= forvar96[(4'h9):(2'h2)];
                      reg132 <= (~|(&reg109[(2'h2):(1'h1)]));
                      reg133 <= ((8'hb1) ?
                          $signed($signed((forvar89 ?
                              forvar40 : reg67))) : {$unsigned(reg86)});
                      reg134 <= ($signed(((reg77 ? forvar89 : reg103) ?
                              $signed(reg102) : $signed((8'h9f)))) ?
                          $signed(($unsigned(reg47) ?
                              {reg72} : $signed((8'hac)))) : reg30);
                    end
                  else
                    begin
                      reg131 <= $signed((~^(~$signed((8'ha1)))));
                      reg132 <= forvar26[(1'h0):(1'h0)];
                      reg133 <= reg53[(1'h1):(1'h1)];
                    end
                  for (forvar135 = (1'h0); (forvar135 < (2'h3)); forvar135 = (forvar135 + (1'h1)))
                    begin
                      reg136 <= reg20[(3'h6):(1'h0)];
                      reg137 <= (-$unsigned(($unsigned((8'ha0)) - $signed(reg133))));
                      reg138 <= (8'hb5);
                      reg139 <= $signed($unsigned((^~forvar113[(3'h6):(3'h4)])));
                    end
                  for (forvar140 = (1'h0); (forvar140 < (2'h3)); forvar140 = (forvar140 + (1'h1)))
                    begin
                      reg141 <= (({$signed(forvar6)} != ((~(8'hb4)) ?
                              $signed(forvar135) : (reg121 ?
                                  (8'hb4) : reg36))) ?
                          reg47 : $signed(forvar16[(3'h6):(2'h3)]));
                      reg142 <= reg70[(4'h8):(3'h4)];
                      reg143 <= forvar113;
                    end
                  reg144 <= ((^(+(|(8'h9f)))) ?
                      (((8'ha2) ? {(8'ha8)} : forvar98[(2'h2):(1'h1)]) ?
                          {(!reg47)} : {$unsigned(forvar76)}) : {(~|reg129)});
                end
              else
                begin
                  if ($unsigned($signed((|(8'h9e)))))
                    begin
                      reg131 <= $unsigned((($signed((8'ha2)) ?
                          (~^reg81) : reg26) ^ {{reg102}}));
                      reg132 <= (^reg67[(3'h4):(1'h0)]);
                      reg133 <= $unsigned($unsigned($unsigned((8'hb2))));
                    end
                  else
                    begin
                      reg131 <= ({reg104} ?
                          $unsigned($unsigned($signed(forvar6))) : reg121);
                      reg132 <= {($signed(reg63) ?
                              (reg116[(4'h8):(1'h1)] ^~ $signed(reg87)) : reg120)};
                      reg133 <= (^$unsigned(($unsigned(forvar19) ?
                          (8'ha7) : reg32[(3'h5):(3'h5)])));
                    end
                  if (reg103[(4'h9):(1'h0)])
                    begin
                      reg134 <= ($signed((~^reg73[(1'h0):(1'h0)])) < forvar11[(3'h6):(2'h2)]);
                      reg135 <= forvar14[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg134 <= ((8'hb6) || {$signed((reg138 ?
                              (8'ha7) : reg74))});
                      reg135 <= forvar88;
                      reg136 <= (forvar14[(2'h3):(1'h1)] >> (~&$unsigned(reg39[(1'h0):(1'h0)])));
                    end
                end
              for (forvar145 = (1'h0); (forvar145 < (1'h0)); forvar145 = (forvar145 + (1'h1)))
                begin
                  if ($signed($signed(reg87[(4'hc):(1'h0)])))
                    begin
                      reg146 <= (reg122 < $signed(reg28));
                      reg147 <= reg24[(2'h2):(1'h1)];
                      reg148 <= $signed($signed($signed((reg128 < forvar27))));
                      reg149 <= {({(reg77 && reg132)} ?
                              $unsigned($unsigned(reg132)) : (reg128[(3'h4):(2'h2)] >> $unsigned(reg115)))};
                    end
                  else
                    begin
                      reg146 <= reg126;
                      reg147 <= $unsigned($signed((&$unsigned(reg44))));
                      reg148 <= ((~&((|reg63) ?
                          (reg75 << reg12) : $unsigned(reg92))) + (^$unsigned($unsigned((8'hba)))));
                      reg149 <= (!(8'hac));
                    end
                  for (forvar150 = (1'h0); (forvar150 < (2'h2)); forvar150 = (forvar150 + (1'h1)))
                    begin
                      reg151 <= reg109[(2'h3):(2'h2)];
                      reg152 <= (|(~&$unsigned(reg63[(2'h3):(1'h0)])));
                      reg153 <= $signed($unsigned((reg10[(2'h2):(2'h2)] & (8'h9d))));
                    end
                  if ({reg80[(1'h1):(1'h0)]})
                    begin
                      reg154 <= (forvar77[(1'h1):(1'h0)] >= ($signed((forvar124 ^ (8'ha6))) ?
                          $unsigned($signed((8'ha6))) : (~$signed(reg129))));
                    end
                  else
                    begin
                      reg154 <= reg117;
                      reg155 <= ($signed($signed((forvar140 ?
                              reg35 : (8'hb0)))) ?
                          forvar114[(2'h3):(1'h0)] : (reg122[(4'hd):(3'h5)] ?
                              forvar59 : ($unsigned(wire3) && (!forvar41))));
                      reg156 <= {(^reg71[(1'h0):(1'h0)])};
                    end
                  reg157 <= $signed({$signed({reg100})});
                end
            end
        end
      if (($signed($unsigned((|reg80))) ?
          wire4[(2'h2):(2'h2)] : (|(&(^~forvar39)))))
        begin
          if (($unsigned(((reg136 ^ reg117) ?
              (~(8'ha2)) : (reg151 != reg13))) >> $signed((|reg38[(1'h0):(1'h0)]))))
            begin
              for (forvar158 = (1'h0); (forvar158 < (1'h0)); forvar158 = (forvar158 + (1'h1)))
                begin
                  if ((~&($unsigned($unsigned(reg31)) <= forvar113[(4'ha):(4'h8)])))
                    begin
                      reg159 <= (wire3[(4'ha):(1'h0)] == (|((reg28 * reg15) ^~ (reg41 ?
                          reg149 : reg137))));
                      reg160 <= $unsigned(forvar21);
                      reg161 <= $unsigned(forvar69[(4'ha):(4'h9)]);
                    end
                  else
                    begin
                      reg159 <= {forvar50};
                      reg160 <= {(reg157 ?
                              reg94 : ((forvar76 << forvar88) ?
                                  reg98[(2'h3):(2'h3)] : (reg48 ?
                                      forvar11 : reg159)))};
                      reg161 <= {(|(reg33 >> $unsigned(reg121)))};
                    end
                end
              if ((8'h9c))
                begin
                  for (forvar162 = (1'h0); (forvar162 < (2'h3)); forvar162 = (forvar162 + (1'h1)))
                    begin
                      reg163 <= $signed((+(|(reg34 ? reg136 : forvar60))));
                      reg164 <= (((reg156 ^~ forvar88[(3'h5):(1'h0)]) ?
                              (~^reg106[(3'h4):(1'h0)]) : $signed($unsigned(reg109))) ?
                          $signed(reg35[(3'h6):(1'h0)]) : ($signed({forvar145}) | $unsigned((forvar113 ?
                              reg12 : (8'hab)))));
                      reg165 <= forvar96[(4'h9):(3'h6)];
                      reg166 <= forvar77[(3'h4):(2'h2)];
                    end
                  for (forvar167 = (1'h0); (forvar167 < (1'h1)); forvar167 = (forvar167 + (1'h1)))
                    begin
                      reg168 <= $unsigned((($unsigned((8'hb6)) >>> forvar107) ?
                          ((~&reg106) << reg23[(3'h6):(1'h0)]) : $unsigned($unsigned(reg154))));
                    end
                end
              else
                begin
                  if ((($signed((-reg58)) ?
                      ({forvar135} ?
                          (!forvar124) : $unsigned(reg8)) : $signed(wire1)) <<< (forvar62[(3'h4):(2'h3)] >= $unsigned(forvar119))))
                    begin
                      reg162 <= (((~|(~reg105)) == (forvar158 & ((8'ha2) ?
                          reg128 : reg71))) == ((reg94[(4'h9):(4'h8)] - $unsigned(reg13)) + ((forvar36 ?
                          (8'ha4) : reg84) + $unsigned(reg70))));
                      reg163 <= $signed($unsigned(reg34[(4'h8):(2'h3)]));
                    end
                  else
                    begin
                      reg162 <= $unsigned(reg132);
                    end
                  if ($unsigned(($unsigned(reg151) != (8'ha7))))
                    begin
                      reg164 <= (8'hb1);
                      reg165 <= (~(reg52 & $unsigned({reg15})));
                      reg166 <= ({($unsigned(reg15) ?
                                  $unsigned(reg79) : reg15[(4'h9):(4'h9)])} ?
                          $unsigned(reg53) : forvar51);
                    end
                  else
                    begin
                      reg164 <= ((forvar6[(2'h2):(1'h1)] ?
                          (reg83 + (|reg11)) : (~(8'hb7))) <<< $signed($unsigned($unsigned(forvar89))));
                    end
                end
            end
          else
            begin
              for (forvar158 = (1'h0); (forvar158 < (2'h2)); forvar158 = (forvar158 + (1'h1)))
                begin
                  for (forvar159 = (1'h0); (forvar159 < (2'h2)); forvar159 = (forvar159 + (1'h1)))
                    begin
                      reg160 <= (reg54[(2'h3):(2'h2)] <<< ((|reg155[(1'h0):(1'h0)]) ?
                          ($signed(forvar159) ?
                              reg152 : (+reg109)) : {wire1[(4'he):(4'he)]}));
                      reg161 <= ((^((reg87 ? reg14 : forvar124) ?
                          $signed(reg20) : (&reg19))) & ((reg12 ?
                              $unsigned(reg41) : {reg27}) ?
                          {$unsigned(forvar36)} : {{forvar27}}));
                    end
                end
              for (forvar162 = (1'h0); (forvar162 < (1'h0)); forvar162 = (forvar162 + (1'h1)))
                begin
                  for (forvar163 = (1'h0); (forvar163 < (1'h1)); forvar163 = (forvar163 + (1'h1)))
                    begin
                      reg164 <= $unsigned(forvar49);
                      reg165 <= $signed((~$unsigned({forvar88})));
                    end
                  for (forvar166 = (1'h0); (forvar166 < (1'h1)); forvar166 = (forvar166 + (1'h1)))
                    begin
                      reg167 <= ((+(!$signed(reg53))) ?
                          (reg56 ?
                              (~(~^(8'ha3))) : (reg75 ?
                                  reg44[(4'h9):(3'h5)] : (&reg84))) : forvar57[(3'h6):(3'h5)]);
                      reg168 <= ($unsigned(reg41[(1'h1):(1'h0)]) ?
                          $signed($signed($signed(reg24))) : {$signed(reg68[(2'h2):(2'h2)])});
                      reg169 <= {reg157[(2'h2):(2'h2)]};
                    end
                  for (forvar170 = (1'h0); (forvar170 < (2'h2)); forvar170 = (forvar170 + (1'h1)))
                    begin
                      reg171 <= (reg23[(1'h1):(1'h1)] > (~&{reg42}));
                      reg172 <= $unsigned((((reg73 ? forvar159 : reg137) ?
                              $unsigned(reg60) : (reg74 ^ forvar49)) ?
                          $signed((forvar51 ? reg32 : (8'hae))) : (~|(8'ha0))));
                    end
                end
            end
        end
      else
        begin
          if ($signed((~^$unsigned(reg157))))
            begin
              for (forvar158 = (1'h0); (forvar158 < (1'h0)); forvar158 = (forvar158 + (1'h1)))
                begin
                  for (forvar159 = (1'h0); (forvar159 < (1'h0)); forvar159 = (forvar159 + (1'h1)))
                    begin
                      reg160 <= (({(reg143 ?
                              reg148 : forvar51)} && (!$unsigned(reg142))) >= forvar150[(2'h3):(2'h2)]);
                      reg161 <= $unsigned(($signed(((8'hb3) ?
                              reg67 : (8'hb7))) ?
                          reg35 : $unsigned(forvar41)));
                      reg162 <= {(reg117 ? forvar163 : reg79)};
                      reg163 <= ($unsigned({reg51}) << forvar30);
                    end
                end
              reg164 <= ($unsigned({$signed(reg152)}) ?
                  reg151[(2'h3):(1'h1)] : $signed(forvar9[(2'h3):(1'h0)]));
              for (forvar165 = (1'h0); (forvar165 < (2'h2)); forvar165 = (forvar165 + (1'h1)))
                begin
                  reg166 <= $unsigned(reg34);
                  for (forvar167 = (1'h0); (forvar167 < (2'h3)); forvar167 = (forvar167 + (1'h1)))
                    begin
                      reg168 <= wire1;
                    end
                end
            end
          else
            begin
              for (forvar158 = (1'h0); (forvar158 < (2'h2)); forvar158 = (forvar158 + (1'h1)))
                begin
                  if ($unsigned(((~&((8'ha4) == reg55)) <<< reg103[(3'h7):(1'h0)])))
                    begin
                      reg159 <= ((~&{(reg132 + reg118)}) | reg38);
                      reg160 <= reg76;
                      reg161 <= reg9;
                    end
                  else
                    begin
                      reg159 <= ((^~reg130[(1'h0):(1'h0)]) ?
                          $signed((!$signed(reg31))) : (($unsigned(reg102) ?
                              $signed(forvar88) : (~^wire0)) ~^ $signed($unsigned(reg72))));
                    end
                  for (forvar162 = (1'h0); (forvar162 < (2'h3)); forvar162 = (forvar162 + (1'h1)))
                    begin
                      reg163 <= $unsigned((&($signed(reg102) ?
                          forvar43 : (reg27 ? forvar18 : reg169))));
                      reg164 <= (($signed((forvar102 * reg53)) | reg28[(2'h2):(1'h1)]) && ($unsigned(reg28) ^ (&$signed((8'hb9)))));
                      reg165 <= ({{forvar119[(1'h1):(1'h1)]}} * (+reg160));
                      reg166 <= ($signed((|(^forvar135))) < (8'hb4));
                    end
                end
              for (forvar167 = (1'h0); (forvar167 < (2'h2)); forvar167 = (forvar167 + (1'h1)))
                begin
                  if ($unsigned($unsigned(({forvar112} ?
                      {reg73} : $signed(reg153)))))
                    begin
                      reg168 <= (8'hb0);
                      reg169 <= reg16;
                    end
                  else
                    begin
                      reg168 <= $unsigned((~|reg124));
                      reg169 <= reg38;
                    end
                  reg170 <= $signed($signed($unsigned($unsigned(reg161))));
                  if ((((8'hb9) ^~ reg172[(1'h1):(1'h0)]) + forvar165))
                    begin
                      reg171 <= ((((^forvar107) | (reg171 | reg171)) ?
                              reg139 : {reg170}) ?
                          $unsigned($unsigned($signed(forvar162))) : (|{$unsigned((8'had))}));
                      reg172 <= ($signed($unsigned(reg143[(3'h7):(3'h6)])) ?
                          reg157 : (!((reg75 ? reg167 : reg122) << reg156)));
                    end
                  else
                    begin
                      reg171 <= (($signed(reg85) ?
                              $unsigned($unsigned((8'ha9))) : forvar102[(3'h6):(2'h2)]) ?
                          $signed(forvar124[(1'h0):(1'h0)]) : ($unsigned(forvar6[(4'hb):(3'h6)]) ?
                              $signed({wire3}) : ((~^forvar59) ?
                                  $signed((8'hba)) : (+reg103))));
                      reg172 <= reg7[(1'h1):(1'h1)];
                      reg173 <= (((~&(&forvar51)) - (^(8'haa))) ?
                          (($signed(forvar46) ?
                                  ((8'ha8) ?
                                      (8'haa) : forvar60) : ((8'hba) - (8'hac))) ?
                              $unsigned($unsigned(reg143)) : reg91[(2'h2):(1'h0)]) : ((~|(forvar83 ?
                                  (8'ha4) : reg122)) ?
                              (+$signed(reg97)) : {$unsigned(reg126)}));
                      reg174 <= ((reg21 ^~ ({reg78} ?
                          reg164[(4'h8):(2'h3)] : (-reg26))) == forvar165[(4'he):(4'h8)]);
                    end
                  for (forvar175 = (1'h0); (forvar175 < (2'h3)); forvar175 = (forvar175 + (1'h1)))
                    begin
                      reg176 <= $signed((((^reg81) < (forvar166 ?
                          reg128 : (8'haf))) && $unsigned((reg169 != reg147))));
                      reg177 <= $signed(($unsigned((^(8'ha2))) ?
                          ($signed(reg144) + forvar44) : ($unsigned(reg122) ?
                              (^forvar7) : (reg70 ? reg9 : reg130))));
                      reg178 <= $unsigned((reg67[(3'h4):(1'h0)] ?
                          $unsigned((forvar83 ~^ reg56)) : reg174[(3'h5):(1'h0)]));
                    end
                end
              for (forvar179 = (1'h0); (forvar179 < (1'h1)); forvar179 = (forvar179 + (1'h1)))
                begin
                  for (forvar180 = (1'h0); (forvar180 < (2'h3)); forvar180 = (forvar180 + (1'h1)))
                    begin
                      reg181 <= reg6;
                    end
                  if ($signed((forvar180 ?
                      reg144[(2'h3):(2'h2)] : $unsigned((+forvar75)))))
                    begin
                      reg182 <= ((^~(-$unsigned(reg44))) ?
                          wire5[(1'h0):(1'h0)] : (8'hb6));
                      reg183 <= reg143;
                    end
                  else
                    begin
                      reg182 <= reg152[(3'h4):(3'h4)];
                      reg183 <= (!(!reg94[(4'h8):(3'h4)]));
                    end
                  for (forvar184 = (1'h0); (forvar184 < (1'h1)); forvar184 = (forvar184 + (1'h1)))
                    begin
                      reg185 <= (({(reg120 ^~ reg181)} != (&forvar167[(1'h0):(1'h0)])) ?
                          (($signed(wire5) >= (-reg53)) ?
                              $signed((reg29 ?
                                  reg63 : reg72)) : reg111) : $unsigned(reg76[(3'h4):(2'h2)]));
                      reg186 <= ((reg182[(3'h6):(3'h4)] ?
                              ($unsigned(forvar163) + reg94) : reg92) ?
                          (8'h9e) : $signed((reg34 ~^ $signed(reg48))));
                    end
                  if ((reg157[(2'h2):(1'h0)] ^ ((+$unsigned((8'hb0))) ?
                      $signed((reg141 ?
                          reg162 : reg29)) : reg79[(3'h4):(2'h2)])))
                    begin
                      reg187 <= reg91;
                    end
                  else
                    begin
                      reg187 <= $signed(reg36[(3'h6):(2'h2)]);
                      reg188 <= reg66;
                    end
                end
              for (forvar189 = (1'h0); (forvar189 < (2'h3)); forvar189 = (forvar189 + (1'h1)))
                begin
                  for (forvar190 = (1'h0); (forvar190 < (1'h1)); forvar190 = (forvar190 + (1'h1)))
                    begin
                      reg191 <= forvar140[(2'h3):(1'h1)];
                    end
                  for (forvar192 = (1'h0); (forvar192 < (2'h3)); forvar192 = (forvar192 + (1'h1)))
                    begin
                      reg193 <= (~|$unsigned(reg91[(3'h6):(3'h4)]));
                      reg194 <= (!reg11[(3'h4):(2'h2)]);
                      reg195 <= (|wire1[(4'he):(4'ha)]);
                    end
                end
            end
          if ((~|$unsigned($signed({reg40}))))
            begin
              for (forvar196 = (1'h0); (forvar196 < (2'h2)); forvar196 = (forvar196 + (1'h1)))
                begin
                  if ($unsigned(($unsigned((forvar135 ?
                      (8'h9e) : reg149)) > (reg108[(3'h5):(1'h1)] < reg160[(2'h2):(1'h0)]))))
                    begin
                      reg197 <= $signed((~&(reg129 ?
                          (reg162 ? reg121 : reg105) : $unsigned(reg30))));
                    end
                  else
                    begin
                      reg197 <= forvar9;
                    end
                  if ((8'hac))
                    begin
                      reg198 <= ((!reg151[(2'h2):(1'h0)]) * $unsigned(forvar51));
                      reg199 <= (-(8'hb0));
                      reg200 <= {(|{$signed(reg44)})};
                    end
                  else
                    begin
                      reg198 <= reg147[(1'h0):(1'h0)];
                    end
                  reg201 <= (reg71[(1'h0):(1'h0)] <= reg81[(4'h8):(3'h4)]);
                end
            end
          else
            begin
              if ($signed((+$signed((~^reg32)))))
                begin
                  for (forvar196 = (1'h0); (forvar196 < (1'h1)); forvar196 = (forvar196 + (1'h1)))
                    begin
                      reg197 <= reg35[(1'h0):(1'h0)];
                      reg198 <= {$signed(((reg71 >> reg24) ? {wire0} : reg77))};
                      reg199 <= ((forvar44[(4'h9):(3'h7)] && $signed((8'h9d))) ?
                          (~&(forvar83 || ((8'ha2) >>> reg164))) : $signed(forvar16[(1'h1):(1'h1)]));
                      reg200 <= (!$unsigned(((~^forvar9) + $unsigned(forvar30))));
                    end
                  for (forvar201 = (1'h0); (forvar201 < (2'h2)); forvar201 = (forvar201 + (1'h1)))
                    begin
                      reg202 <= $signed(reg127[(3'h6):(2'h2)]);
                      reg203 <= ((forvar36[(4'hf):(4'h8)] * (!((8'ha5) ?
                          reg198 : reg83))) & forvar201);
                    end
                end
              else
                begin
                  for (forvar196 = (1'h0); (forvar196 < (2'h2)); forvar196 = (forvar196 + (1'h1)))
                    begin
                      reg197 <= forvar46[(2'h2):(1'h0)];
                      reg198 <= (^~reg193[(2'h3):(1'h0)]);
                      reg199 <= $signed((forvar77[(4'h8):(4'h8)] & (reg183 ?
                          reg34[(3'h5):(1'h1)] : (~|reg87))));
                      reg200 <= $unsigned((!$signed((reg177 ^ reg135))));
                    end
                  if (((((reg155 ? reg48 : reg149) ?
                          $unsigned(forvar98) : reg37[(4'h8):(3'h4)]) ?
                      $unsigned({reg52}) : $unsigned((8'ha5))) * ($unsigned((reg39 ?
                          reg98 : reg8)) ?
                      {reg27[(1'h0):(1'h0)]} : (~|(&reg57)))))
                    begin
                      reg201 <= reg29;
                      reg202 <= ((+((|reg72) || (forvar114 ? reg29 : reg136))) ?
                          {{$unsigned(forvar159)}} : $signed({reg135}));
                    end
                  else
                    begin
                      reg201 <= (((&reg159[(2'h2):(2'h2)]) ~^ reg44[(4'hd):(2'h2)]) < reg127);
                      reg202 <= ($signed(((forvar190 ?
                          reg59 : reg88) && (^reg23))) > {reg161});
                      reg203 <= $signed({(~(reg104 <<< forvar175))});
                      reg204 <= reg87;
                    end
                end
            end
          if ($unsigned((reg110 << {{reg200}})))
            begin
              for (forvar205 = (1'h0); (forvar205 < (1'h0)); forvar205 = (forvar205 + (1'h1)))
                begin
                  if (forvar40)
                    begin
                      reg206 <= (($unsigned((8'hb4)) ?
                          reg198[(2'h3):(1'h1)] : (reg36[(4'h8):(4'h8)] ?
                              forvar43[(2'h2):(1'h1)] : ((8'h9e) ^~ forvar166))) || ((|reg59[(1'h0):(1'h0)]) ?
                          reg135 : $signed(forvar16[(2'h3):(2'h2)])));
                      reg207 <= {(+forvar150)};
                      reg208 <= ($unsigned(((forvar107 << reg33) * (&forvar102))) * ((forvar162[(4'h8):(1'h0)] ?
                          {reg123} : $unsigned(reg163)) | ((forvar165 & reg57) >= {reg73})));
                    end
                  else
                    begin
                      reg206 <= ($unsigned(reg194) ?
                          (~^(^~$signed(reg121))) : ((!$signed(reg136)) + (reg124 != $signed(reg37))));
                    end
                  for (forvar209 = (1'h0); (forvar209 < (2'h2)); forvar209 = (forvar209 + (1'h1)))
                    begin
                      reg210 <= ($unsigned({(-(8'hb6))}) - {forvar69[(3'h7):(2'h3)]});
                      reg211 <= $signed($signed($signed(reg157[(1'h0):(1'h0)])));
                      reg212 <= (-(forvar98 ? reg32 : $unsigned(reg188)));
                      reg213 <= (^$signed(wire3));
                    end
                  if (reg185[(4'ha):(3'h7)])
                    begin
                      reg214 <= {reg101[(2'h2):(1'h0)]};
                      reg215 <= $unsigned((8'haa));
                    end
                  else
                    begin
                      reg214 <= $unsigned(reg74);
                      reg215 <= $unsigned(forvar9);
                      reg216 <= (~forvar7);
                    end
                  for (forvar217 = (1'h0); (forvar217 < (2'h3)); forvar217 = (forvar217 + (1'h1)))
                    begin
                      reg218 <= reg207[(1'h0):(1'h0)];
                      reg219 <= $unsigned(forvar119);
                    end
                end
            end
          else
            begin
              for (forvar205 = (1'h0); (forvar205 < (1'h0)); forvar205 = (forvar205 + (1'h1)))
                begin
                  if (forvar114)
                    begin
                      reg206 <= (((|{reg26}) ?
                          $signed((reg10 ~^ reg195)) : reg176[(2'h2):(1'h1)]) * {reg186});
                      reg207 <= forvar73[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg206 <= reg73[(3'h4):(2'h2)];
                    end
                  for (forvar208 = (1'h0); (forvar208 < (2'h2)); forvar208 = (forvar208 + (1'h1)))
                    begin
                      reg209 <= reg202;
                      reg210 <= (8'ha2);
                    end
                  for (forvar211 = (1'h0); (forvar211 < (1'h1)); forvar211 = (forvar211 + (1'h1)))
                    begin
                      reg212 <= $signed(forvar107);
                      reg213 <= forvar88;
                    end
                  reg214 <= ($unsigned((~^$unsigned(forvar83))) ?
                      reg30[(1'h0):(1'h0)] : (|((wire1 || forvar27) ^ (8'hb9))));
                end
            end
        end
      for (forvar220 = (1'h0); (forvar220 < (1'h1)); forvar220 = (forvar220 + (1'h1)))
        begin
          if (((({(8'ha7)} ? forvar6 : (reg87 == (8'h9c))) ?
                  $unsigned($unsigned((8'haa))) : $signed(forvar57)) ?
              $signed(((reg90 ? reg80 : reg201) ?
                  (reg10 ?
                      reg132 : reg37) : $unsigned((8'hb7)))) : {((reg76 + reg219) ?
                      reg85 : ((8'haf) >>> reg81))}))
            begin
              if ($unsigned($signed((((8'hac) >>> reg210) ~^ $signed(reg130)))))
                begin
                  for (forvar221 = (1'h0); (forvar221 < (2'h2)); forvar221 = (forvar221 + (1'h1)))
                    begin
                      reg222 <= $unsigned((+((+reg56) ?
                          ((8'ha4) || (8'ha4)) : reg136)));
                    end
                end
              else
                begin
                  if (reg137)
                    begin
                      reg221 <= $unsigned(($signed({reg12}) ?
                          reg151[(2'h3):(1'h1)] : $signed({reg88})));
                    end
                  else
                    begin
                      reg221 <= ({reg100} ?
                          $unsigned(($signed(forvar175) + $unsigned(reg171))) : (~&(~$signed((8'hb9)))));
                    end
                  if ($signed(reg95[(2'h3):(1'h0)]))
                    begin
                      reg222 <= forvar114[(2'h3):(1'h1)];
                      reg223 <= $unsigned($unsigned((8'ha1)));
                      reg224 <= (reg111[(4'hd):(3'h5)] ?
                          $signed(reg66[(3'h4):(1'h0)]) : (^~$unsigned($unsigned(reg208))));
                      reg225 <= (8'hb2);
                    end
                  else
                    begin
                      reg222 <= (reg13[(1'h0):(1'h0)] | (8'h9d));
                    end
                  reg226 <= $unsigned((((-(8'hb9)) ?
                          reg125[(3'h4):(2'h3)] : (~reg10)) ?
                      $signed($signed(reg73)) : (~&{reg33})));
                  reg227 <= {((~&(reg160 ?
                          forvar62 : reg122)) + $unsigned(reg79[(2'h3):(1'h0)]))};
                end
              for (forvar228 = (1'h0); (forvar228 < (2'h3)); forvar228 = (forvar228 + (1'h1)))
                begin
                  for (forvar229 = (1'h0); (forvar229 < (1'h0)); forvar229 = (forvar229 + (1'h1)))
                    begin
                      reg230 <= $signed($unsigned(reg198[(2'h2):(2'h2)]));
                      reg231 <= wire1;
                      reg232 <= ({$unsigned(reg95[(4'ha):(1'h0)])} | (forvar69[(3'h4):(3'h4)] < ((!forvar16) ?
                          (forvar73 ?
                              reg146 : (8'hab)) : forvar88[(3'h5):(1'h1)])));
                      reg233 <= ({((~|forvar119) <<< (^~forvar83))} ?
                          ({$unsigned((8'hac))} <= (((8'ha5) > (8'hb3)) ~^ (reg183 ?
                              reg161 : reg170))) : reg206[(3'h4):(1'h0)]);
                    end
                  reg234 <= $unsigned($unsigned((((8'hab) >= reg215) | (8'ha0))));
                  if ({$signed(forvar175)})
                    begin
                      reg235 <= forvar221;
                      reg236 <= reg167;
                      reg237 <= reg133;
                    end
                  else
                    begin
                      reg235 <= (+$unsigned(({forvar88} ~^ $unsigned(reg208))));
                    end
                end
              reg238 <= $signed(((~|(8'ha5)) ?
                  ($unsigned(reg212) ?
                      (forvar220 - reg44) : forvar43) : $unsigned($signed(forvar15))));
            end
          else
            begin
              for (forvar221 = (1'h0); (forvar221 < (2'h2)); forvar221 = (forvar221 + (1'h1)))
                begin
                  for (forvar222 = (1'h0); (forvar222 < (2'h2)); forvar222 = (forvar222 + (1'h1)))
                    begin
                      reg223 <= ((-$signed({reg118})) ?
                          (^$signed(forvar44)) : $unsigned($signed(reg146)));
                    end
                  for (forvar224 = (1'h0); (forvar224 < (2'h3)); forvar224 = (forvar224 + (1'h1)))
                    begin
                      reg225 <= $unsigned($signed((forvar73[(2'h2):(1'h0)] ^~ reg73[(1'h0):(1'h0)])));
                    end
                  if ({((^~(~^reg22)) ^ (reg22 ^ (reg163 ?
                          forvar69 : reg161)))})
                    begin
                      reg226 <= ({$unsigned((reg178 ?
                              reg135 : reg110))} >>> reg149);
                      reg227 <= reg10[(1'h1):(1'h0)];
                      reg228 <= {(^{(reg63 || reg33)})};
                      reg229 <= reg101[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg226 <= reg168;
                      reg227 <= ($signed(forvar140[(4'h9):(2'h3)]) || reg160);
                    end
                  if ({$signed($unsigned(reg153[(3'h5):(2'h2)]))})
                    begin
                      reg230 <= reg228[(1'h0):(1'h0)];
                      reg231 <= $signed((~^forvar62));
                      reg232 <= ($unsigned($unsigned((^reg149))) ?
                          reg51 : $unsigned(reg218[(4'hd):(4'hd)]));
                      reg233 <= ($signed(reg141) ?
                          ($signed((~^reg185)) ~^ (forvar31[(1'h0):(1'h0)] != (!reg32))) : ($signed((reg93 + wire4)) << reg208));
                    end
                  else
                    begin
                      reg230 <= reg39[(3'h5):(2'h2)];
                      reg231 <= $unsigned(reg38[(3'h5):(1'h0)]);
                      reg232 <= forvar69[(2'h2):(2'h2)];
                    end
                end
            end
        end
    end
  assign wire239 = ($unsigned((~(&reg156))) ?
                       reg75 : (({reg229} >>> (8'ha0)) ?
                           reg123 : $signed((~|reg72))));
  assign wire240 = ((~&({reg138} | $signed(reg74))) ?
                       ($signed((reg66 <<< (8'hb5))) ?
                           $unsigned((8'ha7)) : reg95[(3'h7):(1'h1)]) : (reg142[(4'hb):(3'h5)] ?
                           {(reg32 ^ (8'hb6))} : $unsigned(((8'ha5) && reg138))));
  always
    @(posedge clk) begin
      if (reg226[(2'h2):(1'h0)])
        begin
          if ({(^$unsigned($signed(reg61)))})
            begin
              reg241 <= $unsigned(reg31[(2'h3):(2'h2)]);
              for (forvar242 = (1'h0); (forvar242 < (2'h2)); forvar242 = (forvar242 + (1'h1)))
                begin
                  for (forvar243 = (1'h0); (forvar243 < (2'h2)); forvar243 = (forvar243 + (1'h1)))
                    begin
                      reg244 <= (8'ha7);
                      reg245 <= ((reg95[(3'h4):(2'h3)] ?
                              reg19[(3'h6):(1'h1)] : $unsigned(wire3[(4'h9):(3'h4)])) ?
                          (($unsigned((8'had)) + ((8'ha8) ?
                              (8'h9e) : reg85)) << {reg215}) : $signed(reg101[(3'h5):(2'h2)]));
                    end
                  if (reg155[(2'h2):(1'h0)])
                    begin
                      reg246 <= ((+$unsigned(reg76[(2'h2):(1'h0)])) ?
                          (((reg193 ? reg183 : reg155) ?
                              (reg153 || reg146) : (~^reg183)) >>> (~(+reg164))) : ({$signed(reg100)} ?
                              reg31 : (~((8'had) == reg92))));
                    end
                  else
                    begin
                      reg246 <= reg95;
                      reg247 <= (|(+(((8'hb1) ? reg195 : reg185) != reg15)));
                      reg248 <= $unsigned({$signed(reg36[(2'h2):(2'h2)])});
                      reg249 <= (((~$unsigned(reg222)) ?
                          $signed((8'h9c)) : (reg31[(3'h7):(3'h7)] >= $unsigned(reg203))) ^ $signed(reg58));
                    end
                  for (forvar250 = (1'h0); (forvar250 < (2'h3)); forvar250 = (forvar250 + (1'h1)))
                    begin
                      reg251 <= $signed($signed(((reg156 <<< reg17) ?
                          reg12 : $signed(forvar243))));
                    end
                  for (forvar252 = (1'h0); (forvar252 < (2'h2)); forvar252 = (forvar252 + (1'h1)))
                    begin
                      reg253 <= reg136;
                    end
                end
              for (forvar254 = (1'h0); (forvar254 < (1'h0)); forvar254 = (forvar254 + (1'h1)))
                begin
                  reg255 <= {({(~|reg173)} - reg25[(2'h2):(1'h0)])};
                  reg256 <= (reg13[(3'h6):(3'h5)] & (reg21[(2'h2):(2'h2)] ?
                      reg248 : reg133[(2'h3):(2'h2)]));
                  for (forvar257 = (1'h0); (forvar257 < (2'h3)); forvar257 = (forvar257 + (1'h1)))
                    begin
                      reg258 <= {((~&reg70) && $signed($unsigned(reg73)))};
                    end
                  if (reg219[(4'ha):(3'h5)])
                    begin
                      reg259 <= (((!$unsigned(reg39)) << {$signed(reg28)}) ?
                          reg167 : (~^(reg79 ? $unsigned(reg216) : (~|reg33))));
                      reg260 <= reg74;
                      reg261 <= reg72;
                    end
                  else
                    begin
                      reg259 <= (|$signed($unsigned((reg229 ?
                          reg123 : reg228))));
                      reg260 <= $unsigned(reg146[(4'ha):(4'h9)]);
                    end
                end
            end
          else
            begin
              for (forvar241 = (1'h0); (forvar241 < (2'h2)); forvar241 = (forvar241 + (1'h1)))
                begin
                  if (((-$signed(reg195)) ?
                      (!(~^reg88[(4'h9):(3'h4)])) : {$unsigned(((8'hb2) && reg259))}))
                    begin
                      reg242 <= reg253;
                      reg243 <= reg59[(1'h1):(1'h0)];
                      reg244 <= (8'ha0);
                      reg245 <= forvar242;
                    end
                  else
                    begin
                      reg242 <= ((reg85[(1'h0):(1'h0)] == {$unsigned(reg51)}) * (^($signed(reg151) ^ ((8'ha5) ?
                          (8'had) : reg153))));
                      reg243 <= ($unsigned({$signed(reg24)}) ?
                          ((8'hac) || (~{reg23})) : $signed(((^(8'ha6)) ?
                              (reg79 >= reg198) : reg92[(3'h4):(1'h1)])));
                      reg244 <= $unsigned(({$signed(reg209)} < reg141));
                    end
                end
            end
        end
      else
        begin
          for (forvar241 = (1'h0); (forvar241 < (2'h3)); forvar241 = (forvar241 + (1'h1)))
            begin
              if ((^~reg181))
                begin
                  for (forvar242 = (1'h0); (forvar242 < (2'h3)); forvar242 = (forvar242 + (1'h1)))
                    begin
                      reg243 <= $signed((reg203[(2'h2):(1'h1)] ?
                          reg26 : $signed((reg163 ? (8'haf) : reg154))));
                      reg244 <= $signed(((8'hb7) ^~ (-(reg54 ?
                          reg68 : reg165))));
                      reg245 <= reg75[(4'h8):(2'h2)];
                      reg246 <= $signed(((|{reg172}) ^ (reg230 >> reg153[(3'h5):(3'h4)])));
                    end
                  if (((reg37 ? (~^$signed(reg26)) : reg84) >= ((8'hb1) ?
                      ((reg198 ?
                          reg83 : (8'hab)) * {reg79}) : {((8'hae) >>> reg98)})))
                    begin
                      reg247 <= ($signed((+$signed(reg231))) ^ reg55[(3'h4):(3'h4)]);
                      reg248 <= (^~$unsigned(reg238));
                      reg249 <= ((!(^{reg152})) ?
                          reg92[(3'h6):(1'h0)] : (-$unsigned($signed(reg79))));
                      reg250 <= ({(~(^~reg82))} ^~ (reg27 - (8'hb5)));
                    end
                  else
                    begin
                      reg247 <= {(reg222[(3'h4):(1'h1)] < (reg58 <= {reg131}))};
                      reg248 <= ({reg101[(1'h1):(1'h1)]} ?
                          reg206[(3'h5):(1'h1)] : $signed(($signed(reg169) < $unsigned((8'hb4)))));
                      reg249 <= {($signed({reg47}) ^ (8'ha9))};
                      reg250 <= ($unsigned(($signed(reg197) ?
                              (reg91 <= reg6) : $signed(reg128))) ?
                          $signed(($unsigned(reg31) <= reg7)) : ((~^(reg39 < reg261)) ?
                              reg224 : (8'had)));
                    end
                  if (reg186)
                    begin
                      reg251 <= reg26[(4'ha):(3'h5)];
                      reg252 <= $unsigned(((^~reg30[(1'h1):(1'h1)]) ?
                          (~$signed((8'hb8))) : forvar250));
                      reg253 <= reg57;
                    end
                  else
                    begin
                      reg251 <= $signed($signed(((reg187 ? (8'ha1) : reg40) ?
                          (~&reg166) : reg110[(3'h4):(3'h4)])));
                    end
                end
              else
                begin
                  reg242 <= ($unsigned(((8'h9d) && (reg244 >> reg187))) ^ {$signed((reg72 * reg23))});
                end
            end
        end
      if ({(reg172[(3'h5):(3'h4)] ?
              reg22[(3'h5):(2'h3)] : $unsigned($unsigned(reg183)))})
        begin
          if (reg234[(1'h0):(1'h0)])
            begin
              for (forvar262 = (1'h0); (forvar262 < (2'h3)); forvar262 = (forvar262 + (1'h1)))
                begin
                  for (forvar263 = (1'h0); (forvar263 < (1'h0)); forvar263 = (forvar263 + (1'h1)))
                    begin
                      reg264 <= $signed({reg223[(1'h0):(1'h0)]});
                      reg265 <= (reg79 ?
                          reg131 : $unsigned((+$signed(forvar254))));
                      reg266 <= $unsigned($signed($signed(forvar262)));
                    end
                end
              for (forvar267 = (1'h0); (forvar267 < (1'h1)); forvar267 = (forvar267 + (1'h1)))
                begin
                  for (forvar268 = (1'h0); (forvar268 < (2'h2)); forvar268 = (forvar268 + (1'h1)))
                    begin
                      reg269 <= reg169;
                      reg270 <= (~&reg242);
                      reg271 <= (reg172 ?
                          reg213[(3'h5):(3'h4)] : (~^($signed(reg60) >> reg122)));
                    end
                  for (forvar272 = (1'h0); (forvar272 < (2'h3)); forvar272 = (forvar272 + (1'h1)))
                    begin
                      reg273 <= reg155;
                      reg274 <= (~$signed({(!reg209)}));
                      reg275 <= (((reg265[(3'h7):(1'h1)] && ((8'hb7) ?
                          reg55 : reg210)) == $signed(((8'ha1) != reg144))) != $signed($unsigned(reg166[(4'ha):(4'ha)])));
                      reg276 <= {({(^~(8'h9e))} ?
                              $signed(reg74[(3'h7):(3'h5)]) : $unsigned((~reg247)))};
                    end
                end
              for (forvar277 = (1'h0); (forvar277 < (1'h0)); forvar277 = (forvar277 + (1'h1)))
                begin
                  if (($signed(reg181[(4'ha):(3'h6)]) * $unsigned($signed($signed(reg48)))))
                    begin
                      reg278 <= (~(^~$signed($signed((8'h9f)))));
                      reg279 <= (8'ha5);
                    end
                  else
                    begin
                      reg278 <= reg66[(1'h1):(1'h1)];
                    end
                end
              reg280 <= $unsigned(wire4[(1'h1):(1'h1)]);
            end
          else
            begin
              if (($unsigned(((reg163 <= reg244) ?
                      reg185 : (reg152 ? (8'hb7) : reg213))) ?
                  (&(&reg58)) : reg100))
                begin
                  reg262 <= (8'ha7);
                  for (forvar263 = (1'h0); (forvar263 < (2'h3)); forvar263 = (forvar263 + (1'h1)))
                    begin
                      reg264 <= reg146[(3'h5):(3'h4)];
                      reg265 <= reg168;
                      reg266 <= reg66[(3'h6):(3'h4)];
                      reg267 <= ((($unsigned(reg10) ?
                                  (reg13 ?
                                      (8'ha4) : (8'ha2)) : reg99[(3'h5):(1'h0)]) ?
                              (8'hb9) : ((forvar252 ?
                                  reg51 : reg108) <<< $unsigned(reg226))) ?
                          (8'hb3) : {(~|$unsigned(reg110))});
                    end
                  for (forvar268 = (1'h0); (forvar268 < (1'h1)); forvar268 = (forvar268 + (1'h1)))
                    begin
                      reg269 <= reg235;
                      reg270 <= reg111[(4'h9):(4'h9)];
                      reg271 <= reg261[(4'ha):(4'h9)];
                      reg272 <= ((-$unsigned($unsigned(reg237))) >= reg15[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  reg262 <= ((~^$signed((reg103 && reg58))) && $unsigned($signed($signed(reg213))));
                  if (reg103[(3'h5):(1'h0)])
                    begin
                      reg263 <= reg16[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg263 <= $unsigned((reg244[(3'h4):(3'h4)] ?
                          ({reg24} ?
                              (reg229 ~^ reg79) : (reg275 ?
                                  reg64 : reg269)) : (reg97[(3'h6):(1'h1)] >= $signed(reg78))));
                      reg264 <= {reg101[(2'h3):(2'h2)]};
                      reg265 <= reg73[(2'h3):(1'h0)];
                      reg266 <= reg125;
                    end
                  for (forvar267 = (1'h0); (forvar267 < (1'h1)); forvar267 = (forvar267 + (1'h1)))
                    begin
                      reg268 <= reg256[(1'h0):(1'h0)];
                      reg269 <= (reg242 ?
                          $signed($signed($unsigned(reg97))) : {$signed({reg268})});
                    end
                  for (forvar270 = (1'h0); (forvar270 < (1'h0)); forvar270 = (forvar270 + (1'h1)))
                    begin
                      reg271 <= $unsigned($signed($signed((-reg10))));
                      reg272 <= {($unsigned(reg258[(3'h4):(2'h3)]) ?
                              reg268[(2'h2):(1'h1)] : ((reg161 * reg74) ?
                                  (~&forvar242) : (^(8'ha2))))};
                      reg273 <= $signed($signed(forvar268));
                    end
                end
              for (forvar274 = (1'h0); (forvar274 < (2'h3)); forvar274 = (forvar274 + (1'h1)))
                begin
                  for (forvar275 = (1'h0); (forvar275 < (2'h2)); forvar275 = (forvar275 + (1'h1)))
                    begin
                      reg276 <= $signed(reg159);
                    end
                end
            end
          for (forvar281 = (1'h0); (forvar281 < (2'h3)); forvar281 = (forvar281 + (1'h1)))
            begin
              for (forvar282 = (1'h0); (forvar282 < (2'h3)); forvar282 = (forvar282 + (1'h1)))
                begin
                  if (($unsigned($signed((+(8'ha1)))) ?
                      $signed(reg169) : ((reg88[(4'h9):(2'h3)] ?
                              (^~reg263) : ((8'hba) ^~ reg144)) ?
                          {forvar250} : $unsigned((reg234 ? reg63 : reg143)))))
                    begin
                      reg283 <= (reg261[(4'h8):(1'h1)] || {$signed({reg170})});
                    end
                  else
                    begin
                      reg283 <= reg194;
                      reg284 <= $unsigned($unsigned((^~reg24[(3'h4):(1'h0)])));
                      reg285 <= {$unsigned(((reg275 ?
                              reg58 : reg106) + (reg87 - reg154)))};
                    end
                  if (reg92[(3'h4):(2'h3)])
                    begin
                      reg286 <= ({((reg125 ? reg78 : (8'ha9)) - {wire1})} ?
                          {(^$signed(reg229))} : ($unsigned(reg149) ?
                              $signed((reg128 * reg126)) : ((^~(8'had)) ?
                                  $unsigned(forvar252) : reg120)));
                      reg287 <= forvar263;
                    end
                  else
                    begin
                      reg286 <= ($signed((|(8'ha9))) >>> {reg267});
                      reg287 <= $unsigned($signed(reg31));
                      reg288 <= $unsigned(reg169[(3'h7):(2'h3)]);
                    end
                  for (forvar289 = (1'h0); (forvar289 < (1'h0)); forvar289 = (forvar289 + (1'h1)))
                    begin
                      reg290 <= $signed(reg120);
                      reg291 <= $unsigned((^~forvar242));
                      reg292 <= (((~^(reg153 && reg278)) ?
                          $unsigned(reg75) : ($signed(reg245) ?
                              (!reg81) : reg36[(3'h7):(3'h5)])) && reg171[(3'h7):(1'h1)]);
                    end
                  for (forvar293 = (1'h0); (forvar293 < (1'h0)); forvar293 = (forvar293 + (1'h1)))
                    begin
                      reg294 <= (|(reg285 ?
                          wire2[(2'h3):(2'h3)] : ($signed((8'ha1)) ?
                              reg86 : $signed((8'ha5)))));
                    end
                end
            end
        end
      else
        begin
          for (forvar262 = (1'h0); (forvar262 < (1'h1)); forvar262 = (forvar262 + (1'h1)))
            begin
              if ($signed(($signed((reg93 ? reg32 : reg58)) >> (^~(^~reg17)))))
                begin
                  reg263 <= (^reg88[(4'hc):(3'h7)]);
                  reg264 <= reg66;
                  if (reg42[(2'h2):(2'h2)])
                    begin
                      reg265 <= reg280[(4'he):(4'ha)];
                      reg266 <= $unsigned((8'ha5));
                      reg267 <= (^~$unsigned($unsigned((^~reg199))));
                    end
                  else
                    begin
                      reg265 <= $signed($unsigned($unsigned((reg161 && reg253))));
                      reg266 <= ((^((reg78 ? reg42 : (8'ha1)) ?
                          (8'haf) : (forvar277 ^~ reg75))) && (|forvar270[(3'h4):(2'h3)]));
                    end
                  if (($unsigned($signed($unsigned(reg110))) ?
                      (reg51 >= (+(reg27 - (8'ha7)))) : (~&(8'ha8))))
                    begin
                      reg268 <= (reg130 ?
                          $signed(reg51[(2'h3):(2'h2)]) : reg191[(3'h4):(1'h0)]);
                      reg269 <= (reg81 != reg74);
                      reg270 <= $unsigned((^(|(-reg160))));
                    end
                  else
                    begin
                      reg268 <= (&reg182[(4'h9):(4'h9)]);
                      reg269 <= ({(&(reg61 ? (8'ha7) : wire1))} ?
                          reg210 : (reg16[(3'h5):(2'h2)] >>> $unsigned(reg74[(1'h0):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar263 = (1'h0); (forvar263 < (1'h0)); forvar263 = (forvar263 + (1'h1)))
                    begin
                      reg264 <= reg292;
                      reg265 <= $signed(($unsigned($signed(forvar272)) ^~ $unsigned((reg274 != reg67))));
                      reg266 <= ((reg232 ?
                              $signed({(8'hab)}) : $unsigned($unsigned(reg21))) ?
                          $signed(reg71) : $signed(reg286));
                      reg267 <= reg32[(1'h0):(1'h0)];
                    end
                  for (forvar268 = (1'h0); (forvar268 < (2'h2)); forvar268 = (forvar268 + (1'h1)))
                    begin
                      reg269 <= reg106;
                    end
                  for (forvar270 = (1'h0); (forvar270 < (2'h3)); forvar270 = (forvar270 + (1'h1)))
                    begin
                      reg271 <= {((~&((8'hb4) ? (8'hb5) : reg274)) ?
                              (^$unsigned(reg32)) : (8'hb7))};
                      reg272 <= $unsigned(reg33);
                      reg273 <= ((($signed(reg134) ?
                                  $unsigned(reg181) : (|(8'ha9))) ?
                              $signed($signed(reg42)) : reg258) ?
                          ($signed(((8'hae) <= (8'ha9))) ?
                              $unsigned(reg134) : (^((8'hab) ?
                                  reg40 : reg195))) : reg146);
                    end
                end
              for (forvar274 = (1'h0); (forvar274 < (2'h2)); forvar274 = (forvar274 + (1'h1)))
                begin
                  if ($signed($signed($unsigned($signed(reg57)))))
                    begin
                      reg275 <= (8'h9e);
                      reg276 <= reg159[(3'h4):(3'h4)];
                      reg277 <= $unsigned({(8'hae)});
                      reg278 <= (^~reg231[(4'hc):(4'hb)]);
                    end
                  else
                    begin
                      reg275 <= $signed(($unsigned($signed(reg26)) ?
                          (reg160 - (reg56 >> reg233)) : reg14));
                      reg276 <= reg132[(2'h3):(2'h3)];
                      reg277 <= $unsigned({((reg259 ? reg227 : reg57) ?
                              reg264 : ((8'haf) ? reg207 : reg53))});
                      reg278 <= {reg87};
                    end
                end
              for (forvar279 = (1'h0); (forvar279 < (1'h0)); forvar279 = (forvar279 + (1'h1)))
                begin
                  if (({$unsigned(reg243)} ? {(|$unsigned(reg120))} : reg67))
                    begin
                      reg280 <= reg22[(3'h6):(3'h4)];
                      reg281 <= (($signed({forvar263}) ?
                          $unsigned((~|reg75)) : reg246[(3'h5):(1'h1)]) < ($signed((^reg61)) ?
                          $unsigned(reg223[(4'ha):(4'h9)]) : reg77[(1'h0):(1'h0)]));
                      reg282 <= (^~$signed(($signed(reg78) ?
                          ((8'had) ? (8'hb5) : reg28) : $unsigned(reg256))));
                    end
                  else
                    begin
                      reg280 <= (~^$unsigned(reg172));
                      reg281 <= (reg225 ?
                          ((reg275[(1'h0):(1'h0)] << (reg57 ^ reg60)) > reg135) : ($signed((reg201 ?
                              reg199 : reg33)) < ($unsigned(reg283) ?
                              reg226 : reg250)));
                      reg282 <= ((!((^reg165) ^~ reg26[(2'h2):(2'h2)])) <<< ($signed((reg193 ?
                              reg164 : reg37)) ?
                          (8'ha4) : {reg249}));
                    end
                  for (forvar283 = (1'h0); (forvar283 < (1'h0)); forvar283 = (forvar283 + (1'h1)))
                    begin
                      reg284 <= (reg221[(3'h6):(3'h5)] ^~ $signed((8'hb3)));
                      reg285 <= reg47[(2'h2):(1'h0)];
                      reg286 <= $signed(reg125[(1'h0):(1'h0)]);
                    end
                end
              for (forvar287 = (1'h0); (forvar287 < (1'h0)); forvar287 = (forvar287 + (1'h1)))
                begin
                  for (forvar288 = (1'h0); (forvar288 < (2'h2)); forvar288 = (forvar288 + (1'h1)))
                    begin
                      reg289 <= (forvar274 <= (($signed(wire0) | (~|reg187)) ?
                          $unsigned(reg8[(4'ha):(3'h6)]) : $signed((reg80 ?
                              reg79 : reg48))));
                      reg290 <= forvar283;
                      reg291 <= (~(-reg242[(4'ha):(2'h3)]));
                    end
                  if ($unsigned(($unsigned((reg121 ?
                      reg72 : reg11)) << ($unsigned(reg27) << $signed(reg146)))))
                    begin
                      reg292 <= (reg259 ?
                          ((+$signed((8'ha7))) || $signed($signed(reg13))) : $signed({(reg20 ?
                                  reg115 : reg294)}));
                      reg293 <= (+$signed(((reg272 ?
                          reg26 : (8'ha7)) || {reg143})));
                    end
                  else
                    begin
                      reg292 <= forvar287[(3'h7):(1'h0)];
                      reg293 <= $unsigned(reg138[(3'h6):(3'h4)]);
                      reg294 <= (^reg97[(1'h1):(1'h1)]);
                    end
                  if ((($unsigned((8'ha3)) ?
                      $signed($unsigned(forvar243)) : (~{reg218})) + reg42[(1'h0):(1'h0)]))
                    begin
                      reg295 <= $signed((+reg234));
                      reg296 <= $signed($signed($unsigned((reg266 ?
                          reg167 : wire240))));
                      reg297 <= $signed((~|$unsigned($signed(reg10))));
                      reg298 <= {(!($unsigned(reg181) ?
                              reg154[(4'h9):(2'h3)] : (-reg121)))};
                    end
                  else
                    begin
                      reg295 <= (|(reg19[(3'h5):(3'h4)] ?
                          {(~reg73)} : $signed(reg79[(1'h1):(1'h0)])));
                    end
                end
            end
          reg299 <= (|(~reg142));
        end
      reg300 <= (($signed($unsigned(reg61)) | reg288[(4'h8):(3'h4)]) ?
          reg193 : (reg74[(3'h7):(3'h5)] <= (reg37[(3'h7):(2'h3)] || (~^reg295))));
    end
  assign wire301 = (8'ha7);
  assign wire302 = (-((reg45[(1'h1):(1'h1)] ?
                       (reg115 == reg176) : reg29) ^~ reg37[(2'h3):(2'h2)]));
  module303 #() modinst413 (.y(wire412), .wire304(wire2), .wire307(reg146), .clk(clk), .wire308(reg216), .wire305(reg73), .wire306(reg83));
  assign wire414 = (~^reg289);
  assign wire415 = (8'hb6);
  assign wire416 = ($signed(reg194[(3'h6):(3'h4)]) ?
                       ($unsigned($signed(reg143)) <= (-(!wire5))) : ($unsigned((reg94 ?
                           reg120 : (8'hb2))) < $signed($unsigned(reg98))));
  assign wire417 = $signed($unsigned({{(8'ha4)}}));
  assign wire418 = $signed((reg169 ?
                       ($unsigned(reg224) >= (~&reg177)) : {(^~reg121)}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module303
#(parameter param411 = {((~|((8'ha1) - (8'hb0))) ? {((8'hb8) ? (8'hb5) : (8'ha1))} : ((+(8'ha9)) ? (-(8'hab)) : ((8'ha5) >>> (8'ha4))))})
(y, clk, wire308, wire307, wire306, wire305, wire304);
  output wire [(32'h454):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire308;
  input wire [(2'h2):(1'h0)] wire307;
  input wire [(4'h8):(1'h0)] wire306;
  input wire [(4'hb):(1'h0)] wire305;
  input wire signed [(4'hc):(1'h0)] wire304;
  wire signed [(3'h4):(1'h0)] wire410;
  wire [(4'hd):(1'h0)] wire313;
  wire signed [(4'h9):(1'h0)] wire312;
  wire signed [(4'hc):(1'h0)] wire311;
  wire [(4'hd):(1'h0)] wire310;
  wire signed [(3'h6):(1'h0)] wire309;
  reg signed [(5'h10):(1'h0)] reg409 = (1'h0);
  reg [(4'h8):(1'h0)] reg408 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg407 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg406 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg405 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg404 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg403 = (1'h0);
  reg [(3'h5):(1'h0)] reg401 = (1'h0);
  reg [(3'h6):(1'h0)] reg399 = (1'h0);
  reg [(4'he):(1'h0)] reg398 = (1'h0);
  reg [(3'h5):(1'h0)] reg396 = (1'h0);
  reg [(4'he):(1'h0)] reg394 = (1'h0);
  reg [(4'ha):(1'h0)] reg392 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg391 = (1'h0);
  reg [(3'h5):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg389 = (1'h0);
  reg [(3'h5):(1'h0)] reg388 = (1'h0);
  reg [(2'h3):(1'h0)] reg387 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg378 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg386 = (1'h0);
  reg [(4'hf):(1'h0)] reg385 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg384 = (1'h0);
  reg [(3'h5):(1'h0)] reg383 = (1'h0);
  reg [(4'hb):(1'h0)] reg382 = (1'h0);
  reg [(2'h3):(1'h0)] reg381 = (1'h0);
  reg [(3'h7):(1'h0)] reg380 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg379 = (1'h0);
  reg [(3'h7):(1'h0)] reg377 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg376 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg375 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg359 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg362 = (1'h0);
  reg [(2'h2):(1'h0)] reg361 = (1'h0);
  reg [(4'h8):(1'h0)] reg350 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg342 = (1'h0);
  reg [(4'ha):(1'h0)] reg334 = (1'h0);
  reg [(5'h10):(1'h0)] reg325 = (1'h0);
  reg [(4'hb):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg330 = (1'h0);
  reg [(3'h4):(1'h0)] reg372 = (1'h0);
  reg [(4'he):(1'h0)] reg371 = (1'h0);
  reg [(2'h3):(1'h0)] reg370 = (1'h0);
  reg [(5'h10):(1'h0)] reg369 = (1'h0);
  reg [(3'h7):(1'h0)] reg368 = (1'h0);
  reg [(3'h4):(1'h0)] reg367 = (1'h0);
  reg [(4'hc):(1'h0)] reg366 = (1'h0);
  reg [(2'h3):(1'h0)] reg365 = (1'h0);
  reg [(3'h5):(1'h0)] reg364 = (1'h0);
  reg [(5'h10):(1'h0)] reg363 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg360 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg358 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg357 = (1'h0);
  reg [(3'h6):(1'h0)] reg355 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg354 = (1'h0);
  reg [(4'hc):(1'h0)] reg353 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg352 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg351 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg349 = (1'h0);
  reg [(4'hb):(1'h0)] reg348 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg347 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg346 = (1'h0);
  reg [(2'h2):(1'h0)] reg344 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg343 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg341 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg340 = (1'h0);
  reg [(4'ha):(1'h0)] reg339 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg338 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg337 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg336 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg335 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg327 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg333 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg332 = (1'h0);
  reg signed [(4'he):(1'h0)] reg331 = (1'h0);
  reg [(3'h5):(1'h0)] reg329 = (1'h0);
  reg [(4'hd):(1'h0)] reg328 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg326 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg323 = (1'h0);
  reg [(2'h3):(1'h0)] reg322 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg320 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg319 = (1'h0);
  reg [(4'h8):(1'h0)] reg318 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg315 = (1'h0);
  reg [(4'h9):(1'h0)] forvar402 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar400 = (1'h0);
  reg [(4'he):(1'h0)] forvar398 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar397 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar395 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar393 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar386 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar382 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar377 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar378 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar374 = (1'h0);
  reg [(4'he):(1'h0)] forvar373 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar365 = (1'h0);
  reg [(2'h2):(1'h0)] forvar348 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar344 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar340 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar335 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar329 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar328 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar362 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar361 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar359 = (1'h0);
  reg [(3'h7):(1'h0)] forvar356 = (1'h0);
  reg [(4'h9):(1'h0)] forvar350 = (1'h0);
  reg [(3'h5):(1'h0)] forvar339 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar345 = (1'h0);
  reg [(4'h9):(1'h0)] forvar342 = (1'h0);
  reg [(5'h10):(1'h0)] forvar334 = (1'h0);
  reg [(4'hf):(1'h0)] forvar330 = (1'h0);
  reg [(4'ha):(1'h0)] forvar327 = (1'h0);
  reg [(4'hb):(1'h0)] forvar325 = (1'h0);
  reg [(4'hd):(1'h0)] forvar324 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar317 = (1'h0);
  reg [(4'hc):(1'h0)] forvar321 = (1'h0);
  reg [(4'he):(1'h0)] forvar316 = (1'h0);
  reg [(4'h8):(1'h0)] forvar314 = (1'h0);
  assign y = {wire410,
                 wire313,
                 wire312,
                 wire311,
                 wire310,
                 wire309,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg401,
                 reg399,
                 reg398,
                 reg396,
                 reg394,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg378,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg377,
                 reg376,
                 reg375,
                 reg359,
                 reg362,
                 reg361,
                 reg350,
                 reg342,
                 reg334,
                 reg325,
                 reg324,
                 reg330,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 reg360,
                 reg358,
                 reg357,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg344,
                 reg343,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg327,
                 reg333,
                 reg332,
                 reg331,
                 reg329,
                 reg328,
                 reg326,
                 reg323,
                 reg322,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg315,
                 forvar402,
                 forvar400,
                 forvar398,
                 forvar397,
                 forvar395,
                 forvar393,
                 forvar386,
                 forvar382,
                 forvar377,
                 forvar378,
                 forvar374,
                 forvar373,
                 forvar365,
                 forvar348,
                 forvar344,
                 forvar340,
                 forvar335,
                 forvar329,
                 forvar328,
                 forvar362,
                 forvar361,
                 forvar359,
                 forvar356,
                 forvar350,
                 forvar339,
                 forvar345,
                 forvar342,
                 forvar334,
                 forvar330,
                 forvar327,
                 forvar325,
                 forvar324,
                 forvar317,
                 forvar321,
                 forvar316,
                 forvar314,
                 (1'h0)};
  assign wire309 = (^(({wire306} ? wire307 : $signed((8'h9f))) ?
                       {$unsigned(wire306)} : (wire308 ?
                           wire307[(2'h2):(1'h1)] : (~wire307))));
  assign wire310 = $unsigned((wire307 - ((wire305 ^ wire308) != (^(8'hae)))));
  assign wire311 = {(~&(8'ha8))};
  assign wire312 = $signed(wire311[(3'h4):(1'h1)]);
  assign wire313 = wire309;
  always
    @(posedge clk) begin
      for (forvar314 = (1'h0); (forvar314 < (2'h3)); forvar314 = (forvar314 + (1'h1)))
        begin
          reg315 <= $unsigned($signed($signed(wire309)));
          for (forvar316 = (1'h0); (forvar316 < (2'h3)); forvar316 = (forvar316 + (1'h1)))
            begin
              if ((((8'ha6) ?
                      (+{wire307}) : ((wire311 ?
                          wire311 : wire311) - (~^wire306))) ?
                  $signed((wire305[(2'h2):(1'h1)] || {forvar316})) : (~&wire306[(2'h3):(2'h3)])))
                begin
                  if (wire309)
                    begin
                      reg317 <= {($signed({wire307}) ?
                              $signed((~|wire311)) : wire311)};
                      reg318 <= $unsigned($unsigned($unsigned((wire308 ^ wire308))));
                      reg319 <= (^~forvar316[(3'h7):(1'h1)]);
                      reg320 <= (^~(($unsigned((8'hac)) ?
                              (wire308 >>> (8'ha6)) : (wire305 ?
                                  forvar316 : forvar316)) ?
                          (!(forvar316 ?
                              wire307 : wire311)) : $unsigned((wire304 & reg315))));
                    end
                  else
                    begin
                      reg317 <= (wire304 + (^~((wire311 ?
                          (8'hae) : wire309) <= (&wire307))));
                      reg318 <= ({reg319} ?
                          ($signed(wire306[(2'h2):(1'h1)]) ?
                              forvar316 : forvar316[(4'he):(3'h4)]) : ((^~{wire305}) ?
                              ($unsigned(wire306) ^ $signed(wire305)) : forvar314[(2'h2):(2'h2)]));
                      reg319 <= {forvar316};
                    end
                  for (forvar321 = (1'h0); (forvar321 < (1'h0)); forvar321 = (forvar321 + (1'h1)))
                    begin
                      reg322 <= wire307[(1'h0):(1'h0)];
                      reg323 <= $signed((&reg317[(3'h4):(1'h1)]));
                    end
                end
              else
                begin
                  for (forvar317 = (1'h0); (forvar317 < (2'h2)); forvar317 = (forvar317 + (1'h1)))
                    begin
                      reg318 <= $signed(((8'ha6) ^ $signed($unsigned(reg320))));
                    end
                end
            end
        end
      if ($unsigned(forvar317))
        begin
          for (forvar324 = (1'h0); (forvar324 < (1'h0)); forvar324 = (forvar324 + (1'h1)))
            begin
              if (forvar321[(3'h6):(1'h1)])
                begin
                  for (forvar325 = (1'h0); (forvar325 < (2'h3)); forvar325 = (forvar325 + (1'h1)))
                    begin
                      reg326 <= forvar317[(3'h6):(3'h4)];
                    end
                  for (forvar327 = (1'h0); (forvar327 < (1'h1)); forvar327 = (forvar327 + (1'h1)))
                    begin
                      reg328 <= ({(^~$signed(forvar316))} > $unsigned(reg322));
                      reg329 <= reg323[(2'h2):(1'h1)];
                    end
                  for (forvar330 = (1'h0); (forvar330 < (2'h3)); forvar330 = (forvar330 + (1'h1)))
                    begin
                      reg331 <= $unsigned(wire312);
                      reg332 <= $signed($unsigned({(reg323 ?
                              wire305 : forvar314)}));
                    end
                  reg333 <= (8'hb1);
                end
              else
                begin
                  for (forvar325 = (1'h0); (forvar325 < (1'h0)); forvar325 = (forvar325 + (1'h1)))
                    begin
                      reg326 <= (reg331[(3'h5):(3'h4)] | ((8'hba) && reg319[(3'h5):(2'h2)]));
                      reg327 <= reg318;
                    end
                end
              if (wire310[(4'hc):(2'h3)])
                begin
                  for (forvar334 = (1'h0); (forvar334 < (1'h0)); forvar334 = (forvar334 + (1'h1)))
                    begin
                      reg335 <= ($signed(((&wire313) ?
                              (-reg331) : $unsigned(reg333))) ?
                          ($unsigned((reg333 <<< forvar324)) ?
                              (8'ha5) : ((~reg331) + (+wire312))) : forvar317);
                      reg336 <= (~(!(^forvar325)));
                      reg337 <= $unsigned(wire312[(3'h7):(1'h1)]);
                      reg338 <= reg331;
                    end
                  if ((~&(8'ha0)))
                    begin
                      reg339 <= {({(forvar316 ? reg328 : reg329)} ?
                              $unsigned($unsigned(forvar334)) : reg317[(3'h5):(2'h2)])};
                      reg340 <= (reg322[(1'h0):(1'h0)] ^~ $unsigned(forvar321[(2'h2):(1'h0)]));
                      reg341 <= $signed($unsigned((~|(~forvar316))));
                    end
                  else
                    begin
                      reg339 <= reg332;
                      reg340 <= (8'had);
                    end
                  for (forvar342 = (1'h0); (forvar342 < (1'h0)); forvar342 = (forvar342 + (1'h1)))
                    begin
                      reg343 <= (wire312 != ($signed(forvar330) ?
                          (reg320[(3'h7):(3'h6)] ?
                              (reg320 && (8'had)) : $unsigned(wire313)) : reg338[(1'h1):(1'h1)]));
                      reg344 <= $unsigned({(~(-wire306))});
                    end
                  for (forvar345 = (1'h0); (forvar345 < (1'h0)); forvar345 = (forvar345 + (1'h1)))
                    begin
                      reg346 <= (forvar327 ? (8'hb7) : (reg320 ~^ (~^wire311)));
                      reg347 <= $unsigned(reg339);
                      reg348 <= $signed($signed(reg329));
                      reg349 <= $unsigned({$signed($unsigned(reg322))});
                    end
                end
              else
                begin
                  for (forvar334 = (1'h0); (forvar334 < (2'h3)); forvar334 = (forvar334 + (1'h1)))
                    begin
                      reg335 <= $unsigned((8'hb2));
                      reg336 <= {$signed({(wire305 ^~ reg344)})};
                      reg337 <= (($signed($unsigned((8'hac))) ?
                              $unsigned($signed(forvar324)) : ((reg328 ?
                                      reg344 : forvar314) ?
                                  (~^(8'ha6)) : (-(8'ha6)))) ?
                          (8'h9c) : wire308);
                      reg338 <= (wire308[(4'hb):(4'h8)] ?
                          (^~$signed((reg333 << forvar324))) : $signed($unsigned((reg347 >= (8'ha5)))));
                    end
                  for (forvar339 = (1'h0); (forvar339 < (1'h1)); forvar339 = (forvar339 + (1'h1)))
                    begin
                      reg340 <= $signed(forvar339);
                      reg341 <= reg344[(2'h2):(1'h1)];
                    end
                end
              if (reg340[(2'h3):(1'h1)])
                begin
                  for (forvar350 = (1'h0); (forvar350 < (1'h1)); forvar350 = (forvar350 + (1'h1)))
                    begin
                      reg351 <= $signed(($unsigned((reg322 != wire309)) & forvar316[(3'h5):(3'h5)]));
                      reg352 <= $signed(reg320[(4'h8):(2'h2)]);
                    end
                  if (reg349)
                    begin
                      reg353 <= reg340[(3'h4):(3'h4)];
                      reg354 <= $signed({((reg336 ?
                              reg323 : forvar317) < (forvar334 ?
                              forvar327 : reg323))});
                      reg355 <= (~($unsigned((^~wire304)) || {(reg333 >>> wire305)}));
                    end
                  else
                    begin
                      reg353 <= reg331[(4'h9):(3'h7)];
                      reg354 <= ($unsigned((((8'ha3) ?
                              forvar339 : wire309) << $unsigned(reg338))) ?
                          $signed(($unsigned(reg351) ?
                              $signed(reg318) : {forvar334})) : $signed({(+reg340)}));
                    end
                  for (forvar356 = (1'h0); (forvar356 < (2'h3)); forvar356 = (forvar356 + (1'h1)))
                    begin
                      reg357 <= ($unsigned((^reg315)) ?
                          $unsigned(forvar317[(3'h4):(1'h1)]) : $unsigned($unsigned((reg341 ?
                              reg317 : reg318))));
                    end
                end
              else
                begin
                  for (forvar350 = (1'h0); (forvar350 < (2'h2)); forvar350 = (forvar350 + (1'h1)))
                    begin
                      reg351 <= reg341;
                      reg352 <= reg357;
                      reg353 <= (reg353[(4'h8):(2'h2)] & reg323[(2'h3):(2'h3)]);
                    end
                end
              reg358 <= {reg331[(3'h7):(3'h7)]};
            end
          for (forvar359 = (1'h0); (forvar359 < (1'h1)); forvar359 = (forvar359 + (1'h1)))
            begin
              reg360 <= {(($signed(forvar316) ?
                          forvar325[(2'h2):(2'h2)] : $signed(reg337)) ?
                      $signed((reg320 >> reg352)) : (~^(8'ha5)))};
              for (forvar361 = (1'h0); (forvar361 < (2'h2)); forvar361 = (forvar361 + (1'h1)))
                begin
                  for (forvar362 = (1'h0); (forvar362 < (1'h0)); forvar362 = (forvar362 + (1'h1)))
                    begin
                      reg363 <= reg358;
                      reg364 <= reg348;
                      reg365 <= reg357[(4'he):(4'hd)];
                    end
                  reg366 <= $signed($unsigned(reg358[(1'h1):(1'h1)]));
                  reg367 <= $unsigned({(~forvar325)});
                  if (reg332[(1'h0):(1'h0)])
                    begin
                      reg368 <= (^~{({wire310} ?
                              (forvar361 || reg347) : forvar350[(2'h2):(1'h1)])});
                      reg369 <= (($signed((~(8'hae))) ?
                          ((forvar327 ? reg349 : reg355) ?
                              ((8'hb0) + reg347) : ((8'hb1) <<< (8'ha2))) : (-(~reg357))) ^~ (({reg341} ?
                          $unsigned(reg320) : ((8'ha8) >= forvar350)) > $signed((reg346 >> reg336))));
                      reg370 <= wire313[(4'hc):(3'h7)];
                      reg371 <= $unsigned((-wire311));
                    end
                  else
                    begin
                      reg368 <= $signed($unsigned($unsigned((reg336 & forvar359))));
                      reg369 <= $unsigned($unsigned((~&((8'hb0) | reg349))));
                      reg370 <= (reg360 ?
                          $unsigned(({reg347} ?
                              (~|wire307) : (reg336 ^~ wire308))) : (~|reg323[(2'h2):(1'h1)]));
                    end
                end
              reg372 <= ((((-reg344) ~^ $unsigned(reg323)) ?
                      reg343[(1'h0):(1'h0)] : ($signed(forvar330) + wire310)) ?
                  {$unsigned(reg327[(1'h1):(1'h0)])} : $signed(reg338[(1'h1):(1'h0)]));
            end
        end
      else
        begin
          if ((8'hac))
            begin
              for (forvar324 = (1'h0); (forvar324 < (2'h3)); forvar324 = (forvar324 + (1'h1)))
                begin
                  for (forvar325 = (1'h0); (forvar325 < (1'h0)); forvar325 = (forvar325 + (1'h1)))
                    begin
                      reg326 <= wire311;
                      reg327 <= wire306;
                    end
                  for (forvar328 = (1'h0); (forvar328 < (2'h3)); forvar328 = (forvar328 + (1'h1)))
                    begin
                      reg329 <= $unsigned($signed((reg368[(3'h4):(1'h0)] * (~|reg331))));
                      reg330 <= {(reg369[(4'he):(4'hd)] && (~|$signed(reg338)))};
                    end
                end
              reg331 <= $unsigned(reg337);
            end
          else
            begin
              if ((^$signed(((8'hb5) ? reg341 : $signed(reg368)))))
                begin
                  reg324 <= (reg368 ?
                      reg323[(1'h0):(1'h0)] : $unsigned($signed({wire311})));
                  if ((^~$unsigned($signed(forvar339[(3'h4):(2'h2)]))))
                    begin
                      reg325 <= (8'hab);
                      reg326 <= reg372[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg325 <= (!(8'ha5));
                    end
                  if ((((^~(forvar321 ? wire305 : forvar317)) <= wire309) ?
                      $unsigned(((forvar327 ^~ reg371) >> $unsigned(reg329))) : (+((reg363 ?
                              reg329 : (8'hb3)) ?
                          reg346[(2'h2):(1'h1)] : {forvar359}))))
                    begin
                      reg327 <= ($unsigned($signed(((8'hb0) ?
                          forvar342 : forvar339))) <= $unsigned(reg324[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg327 <= (+((+reg364) - $signed((wire305 ?
                          reg348 : reg369))));
                      reg328 <= reg323[(2'h3):(1'h0)];
                    end
                  for (forvar329 = (1'h0); (forvar329 < (1'h0)); forvar329 = (forvar329 + (1'h1)))
                    begin
                      reg330 <= forvar356;
                    end
                end
              else
                begin
                  reg324 <= reg341;
                  if (($signed(reg358[(4'hb):(3'h6)]) <= reg338))
                    begin
                      reg325 <= $signed($unsigned($signed((|reg327))));
                      reg326 <= reg324;
                      reg327 <= $signed((^~(+$signed((8'hb8)))));
                    end
                  else
                    begin
                      reg325 <= $unsigned($signed($signed((forvar334 + wire310))));
                      reg326 <= wire306[(3'h7):(2'h2)];
                    end
                  if (wire309)
                    begin
                      reg328 <= reg370[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg328 <= reg318[(1'h1):(1'h0)];
                      reg329 <= ((^reg322) != reg332);
                      reg330 <= ((({forvar328} ?
                          forvar321 : (reg338 ?
                              reg323 : forvar362)) == (~^reg368)) == reg340[(2'h3):(2'h3)]);
                    end
                end
              if (wire312[(3'h4):(3'h4)])
                begin
                  if ($unsigned(($signed($unsigned(reg320)) ?
                      {$signed(reg322)} : (|(^~reg347)))))
                    begin
                      reg331 <= (~forvar328);
                      reg332 <= (reg328 ? reg336 : (!(~&forvar314)));
                    end
                  else
                    begin
                      reg331 <= (^(((^~wire307) | (wire310 >= reg372)) ^~ (forvar314 ?
                          $unsigned(reg358) : $unsigned(reg370))));
                      reg332 <= forvar330;
                      reg333 <= (reg317 ?
                          (reg372 ?
                              $signed((forvar314 * wire306)) : (reg319[(3'h7):(1'h0)] | (wire310 ?
                                  reg351 : reg349))) : forvar314);
                      reg334 <= (((8'hb8) ?
                              reg365[(1'h0):(1'h0)] : ((~&forvar324) ?
                                  {reg372} : (reg344 == wire304))) ?
                          {reg337[(1'h1):(1'h1)]} : ({(reg343 ?
                                      wire309 : wire305)} ?
                              forvar321[(1'h0):(1'h0)] : $unsigned((reg369 ?
                                  reg327 : (8'hab)))));
                    end
                  for (forvar335 = (1'h0); (forvar335 < (2'h2)); forvar335 = (forvar335 + (1'h1)))
                    begin
                      reg336 <= wire313;
                      reg337 <= (reg363[(3'h4):(2'h3)] ?
                          {((forvar321 ? wire311 : (8'ha4)) ?
                                  reg318 : forvar339[(2'h3):(1'h1)])} : reg357);
                      reg338 <= $signed(reg351[(3'h6):(3'h5)]);
                      reg339 <= forvar325;
                    end
                  for (forvar340 = (1'h0); (forvar340 < (2'h3)); forvar340 = (forvar340 + (1'h1)))
                    begin
                      reg341 <= $unsigned((((reg346 == reg341) ?
                          forvar314[(2'h2):(1'h1)] : forvar356[(3'h4):(1'h0)]) >= ((~(8'hae)) ?
                          $signed(forvar325) : (~^forvar330))));
                      reg342 <= forvar314;
                      reg343 <= ($unsigned(((forvar345 ? (8'ha0) : forvar342) ?
                          wire312[(1'h1):(1'h1)] : reg372)) >= (|{(8'h9d)}));
                    end
                end
              else
                begin
                  if (reg333)
                    begin
                      reg331 <= (reg322 && (~^(~|reg328[(4'hb):(4'hb)])));
                    end
                  else
                    begin
                      reg331 <= ($unsigned(forvar317[(3'h4):(1'h0)]) ?
                          (($unsigned(forvar359) ^ ((8'haf) ^~ reg335)) == $signed(reg323)) : reg340);
                      reg332 <= $unsigned((((8'ha3) << reg347[(3'h7):(1'h1)]) ?
                          forvar342[(3'h6):(3'h6)] : $unsigned((~|reg326))));
                      reg333 <= $unsigned((~forvar334));
                      reg334 <= $signed((8'hb8));
                    end
                  for (forvar335 = (1'h0); (forvar335 < (2'h2)); forvar335 = (forvar335 + (1'h1)))
                    begin
                      reg336 <= reg333;
                    end
                  if (($unsigned((wire305[(1'h1):(1'h0)] >= reg352)) ~^ {(+(wire305 ^ reg325))}))
                    begin
                      reg337 <= $unsigned($unsigned((~|$signed(reg366))));
                      reg338 <= (reg325 ?
                          forvar324[(4'hc):(1'h0)] : $unsigned($unsigned((reg348 ?
                              reg367 : (8'ha9)))));
                      reg339 <= ($signed(((reg368 ?
                          reg338 : reg331) | (forvar356 >= forvar316))) >> (reg325[(3'h7):(1'h1)] >= ((|reg358) ?
                          (~^reg339) : $unsigned((8'haa)))));
                    end
                  else
                    begin
                      reg337 <= reg341[(2'h3):(1'h0)];
                    end
                end
            end
          for (forvar344 = (1'h0); (forvar344 < (1'h0)); forvar344 = (forvar344 + (1'h1)))
            begin
              for (forvar345 = (1'h0); (forvar345 < (2'h3)); forvar345 = (forvar345 + (1'h1)))
                begin
                  reg346 <= wire309[(2'h3):(2'h3)];
                end
            end
          reg347 <= ((8'ha2) ?
              {wire312[(1'h1):(1'h1)]} : $signed(wire313[(1'h0):(1'h0)]));
          for (forvar348 = (1'h0); (forvar348 < (2'h3)); forvar348 = (forvar348 + (1'h1)))
            begin
              if ((wire311[(4'hb):(2'h2)] * ((wire306[(1'h1):(1'h1)] ?
                  $unsigned(forvar316) : reg338) & reg355[(2'h2):(1'h0)])))
                begin
                  if ($signed(reg353[(1'h0):(1'h0)]))
                    begin
                      reg349 <= {reg338};
                      reg350 <= ((wire307[(2'h2):(1'h0)] <<< (~^(^~reg355))) >> $signed($signed(reg371[(4'hc):(1'h0)])));
                      reg351 <= forvar339[(1'h1):(1'h1)];
                      reg352 <= forvar324[(3'h5):(1'h0)];
                    end
                  else
                    begin
                      reg349 <= (reg358 > reg366[(2'h3):(1'h0)]);
                      reg350 <= $unsigned(reg343);
                      reg351 <= (((~&reg351) ^~ $signed((reg317 ?
                          (8'hb8) : (8'ha3)))) == wire311);
                    end
                  if ($signed(($signed(reg349) << {$signed((8'ha9))})))
                    begin
                      reg353 <= ($signed(reg334[(4'h9):(1'h0)]) ?
                          ((^~(forvar314 * wire306)) ~^ {(|reg335)}) : $signed($signed($unsigned(reg370))));
                      reg354 <= $unsigned($unsigned(((reg357 ?
                              reg322 : reg324) ?
                          (8'hb0) : $unsigned(forvar340))));
                      reg355 <= $signed($unsigned(reg341));
                    end
                  else
                    begin
                      reg353 <= $unsigned($signed(reg358));
                      reg354 <= reg368;
                      reg355 <= forvar345;
                    end
                  for (forvar356 = (1'h0); (forvar356 < (1'h0)); forvar356 = (forvar356 + (1'h1)))
                    begin
                      reg357 <= (forvar350[(1'h1):(1'h0)] ?
                          (((~|reg334) < $signed(reg370)) ?
                              ((forvar314 != (8'ha0)) ?
                                  reg370[(2'h2):(1'h0)] : (reg353 ?
                                      reg350 : (8'h9d))) : reg322) : $signed(forvar327[(4'h8):(3'h6)]));
                      reg358 <= ((((reg325 << (8'haf)) == (reg325 ?
                              (8'h9f) : reg338)) ?
                          {(wire309 ^ (8'had))} : reg330[(5'h10):(3'h6)]) << {reg354});
                    end
                end
              else
                begin
                  if (reg354)
                    begin
                      reg349 <= forvar344[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg349 <= (~(reg338 ?
                          forvar350[(3'h5):(3'h5)] : forvar344));
                    end
                  if ($unsigned((reg342[(2'h2):(2'h2)] ?
                      $unsigned(wire309) : (&{forvar344}))))
                    begin
                      reg350 <= $signed((~&$unsigned(((8'hb1) == reg351))));
                      reg351 <= $signed(forvar348);
                    end
                  else
                    begin
                      reg350 <= $unsigned(forvar342);
                      reg351 <= ((($unsigned(reg352) ?
                              $unsigned(wire304) : (forvar335 ^~ (8'haa))) ?
                          (~{reg358}) : $unsigned($signed(reg367))) + (({forvar344} | (reg346 ?
                              forvar330 : forvar361)) ?
                          reg328 : reg324));
                    end
                end
              if ($signed((reg332[(2'h3):(1'h1)] & forvar345[(1'h0):(1'h0)])))
                begin
                  for (forvar359 = (1'h0); (forvar359 < (1'h1)); forvar359 = (forvar359 + (1'h1)))
                    begin
                      reg360 <= $signed({$signed((&forvar356))});
                      reg361 <= wire306[(3'h5):(1'h0)];
                      reg362 <= forvar344;
                      reg363 <= reg365;
                    end
                  reg364 <= reg339[(4'h9):(3'h7)];
                  for (forvar365 = (1'h0); (forvar365 < (1'h1)); forvar365 = (forvar365 + (1'h1)))
                    begin
                      reg366 <= reg327[(1'h1):(1'h1)];
                      reg367 <= ({(~^{reg327})} ~^ $unsigned($unsigned(wire305[(1'h1):(1'h1)])));
                    end
                end
              else
                begin
                  if ((reg329[(3'h5):(2'h3)] && wire306))
                    begin
                      reg359 <= $signed($signed((wire307[(1'h0):(1'h0)] <= reg351[(3'h6):(1'h0)])));
                      reg360 <= $unsigned(forvar359);
                      reg361 <= $unsigned($unsigned(reg315[(2'h2):(2'h2)]));
                      reg362 <= reg326;
                    end
                  else
                    begin
                      reg359 <= ({$signed($signed(forvar362))} != forvar317);
                      reg360 <= forvar344[(1'h1):(1'h1)];
                    end
                end
            end
        end
      if (((|$unsigned($signed(wire313))) ?
          {(^~reg368)} : forvar344[(2'h2):(1'h1)]))
        begin
          for (forvar373 = (1'h0); (forvar373 < (2'h3)); forvar373 = (forvar373 + (1'h1)))
            begin
              for (forvar374 = (1'h0); (forvar374 < (1'h0)); forvar374 = (forvar374 + (1'h1)))
                begin
                  if (forvar316[(4'hb):(4'h9)])
                    begin
                      reg375 <= reg341[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg375 <= (~&(~&($unsigned(reg327) ~^ $signed(reg371))));
                      reg376 <= $signed($signed((~$signed(forvar321))));
                      reg377 <= {(8'h9d)};
                    end
                  for (forvar378 = (1'h0); (forvar378 < (2'h2)); forvar378 = (forvar378 + (1'h1)))
                    begin
                      reg379 <= (((^reg375) < forvar316[(4'ha):(3'h4)]) ?
                          (-(-$signed(reg359))) : $unsigned(reg367[(2'h3):(2'h2)]));
                      reg380 <= forvar316;
                      reg381 <= ((reg360[(3'h7):(2'h2)] ~^ reg370[(2'h3):(2'h3)]) ?
                          forvar359 : (~reg353));
                      reg382 <= forvar328;
                    end
                  if (reg346[(1'h0):(1'h0)])
                    begin
                      reg383 <= forvar344[(3'h4):(2'h3)];
                      reg384 <= (reg347 ?
                          ((-(reg320 << reg319)) ?
                              wire305 : $signed({(8'h9e)})) : (($unsigned(reg375) <= forvar330[(1'h1):(1'h0)]) ?
                              reg318[(2'h3):(1'h0)] : ({reg380} & reg368)));
                      reg385 <= (+$signed(forvar321));
                      reg386 <= (forvar378 != (|((-(8'hb4)) ?
                          (^~(8'ha5)) : $signed(reg333))));
                    end
                  else
                    begin
                      reg383 <= forvar373[(4'hc):(3'h6)];
                      reg384 <= $signed((+$signed((reg381 <<< (8'ha1)))));
                    end
                end
            end
        end
      else
        begin
          for (forvar373 = (1'h0); (forvar373 < (2'h3)); forvar373 = (forvar373 + (1'h1)))
            begin
              for (forvar374 = (1'h0); (forvar374 < (2'h3)); forvar374 = (forvar374 + (1'h1)))
                begin
                  if ($signed($unsigned((reg383[(2'h2):(1'h1)] ?
                      (forvar362 ? reg355 : forvar344) : (~|(8'h9d))))))
                    begin
                      reg375 <= (wire306[(3'h6):(2'h2)] || (((forvar330 ?
                              forvar329 : forvar365) ?
                          {reg315} : (8'ha6)) == $signed($signed(reg357))));
                      reg376 <= reg375;
                    end
                  else
                    begin
                      reg375 <= $signed((wire307[(1'h0):(1'h0)] ^~ reg386[(2'h2):(1'h1)]));
                      reg376 <= {{reg363}};
                    end
                  for (forvar377 = (1'h0); (forvar377 < (2'h2)); forvar377 = (forvar377 + (1'h1)))
                    begin
                      reg378 <= reg346[(1'h0):(1'h0)];
                      reg379 <= {forvar348[(2'h2):(1'h1)]};
                      reg380 <= (~^(&reg359));
                      reg381 <= {$unsigned(($signed(forvar378) ^ forvar339[(2'h2):(1'h0)]))};
                    end
                end
              for (forvar382 = (1'h0); (forvar382 < (2'h2)); forvar382 = (forvar382 + (1'h1)))
                begin
                  if ($signed($signed((reg319 ?
                      (reg376 ? reg335 : (8'h9f)) : forvar339))))
                    begin
                      reg383 <= (reg358 == ($signed((~|wire307)) ?
                          $unsigned((~^(8'had))) : ((forvar356 << reg365) || (forvar345 >>> reg340))));
                      reg384 <= (~{{reg381[(1'h1):(1'h0)]}});
                      reg385 <= wire312;
                    end
                  else
                    begin
                      reg383 <= ($signed(forvar362[(4'he):(1'h1)]) ?
                          ($signed((-forvar321)) ?
                              (|$signed(reg353)) : reg349) : (^forvar330));
                    end
                  for (forvar386 = (1'h0); (forvar386 < (1'h0)); forvar386 = (forvar386 + (1'h1)))
                    begin
                      reg387 <= $unsigned(reg366[(1'h0):(1'h0)]);
                      reg388 <= reg331[(4'hc):(1'h0)];
                    end
                  if (((&forvar382[(3'h4):(1'h0)]) | $signed(forvar359)))
                    begin
                      reg389 <= forvar339;
                      reg390 <= $signed({($signed(reg384) ?
                              (reg367 ?
                                  wire307 : (8'had)) : (reg365 >>> forvar342))});
                      reg391 <= $unsigned(forvar359);
                      reg392 <= $unsigned((((reg320 ? reg331 : reg331) ?
                              reg377 : $signed(wire305)) ?
                          reg322[(2'h3):(2'h3)] : ($unsigned(reg340) <= (reg364 < reg317))));
                    end
                  else
                    begin
                      reg389 <= {(~&{reg360[(1'h0):(1'h0)]})};
                      reg390 <= (^~(^((reg334 != reg375) ?
                          (forvar342 ? reg343 : reg387) : (-forvar324))));
                      reg391 <= (~^($unsigned((reg364 ?
                          forvar359 : forvar382)) || $unsigned((reg392 != forvar386))));
                    end
                end
              for (forvar393 = (1'h0); (forvar393 < (1'h0)); forvar393 = (forvar393 + (1'h1)))
                begin
                  reg394 <= ((~&wire306[(3'h6):(1'h1)]) != {$signed((|reg385))});
                  for (forvar395 = (1'h0); (forvar395 < (1'h0)); forvar395 = (forvar395 + (1'h1)))
                    begin
                      reg396 <= $unsigned(($signed(forvar344[(3'h4):(2'h2)]) ?
                          ($signed(reg318) ?
                              reg339[(1'h0):(1'h0)] : $signed((8'hb8))) : reg389[(4'he):(1'h1)]));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar397 = (1'h0); (forvar397 < (2'h3)); forvar397 = (forvar397 + (1'h1)))
        begin
          if (({reg342} ?
              $unsigned((reg370[(2'h3):(2'h3)] << $unsigned(reg318))) : ($unsigned($signed((8'ha4))) && (8'haa))))
            begin
              reg398 <= (~&(~&$unsigned($signed(reg339))));
            end
          else
            begin
              for (forvar398 = (1'h0); (forvar398 < (1'h0)); forvar398 = (forvar398 + (1'h1)))
                begin
                  reg399 <= reg364[(3'h4):(3'h4)];
                  for (forvar400 = (1'h0); (forvar400 < (1'h1)); forvar400 = (forvar400 + (1'h1)))
                    begin
                      reg401 <= (reg379 == (-$unsigned($unsigned(reg317))));
                    end
                end
              for (forvar402 = (1'h0); (forvar402 < (2'h3)); forvar402 = (forvar402 + (1'h1)))
                begin
                  if ($signed((-reg350)))
                    begin
                      reg403 <= (reg364[(3'h4):(2'h2)] != reg358[(3'h4):(3'h4)]);
                      reg404 <= {($signed($unsigned(reg348)) ?
                              $unsigned(reg323[(1'h1):(1'h1)]) : $signed($unsigned(reg362)))};
                      reg405 <= (^~(+((-reg361) ^~ (reg403 >= reg329))));
                      reg406 <= $unsigned(({(~wire308)} ?
                          $signed((reg336 ?
                              (8'had) : (8'hb8))) : $signed(reg334)));
                    end
                  else
                    begin
                      reg403 <= $unsigned($unsigned(((reg343 ?
                              reg351 : reg348) ?
                          reg329[(1'h1):(1'h1)] : $signed(reg346))));
                    end
                  if (reg366[(3'h4):(3'h4)])
                    begin
                      reg407 <= $signed(reg369[(3'h7):(1'h1)]);
                      reg408 <= $signed($signed(forvar397));
                      reg409 <= $signed(($signed($unsigned(reg354)) ?
                          (~reg385[(4'he):(3'h5)]) : {((8'haf) ^ reg404)}));
                    end
                  else
                    begin
                      reg407 <= ((^~$unsigned(((8'ha4) ~^ reg337))) ?
                          $signed((~&$unsigned(reg399))) : (reg349 <= wire309));
                      reg408 <= reg388[(3'h5):(3'h5)];
                      reg409 <= $unsigned(reg404[(2'h3):(2'h3)]);
                    end
                end
            end
        end
    end
  assign wire410 = reg382;
endmodule