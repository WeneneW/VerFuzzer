(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'hab3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire0;
  input wire [(4'he):(1'h0)] wire1;
  input wire [(5'h10):(1'h0)] wire2;
  input wire signed [(2'h2):(1'h0)] wire3;
  wire signed [(5'h10):(1'h0)] wire1065;
  wire signed [(3'h5):(1'h0)] wire1064;
  wire [(4'h8):(1'h0)] wire836;
  wire [(4'h8):(1'h0)] wire4;
  wire [(5'h10):(1'h0)] wire5;
  wire [(3'h5):(1'h0)] wire834;
  reg signed [(4'h8):(1'h0)] reg1063 = (1'h0);
  reg [(4'hb):(1'h0)] reg1062 = (1'h0);
  reg [(3'h5):(1'h0)] reg1057 = (1'h0);
  reg [(4'hc):(1'h0)] reg1061 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1060 = (1'h0);
  reg [(4'ha):(1'h0)] reg1059 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1058 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1056 = (1'h0);
  reg [(4'hc):(1'h0)] reg1055 = (1'h0);
  reg [(4'hc):(1'h0)] reg1054 = (1'h0);
  reg [(4'h8):(1'h0)] reg1053 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1052 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1051 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1050 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1049 = (1'h0);
  reg [(4'ha):(1'h0)] reg1048 = (1'h0);
  reg [(4'hd):(1'h0)] reg1046 = (1'h0);
  reg [(4'hc):(1'h0)] reg1044 = (1'h0);
  reg [(3'h5):(1'h0)] reg1037 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1047 = (1'h0);
  reg [(4'he):(1'h0)] reg1045 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1043 = (1'h0);
  reg [(2'h2):(1'h0)] reg1042 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1041 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1040 = (1'h0);
  reg [(4'hb):(1'h0)] reg1039 = (1'h0);
  reg [(4'hd):(1'h0)] reg1038 = (1'h0);
  reg [(4'h8):(1'h0)] reg1036 = (1'h0);
  reg [(4'he):(1'h0)] reg1035 = (1'h0);
  reg [(4'h9):(1'h0)] reg1034 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1031 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1030 = (1'h0);
  reg [(2'h2):(1'h0)] reg1029 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1028 = (1'h0);
  reg [(2'h3):(1'h0)] reg1027 = (1'h0);
  reg [(3'h5):(1'h0)] reg1026 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1025 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1024 = (1'h0);
  reg [(4'ha):(1'h0)] reg1023 = (1'h0);
  reg [(4'hf):(1'h0)] reg1022 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1021 = (1'h0);
  reg [(2'h3):(1'h0)] reg1020 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1019 = (1'h0);
  reg [(3'h7):(1'h0)] reg1014 = (1'h0);
  reg [(4'hc):(1'h0)] reg1002 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg986 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg981 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1017 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1016 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1015 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1013 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1010 = (1'h0);
  reg [(4'h9):(1'h0)] reg1007 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1011 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1009 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1008 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1006 = (1'h0);
  reg [(4'hb):(1'h0)] reg1005 = (1'h0);
  reg [(4'hc):(1'h0)] reg1004 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1003 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg999 = (1'h0);
  reg [(4'h9):(1'h0)] reg995 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg992 = (1'h0);
  reg [(4'hf):(1'h0)] reg1001 = (1'h0);
  reg [(4'he):(1'h0)] reg1000 = (1'h0);
  reg [(4'h8):(1'h0)] reg998 = (1'h0);
  reg [(4'hd):(1'h0)] reg997 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg996 = (1'h0);
  reg signed [(4'he):(1'h0)] reg994 = (1'h0);
  reg signed [(4'he):(1'h0)] reg993 = (1'h0);
  reg [(4'hd):(1'h0)] reg991 = (1'h0);
  reg [(4'hb):(1'h0)] reg990 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg989 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg988 = (1'h0);
  reg [(4'hd):(1'h0)] reg987 = (1'h0);
  reg [(2'h2):(1'h0)] reg985 = (1'h0);
  reg [(4'he):(1'h0)] reg984 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg983 = (1'h0);
  reg [(4'h9):(1'h0)] reg982 = (1'h0);
  reg signed [(4'he):(1'h0)] reg980 = (1'h0);
  reg [(4'hb):(1'h0)] reg979 = (1'h0);
  reg [(2'h2):(1'h0)] reg978 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg977 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg975 = (1'h0);
  reg [(4'h9):(1'h0)] reg976 = (1'h0);
  reg [(4'h9):(1'h0)] reg974 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg973 = (1'h0);
  reg [(4'he):(1'h0)] reg972 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg971 = (1'h0);
  reg [(3'h7):(1'h0)] reg970 = (1'h0);
  reg [(4'h8):(1'h0)] reg968 = (1'h0);
  reg [(4'he):(1'h0)] reg963 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg958 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg957 = (1'h0);
  reg [(4'h9):(1'h0)] reg954 = (1'h0);
  reg [(3'h4):(1'h0)] reg943 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg942 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg935 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg940 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg937 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg934 = (1'h0);
  reg [(4'hc):(1'h0)] reg918 = (1'h0);
  reg [(4'h8):(1'h0)] reg917 = (1'h0);
  reg [(5'h10):(1'h0)] reg915 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg907 = (1'h0);
  reg [(5'h10):(1'h0)] reg967 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg966 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg965 = (1'h0);
  reg [(3'h4):(1'h0)] reg964 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg962 = (1'h0);
  reg [(4'hd):(1'h0)] reg961 = (1'h0);
  reg [(4'he):(1'h0)] reg960 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg959 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg956 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg955 = (1'h0);
  reg [(4'hd):(1'h0)] reg953 = (1'h0);
  reg [(4'hb):(1'h0)] reg952 = (1'h0);
  reg [(3'h6):(1'h0)] reg951 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg950 = (1'h0);
  reg [(3'h4):(1'h0)] reg949 = (1'h0);
  reg [(4'h9):(1'h0)] reg948 = (1'h0);
  reg [(3'h5):(1'h0)] reg947 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg946 = (1'h0);
  reg [(4'ha):(1'h0)] reg945 = (1'h0);
  reg [(5'h10):(1'h0)] reg944 = (1'h0);
  reg signed [(4'he):(1'h0)] reg941 = (1'h0);
  reg [(4'he):(1'h0)] reg939 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg938 = (1'h0);
  reg [(4'he):(1'h0)] reg936 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg925 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg933 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg932 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg931 = (1'h0);
  reg [(3'h4):(1'h0)] reg930 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg929 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg928 = (1'h0);
  reg [(3'h7):(1'h0)] reg927 = (1'h0);
  reg [(5'h10):(1'h0)] reg926 = (1'h0);
  reg [(2'h3):(1'h0)] reg924 = (1'h0);
  reg [(4'hf):(1'h0)] reg923 = (1'h0);
  reg [(4'hb):(1'h0)] reg922 = (1'h0);
  reg [(3'h5):(1'h0)] reg921 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg920 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg919 = (1'h0);
  reg [(3'h6):(1'h0)] reg916 = (1'h0);
  reg [(5'h10):(1'h0)] reg914 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg913 = (1'h0);
  reg [(3'h4):(1'h0)] reg912 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg911 = (1'h0);
  reg [(3'h5):(1'h0)] reg910 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg909 = (1'h0);
  reg [(4'he):(1'h0)] reg908 = (1'h0);
  reg [(2'h3):(1'h0)] reg906 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg905 = (1'h0);
  reg [(3'h4):(1'h0)] reg904 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg903 = (1'h0);
  reg [(3'h5):(1'h0)] reg902 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg900 = (1'h0);
  reg [(5'h10):(1'h0)] reg899 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg898 = (1'h0);
  reg [(3'h4):(1'h0)] reg897 = (1'h0);
  reg [(4'hb):(1'h0)] reg896 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg895 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg894 = (1'h0);
  reg [(3'h7):(1'h0)] reg893 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg891 = (1'h0);
  reg [(3'h6):(1'h0)] reg890 = (1'h0);
  reg [(3'h5):(1'h0)] reg889 = (1'h0);
  reg [(4'ha):(1'h0)] reg886 = (1'h0);
  reg [(4'hc):(1'h0)] reg885 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg884 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg883 = (1'h0);
  reg [(2'h2):(1'h0)] reg882 = (1'h0);
  reg [(4'hf):(1'h0)] reg881 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg879 = (1'h0);
  reg [(2'h2):(1'h0)] reg878 = (1'h0);
  reg [(4'hc):(1'h0)] reg877 = (1'h0);
  reg [(3'h6):(1'h0)] reg875 = (1'h0);
  reg [(3'h4):(1'h0)] reg874 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg873 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg872 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg870 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg868 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg867 = (1'h0);
  reg [(4'hb):(1'h0)] reg866 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg865 = (1'h0);
  reg [(3'h6):(1'h0)] reg838 = (1'h0);
  reg [(3'h6):(1'h0)] reg862 = (1'h0);
  reg [(4'hb):(1'h0)] reg861 = (1'h0);
  reg [(4'h9):(1'h0)] reg860 = (1'h0);
  reg [(3'h4):(1'h0)] reg859 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg858 = (1'h0);
  reg signed [(4'he):(1'h0)] reg857 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg856 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg855 = (1'h0);
  reg [(3'h6):(1'h0)] reg854 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg853 = (1'h0);
  reg [(4'hc):(1'h0)] reg852 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg850 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg849 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg848 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg847 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg846 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg845 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg844 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg843 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg842 = (1'h0);
  reg [(4'hb):(1'h0)] reg841 = (1'h0);
  reg signed [(4'he):(1'h0)] reg840 = (1'h0);
  reg signed [(4'he):(1'h0)] reg839 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1052 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1057 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1043 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1038 = (1'h0);
  reg [(4'he):(1'h0)] forvar1046 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1044 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1037 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1033 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1032 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1028 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1024 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1022 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1018 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1013 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1011 = (1'h0);
  reg [(4'he):(1'h0)] forvar998 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar993 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar990 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar984 = (1'h0);
  reg [(4'ha):(1'h0)] forvar979 = (1'h0);
  reg [(4'ha):(1'h0)] forvar978 = (1'h0);
  reg [(4'hc):(1'h0)] forvar977 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1014 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1005 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1010 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1007 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1002 = (1'h0);
  reg [(4'hd):(1'h0)] forvar994 = (1'h0);
  reg [(4'he):(1'h0)] forvar999 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar995 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar992 = (1'h0);
  reg [(4'h9):(1'h0)] forvar986 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar981 = (1'h0);
  reg [(4'hc):(1'h0)] forvar971 = (1'h0);
  reg [(4'h8):(1'h0)] forvar975 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar969 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar967 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar966 = (1'h0);
  reg [(4'he):(1'h0)] forvar965 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar959 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar956 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar955 = (1'h0);
  reg [(3'h7):(1'h0)] forvar948 = (1'h0);
  reg [(3'h7):(1'h0)] forvar947 = (1'h0);
  reg [(4'hd):(1'h0)] forvar946 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar944 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar927 = (1'h0);
  reg [(2'h2):(1'h0)] forvar921 = (1'h0);
  reg [(5'h10):(1'h0)] forvar938 = (1'h0);
  reg [(4'hf):(1'h0)] forvar933 = (1'h0);
  reg [(3'h7):(1'h0)] forvar920 = (1'h0);
  reg [(4'hf):(1'h0)] forvar928 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar924 = (1'h0);
  reg [(2'h3):(1'h0)] forvar919 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar916 = (1'h0);
  reg [(3'h5):(1'h0)] forvar912 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar963 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar958 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar957 = (1'h0);
  reg [(2'h2):(1'h0)] forvar954 = (1'h0);
  reg [(3'h5):(1'h0)] forvar943 = (1'h0);
  reg [(3'h7):(1'h0)] forvar942 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar940 = (1'h0);
  reg [(2'h2):(1'h0)] forvar937 = (1'h0);
  reg [(3'h5):(1'h0)] forvar935 = (1'h0);
  reg [(4'h8):(1'h0)] forvar934 = (1'h0);
  reg [(4'hc):(1'h0)] forvar922 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar925 = (1'h0);
  reg [(3'h7):(1'h0)] forvar918 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar917 = (1'h0);
  reg [(4'hb):(1'h0)] forvar908 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar915 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar907 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar901 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar900 = (1'h0);
  reg [(3'h5):(1'h0)] forvar892 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar888 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar887 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar883 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar880 = (1'h0);
  reg [(3'h7):(1'h0)] forvar876 = (1'h0);
  reg [(4'he):(1'h0)] forvar871 = (1'h0);
  reg [(4'he):(1'h0)] forvar869 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar864 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar863 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar847 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar844 = (1'h0);
  reg [(5'h10):(1'h0)] forvar842 = (1'h0);
  reg [(3'h7):(1'h0)] forvar858 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar851 = (1'h0);
  reg [(2'h2):(1'h0)] forvar838 = (1'h0);
  reg [(4'he):(1'h0)] forvar837 = (1'h0);
  assign y = {wire1065,
                 wire1064,
                 wire836,
                 wire4,
                 wire5,
                 wire834,
                 reg1063,
                 reg1062,
                 reg1057,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 reg1056,
                 reg1055,
                 reg1054,
                 reg1053,
                 reg1052,
                 reg1051,
                 reg1050,
                 reg1049,
                 reg1048,
                 reg1046,
                 reg1044,
                 reg1037,
                 reg1047,
                 reg1045,
                 reg1043,
                 reg1042,
                 reg1041,
                 reg1040,
                 reg1039,
                 reg1038,
                 reg1036,
                 reg1035,
                 reg1034,
                 reg1031,
                 reg1030,
                 reg1029,
                 reg1028,
                 reg1027,
                 reg1026,
                 reg1025,
                 reg1024,
                 reg1023,
                 reg1022,
                 reg1021,
                 reg1020,
                 reg1019,
                 reg1014,
                 reg1002,
                 reg986,
                 reg981,
                 reg1017,
                 reg1016,
                 reg1015,
                 reg1013,
                 reg1012,
                 reg1010,
                 reg1007,
                 reg1011,
                 reg1009,
                 reg1008,
                 reg1006,
                 reg1005,
                 reg1004,
                 reg1003,
                 reg999,
                 reg995,
                 reg992,
                 reg1001,
                 reg1000,
                 reg998,
                 reg997,
                 reg996,
                 reg994,
                 reg993,
                 reg991,
                 reg990,
                 reg989,
                 reg988,
                 reg987,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 reg980,
                 reg979,
                 reg978,
                 reg977,
                 reg975,
                 reg976,
                 reg974,
                 reg973,
                 reg972,
                 reg971,
                 reg970,
                 reg968,
                 reg963,
                 reg958,
                 reg957,
                 reg954,
                 reg943,
                 reg942,
                 reg935,
                 reg940,
                 reg937,
                 reg934,
                 reg918,
                 reg917,
                 reg915,
                 reg907,
                 reg967,
                 reg966,
                 reg965,
                 reg964,
                 reg962,
                 reg961,
                 reg960,
                 reg959,
                 reg956,
                 reg955,
                 reg953,
                 reg952,
                 reg951,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 reg946,
                 reg945,
                 reg944,
                 reg941,
                 reg939,
                 reg938,
                 reg936,
                 reg925,
                 reg933,
                 reg932,
                 reg931,
                 reg930,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 reg924,
                 reg923,
                 reg922,
                 reg921,
                 reg920,
                 reg919,
                 reg916,
                 reg914,
                 reg913,
                 reg912,
                 reg911,
                 reg910,
                 reg909,
                 reg908,
                 reg906,
                 reg905,
                 reg904,
                 reg903,
                 reg902,
                 reg900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg891,
                 reg890,
                 reg889,
                 reg886,
                 reg885,
                 reg884,
                 reg883,
                 reg882,
                 reg881,
                 reg879,
                 reg878,
                 reg877,
                 reg875,
                 reg874,
                 reg873,
                 reg872,
                 reg870,
                 reg868,
                 reg867,
                 reg866,
                 reg865,
                 reg838,
                 reg862,
                 reg861,
                 reg860,
                 reg859,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 reg852,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 reg846,
                 reg845,
                 reg844,
                 reg843,
                 reg842,
                 reg841,
                 reg840,
                 reg839,
                 forvar1052,
                 forvar1057,
                 forvar1043,
                 forvar1038,
                 forvar1046,
                 forvar1044,
                 forvar1037,
                 forvar1033,
                 forvar1032,
                 forvar1028,
                 forvar1024,
                 forvar1022,
                 forvar1018,
                 forvar1013,
                 forvar1011,
                 forvar998,
                 forvar993,
                 forvar990,
                 forvar984,
                 forvar979,
                 forvar978,
                 forvar977,
                 forvar1014,
                 forvar1005,
                 forvar1010,
                 forvar1007,
                 forvar1002,
                 forvar994,
                 forvar999,
                 forvar995,
                 forvar992,
                 forvar986,
                 forvar981,
                 forvar971,
                 forvar975,
                 forvar969,
                 forvar967,
                 forvar966,
                 forvar965,
                 forvar959,
                 forvar956,
                 forvar955,
                 forvar948,
                 forvar947,
                 forvar946,
                 forvar944,
                 forvar927,
                 forvar921,
                 forvar938,
                 forvar933,
                 forvar920,
                 forvar928,
                 forvar924,
                 forvar919,
                 forvar916,
                 forvar912,
                 forvar963,
                 forvar958,
                 forvar957,
                 forvar954,
                 forvar943,
                 forvar942,
                 forvar940,
                 forvar937,
                 forvar935,
                 forvar934,
                 forvar922,
                 forvar925,
                 forvar918,
                 forvar917,
                 forvar908,
                 forvar915,
                 forvar907,
                 forvar901,
                 forvar900,
                 forvar892,
                 forvar888,
                 forvar887,
                 forvar883,
                 forvar880,
                 forvar876,
                 forvar871,
                 forvar869,
                 forvar864,
                 forvar863,
                 forvar847,
                 forvar844,
                 forvar842,
                 forvar858,
                 forvar851,
                 forvar838,
                 forvar837,
                 (1'h0)};
  assign wire4 = wire0;
  assign wire5 = (($unsigned(wire2) << $signed((wire2 & wire4))) >= $unsigned(($signed((8'haa)) ?
                     wire3[(2'h2):(2'h2)] : $unsigned((8'hac)))));
  module6 #() modinst835 (wire834, clk, wire2, wire5, wire4, wire1, wire0);
  assign wire836 = wire5;
  always
    @(posedge clk) begin
      for (forvar837 = (1'h0); (forvar837 < (1'h1)); forvar837 = (forvar837 + (1'h1)))
        begin
          if ((8'hb7))
            begin
              for (forvar838 = (1'h0); (forvar838 < (2'h2)); forvar838 = (forvar838 + (1'h1)))
                begin
                  if (wire3[(2'h2):(2'h2)])
                    begin
                      reg839 <= wire834;
                      reg840 <= $signed((wire4[(3'h4):(1'h1)] ^~ (wire1 ?
                          $signed(reg839) : $signed(reg839))));
                      reg841 <= ($unsigned(wire5) ?
                          reg840[(3'h6):(2'h2)] : wire836);
                      reg842 <= wire2;
                    end
                  else
                    begin
                      reg839 <= $unsigned(wire834[(3'h4):(1'h1)]);
                    end
                  if ($unsigned($signed(wire1)))
                    begin
                      reg843 <= (&$signed(forvar837[(3'h6):(2'h3)]));
                      reg844 <= (~^wire0);
                      reg845 <= (!$unsigned((|(wire1 >> reg841))));
                      reg846 <= ((({wire1} <<< reg841[(3'h7):(1'h0)]) < $unsigned(wire836[(3'h7):(3'h5)])) ?
                          $unsigned(((forvar838 ?
                              wire1 : reg845) ^~ $signed(forvar838))) : (8'ha1));
                    end
                  else
                    begin
                      reg843 <= ((~^$unsigned($signed(reg839))) && (~&((reg845 ?
                              reg841 : forvar838) ?
                          $signed(wire2) : (&(8'hb5)))));
                    end
                  if (((~^(|((8'hb6) ? wire836 : forvar837))) ?
                      (wire2 >= $signed(forvar837[(4'h8):(1'h0)])) : wire834))
                    begin
                      reg847 <= $unsigned((~|($unsigned(reg839) ^ {(8'hb0)})));
                      reg848 <= $signed({{(8'haf)}});
                    end
                  else
                    begin
                      reg847 <= ((^reg842) || reg844);
                      reg848 <= ($unsigned(reg841[(1'h0):(1'h0)]) + (~|$signed((forvar838 ?
                          wire5 : wire5))));
                      reg849 <= reg841;
                      reg850 <= $unsigned($unsigned(($unsigned(reg849) >= (wire3 ?
                          wire1 : wire3))));
                    end
                  for (forvar851 = (1'h0); (forvar851 < (1'h1)); forvar851 = (forvar851 + (1'h1)))
                    begin
                      reg852 <= reg841[(2'h3):(2'h3)];
                      reg853 <= $unsigned(forvar851);
                    end
                end
              if ($unsigned(wire3))
                begin
                  if (($signed((&reg849)) ^ ($unsigned(reg848[(3'h6):(3'h4)]) >> $signed($signed(forvar851)))))
                    begin
                      reg854 <= $unsigned(((forvar837[(1'h0):(1'h0)] & reg840[(3'h4):(2'h2)]) ~^ ((!reg843) ^ $unsigned(wire834))));
                      reg855 <= reg852[(1'h0):(1'h0)];
                      reg856 <= ((reg839[(4'h9):(2'h2)] ^~ $unsigned(reg841)) ?
                          forvar837[(3'h7):(3'h7)] : reg855);
                      reg857 <= ($unsigned($unsigned((8'hb5))) ?
                          ((8'ha0) << reg856) : reg848[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg854 <= {((reg850[(4'ha):(2'h2)] ?
                              reg843 : $signed(reg849)) < $unsigned({reg843}))};
                      reg855 <= $unsigned($unsigned(forvar837[(4'hc):(4'hc)]));
                    end
                  if ($unsigned(forvar851[(2'h2):(2'h2)]))
                    begin
                      reg858 <= ((reg840[(4'he):(1'h1)] ?
                          $signed((reg841 != wire836)) : reg839) + ((&reg856) && {{wire3}}));
                    end
                  else
                    begin
                      reg858 <= reg847[(4'hb):(4'hb)];
                      reg859 <= {$signed(($unsigned(wire3) ?
                              $signed((8'ha7)) : $unsigned(reg845)))};
                      reg860 <= ((&(wire3[(1'h0):(1'h0)] ?
                          (reg848 ?
                              reg844 : forvar838) : wire5[(1'h1):(1'h1)])) != (wire3[(2'h2):(1'h0)] >> ($signed(reg849) | (8'hb0))));
                    end
                  if ($unsigned((reg850 ?
                      $unsigned({reg842}) : $signed((!wire5)))))
                    begin
                      reg861 <= $unsigned((!$unsigned($unsigned(reg854))));
                      reg862 <= $signed($unsigned((!$signed(reg848))));
                    end
                  else
                    begin
                      reg861 <= $signed(forvar837[(4'h9):(3'h6)]);
                    end
                end
              else
                begin
                  if ($unsigned($signed($signed((reg844 || reg862)))))
                    begin
                      reg854 <= $unsigned((^~wire834[(2'h2):(1'h1)]));
                      reg855 <= ((wire0 || (~&reg840)) ?
                          $signed(reg840[(2'h3):(1'h1)]) : {($unsigned((8'ha6)) ?
                                  (^(8'hb5)) : reg845[(1'h1):(1'h0)])});
                    end
                  else
                    begin
                      reg854 <= (!($signed((~&reg857)) ?
                          reg850 : (reg861[(3'h4):(1'h0)] * (wire1 << wire1))));
                      reg855 <= reg849[(3'h7):(3'h4)];
                      reg856 <= (+(reg839[(4'hc):(4'hc)] <= $signed((reg861 && reg844))));
                      reg857 <= (|(-($signed(reg846) ?
                          reg845 : $unsigned(wire836))));
                    end
                  for (forvar858 = (1'h0); (forvar858 < (2'h2)); forvar858 = (forvar858 + (1'h1)))
                    begin
                      reg859 <= forvar858[(3'h4):(2'h2)];
                      reg860 <= reg839;
                      reg861 <= $signed($unsigned(({reg850} ~^ wire1[(4'ha):(4'ha)])));
                    end
                end
            end
          else
            begin
              if (wire1)
                begin
                  for (forvar838 = (1'h0); (forvar838 < (2'h2)); forvar838 = (forvar838 + (1'h1)))
                    begin
                      reg839 <= {$unsigned(reg861)};
                      reg840 <= (($signed(reg858) ? forvar851 : reg861) ?
                          $signed($unsigned(reg846[(2'h2):(2'h2)])) : $signed(((reg855 ?
                                  reg860 : wire0) ?
                              reg839 : $unsigned(reg843))));
                      reg841 <= reg848;
                      reg842 <= forvar851;
                    end
                end
              else
                begin
                  if ($unsigned({(~^{(8'hba)})}))
                    begin
                      reg838 <= wire834;
                    end
                  else
                    begin
                      reg838 <= $signed((reg840 != ($signed(reg839) ?
                          reg853[(3'h5):(1'h0)] : reg843[(2'h3):(1'h0)])));
                      reg839 <= reg839;
                      reg840 <= (~^$unsigned({forvar858}));
                      reg841 <= reg841;
                    end
                  for (forvar842 = (1'h0); (forvar842 < (2'h2)); forvar842 = (forvar842 + (1'h1)))
                    begin
                      reg843 <= reg839[(4'hb):(4'hb)];
                    end
                  for (forvar844 = (1'h0); (forvar844 < (2'h3)); forvar844 = (forvar844 + (1'h1)))
                    begin
                      reg845 <= (reg849[(2'h3):(1'h0)] ?
                          reg854 : reg859[(2'h2):(1'h1)]);
                      reg846 <= (reg840 ?
                          (reg842[(2'h3):(2'h3)] | (((8'haf) ~^ wire0) != (forvar837 ?
                              reg854 : forvar838))) : (|$signed(wire836)));
                    end
                  for (forvar847 = (1'h0); (forvar847 < (1'h1)); forvar847 = (forvar847 + (1'h1)))
                    begin
                      reg848 <= (((8'h9f) || ($unsigned(reg853) ^ reg854[(2'h2):(1'h0)])) ?
                          {(wire1 - (forvar851 ?
                                  wire0 : reg843))} : (^~$unsigned((+forvar858))));
                      reg849 <= forvar838[(1'h0):(1'h0)];
                    end
                end
            end
          for (forvar863 = (1'h0); (forvar863 < (2'h2)); forvar863 = (forvar863 + (1'h1)))
            begin
              for (forvar864 = (1'h0); (forvar864 < (2'h2)); forvar864 = (forvar864 + (1'h1)))
                begin
                  if (reg842)
                    begin
                      reg865 <= ((^~forvar864) ? reg846 : reg849);
                      reg866 <= (~|$unsigned((~^(reg839 ? (8'hb4) : (8'ha6)))));
                    end
                  else
                    begin
                      reg865 <= ($unsigned($unsigned($unsigned(reg857))) && ((8'ha6) ?
                          ($unsigned(reg857) < (reg838 ?
                              reg849 : reg858)) : ((forvar847 ?
                                  reg845 : reg840) ?
                              $signed(reg861) : (-forvar837))));
                      reg866 <= $unsigned(($unsigned($unsigned((8'ha9))) > $unsigned(reg857)));
                      reg867 <= $signed(((&(+reg846)) ?
                          forvar851[(2'h3):(2'h3)] : ($unsigned(reg854) && (&reg862))));
                      reg868 <= $unsigned((reg854 ?
                          (~^$unsigned((8'ha6))) : ((~^reg857) << {(8'hb1)})));
                    end
                  for (forvar869 = (1'h0); (forvar869 < (1'h0)); forvar869 = (forvar869 + (1'h1)))
                    begin
                      reg870 <= $unsigned((((8'hae) <= ((8'h9c) ~^ forvar851)) + $signed(wire5[(4'h9):(1'h0)])));
                    end
                  for (forvar871 = (1'h0); (forvar871 < (1'h1)); forvar871 = (forvar871 + (1'h1)))
                    begin
                      reg872 <= (8'ha8);
                      reg873 <= ($signed((forvar864[(3'h4):(3'h4)] == ((8'hb6) ^ wire836))) ?
                          $unsigned(reg853[(1'h0):(1'h0)]) : $unsigned(((wire4 ?
                                  reg859 : wire2) ?
                              $signed((8'had)) : $signed(reg856))));
                      reg874 <= {forvar847};
                      reg875 <= reg859;
                    end
                end
              for (forvar876 = (1'h0); (forvar876 < (1'h1)); forvar876 = (forvar876 + (1'h1)))
                begin
                  if ($unsigned(reg839[(1'h0):(1'h0)]))
                    begin
                      reg877 <= (reg861[(4'h9):(1'h1)] ?
                          (reg840[(3'h6):(2'h3)] ?
                              reg841[(3'h4):(1'h1)] : (-(reg853 ?
                                  reg853 : reg874))) : ({(~|forvar858)} ?
                              ($signed(forvar863) & $signed(reg861)) : ({reg845} ?
                                  {forvar844} : {forvar864})));
                      reg878 <= (~^$unsigned($unsigned((!reg849))));
                    end
                  else
                    begin
                      reg877 <= (^(8'ha3));
                      reg878 <= ((8'ha5) >>> forvar869[(3'h5):(3'h4)]);
                    end
                end
              reg879 <= ((+(reg868[(2'h3):(1'h1)] ?
                      (reg874 | reg841) : forvar851[(3'h4):(2'h2)])) ?
                  reg841 : $signed(reg847[(4'ha):(3'h5)]));
            end
          for (forvar880 = (1'h0); (forvar880 < (2'h3)); forvar880 = (forvar880 + (1'h1)))
            begin
              if (forvar880)
                begin
                  if ($signed($signed({reg878})))
                    begin
                      reg881 <= $unsigned(forvar880);
                    end
                  else
                    begin
                      reg881 <= $unsigned(({$unsigned(reg850)} ^ reg850[(3'h7):(2'h3)]));
                      reg882 <= (+(reg856 != $signed(reg856[(2'h3):(2'h2)])));
                      reg883 <= $signed((^~{(reg844 && reg879)}));
                      reg884 <= ($signed(reg868[(4'hc):(4'hc)]) ?
                          forvar847 : ($unsigned(reg868) ?
                              ((8'ha9) ?
                                  $signed(reg839) : $signed(reg873)) : (8'ha8)));
                    end
                end
              else
                begin
                  if (reg868)
                    begin
                      reg881 <= reg857;
                      reg882 <= (forvar837 > ($signed((wire0 ?
                          reg883 : wire834)) + ((forvar863 & reg867) ?
                          (~forvar864) : (-forvar847))));
                    end
                  else
                    begin
                      reg881 <= $unsigned($signed($signed(reg845[(1'h0):(1'h0)])));
                    end
                  for (forvar883 = (1'h0); (forvar883 < (2'h2)); forvar883 = (forvar883 + (1'h1)))
                    begin
                      reg884 <= ({$signed((reg881 && reg850))} || {$unsigned({reg840})});
                      reg885 <= $signed(reg861);
                      reg886 <= $signed(((+(^reg855)) != ((wire1 ?
                              reg850 : wire836) ?
                          $signed((8'h9e)) : reg849[(1'h0):(1'h0)])));
                    end
                end
              for (forvar887 = (1'h0); (forvar887 < (1'h1)); forvar887 = (forvar887 + (1'h1)))
                begin
                  for (forvar888 = (1'h0); (forvar888 < (1'h1)); forvar888 = (forvar888 + (1'h1)))
                    begin
                      reg889 <= ((|(8'hb0)) ?
                          ({(forvar838 ? reg881 : forvar838)} ^ ({forvar842} ?
                              $signed(wire0) : reg877[(1'h0):(1'h0)])) : ($unsigned(reg886) < reg885[(1'h1):(1'h1)]));
                      reg890 <= (~^{reg843});
                      reg891 <= (!$signed(forvar871));
                    end
                  for (forvar892 = (1'h0); (forvar892 < (2'h3)); forvar892 = (forvar892 + (1'h1)))
                    begin
                      reg893 <= (^~(8'hb3));
                      reg894 <= (forvar869[(3'h5):(2'h3)] <= $unsigned({reg857}));
                      reg895 <= $unsigned($signed((^$signed((8'ha4)))));
                    end
                  if ({$unsigned(($unsigned(reg889) >> (forvar864 ?
                          wire834 : forvar869)))})
                    begin
                      reg896 <= reg875[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg896 <= (~($unsigned((~reg860)) <<< (wire0[(4'he):(4'h8)] & reg860[(1'h0):(1'h0)])));
                      reg897 <= $signed(forvar844[(1'h0):(1'h0)]);
                      reg898 <= $signed(($signed(reg852[(2'h3):(1'h1)]) ?
                          $signed((-reg852)) : ((reg838 ? (8'hb4) : reg897) ?
                              (reg890 - reg849) : $unsigned(forvar887))));
                    end
                  reg899 <= $unsigned($signed((~&wire2[(3'h4):(2'h2)])));
                end
            end
          if ($signed(reg862))
            begin
              reg900 <= (8'hb0);
            end
          else
            begin
              for (forvar900 = (1'h0); (forvar900 < (1'h1)); forvar900 = (forvar900 + (1'h1)))
                begin
                  for (forvar901 = (1'h0); (forvar901 < (1'h0)); forvar901 = (forvar901 + (1'h1)))
                    begin
                      reg902 <= (reg878 - reg844[(2'h2):(1'h0)]);
                      reg903 <= $unsigned(forvar901[(3'h5):(2'h3)]);
                    end
                  reg904 <= ((-reg866[(4'ha):(1'h0)]) ?
                      $unsigned(((reg897 <<< reg855) ?
                          reg861 : $unsigned((8'hac)))) : forvar900);
                  if ({forvar842[(4'hb):(2'h3)]})
                    begin
                      reg905 <= $unsigned(($signed((+reg903)) ?
                          reg899[(5'h10):(4'h9)] : $unsigned({(8'hb4)})));
                      reg906 <= reg858;
                    end
                  else
                    begin
                      reg905 <= (reg848 << {(~$unsigned(reg895))});
                      reg906 <= (forvar864[(3'h6):(1'h0)] ^ $unsigned(forvar838));
                    end
                end
            end
        end
      if ({$unsigned(reg877[(4'hb):(3'h5)])})
        begin
          for (forvar907 = (1'h0); (forvar907 < (2'h2)); forvar907 = (forvar907 + (1'h1)))
            begin
              if ((|reg883[(3'h6):(3'h5)]))
                begin
                  if (forvar869)
                    begin
                      reg908 <= $unsigned(forvar892);
                      reg909 <= reg875[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg908 <= ((($signed(reg840) ^~ (^forvar907)) <= $signed({wire1})) >= reg874[(2'h2):(2'h2)]);
                      reg909 <= ((^~reg873) ?
                          (~^reg856) : forvar888[(2'h2):(2'h2)]);
                      reg910 <= $signed($unsigned(({forvar837} ?
                          ((8'ha4) ? reg881 : forvar864) : reg890)));
                      reg911 <= (forvar864[(3'h7):(3'h5)] ?
                          (&reg857) : reg879[(2'h2):(1'h1)]);
                    end
                  if ($signed(($signed((~reg872)) ^ reg883)))
                    begin
                      reg912 <= ($signed($signed(reg904)) ?
                          (-((8'ha2) ?
                              (reg857 ?
                                  forvar863 : reg841) : {reg852})) : forvar863);
                      reg913 <= $signed(reg874[(2'h3):(1'h1)]);
                      reg914 <= $unsigned($unsigned((reg902[(3'h4):(2'h3)] & reg872)));
                    end
                  else
                    begin
                      reg912 <= ((8'haf) ?
                          $signed(((&(8'hb3)) && (~&reg872))) : (forvar863[(4'hb):(1'h0)] ?
                              (&(wire2 ? (8'hb2) : forvar888)) : (!reg867)));
                    end
                  for (forvar915 = (1'h0); (forvar915 < (2'h3)); forvar915 = (forvar915 + (1'h1)))
                    begin
                      reg916 <= reg838[(3'h6):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar908 = (1'h0); (forvar908 < (1'h0)); forvar908 = (forvar908 + (1'h1)))
                    begin
                      reg909 <= ($unsigned((^{forvar864})) - reg911[(3'h6):(2'h3)]);
                      reg910 <= ((~^($signed(reg859) ?
                              (reg914 ?
                                  reg853 : (8'hab)) : $unsigned(reg875))) ?
                          $signed(((reg885 < reg899) ?
                              $signed(reg875) : (reg853 < reg866))) : forvar863[(3'h5):(1'h0)]);
                      reg911 <= wire3;
                    end
                  if (reg843)
                    begin
                      reg912 <= $unsigned({reg875});
                    end
                  else
                    begin
                      reg912 <= ($signed($unsigned($unsigned(reg865))) >= (($signed(forvar900) ?
                              (reg844 == (8'hb6)) : reg872) ?
                          $signed(reg882) : ((^~reg855) ?
                              (8'hb7) : {(8'hae)})));
                      reg913 <= ($signed((!(!reg865))) != $unsigned(forvar883));
                      reg914 <= $signed((((8'hb6) >>> (reg870 || reg904)) <<< $signed(reg859)));
                    end
                end
              for (forvar917 = (1'h0); (forvar917 < (1'h1)); forvar917 = (forvar917 + (1'h1)))
                begin
                  for (forvar918 = (1'h0); (forvar918 < (2'h2)); forvar918 = (forvar918 + (1'h1)))
                    begin
                      reg919 <= $unsigned({(-(reg885 == (8'h9f)))});
                      reg920 <= $signed(reg908);
                      reg921 <= (-reg886[(3'h4):(2'h2)]);
                    end
                end
              if ((((reg897[(2'h2):(1'h0)] <= $unsigned(reg895)) ?
                      ($unsigned(reg909) & ((8'h9e) && reg844)) : (^((8'ha2) ?
                          forvar917 : reg895))) ?
                  $signed(($signed(reg884) || (reg861 & forvar864))) : forvar863[(4'he):(2'h2)]))
                begin
                  if (reg877[(3'h4):(2'h2)])
                    begin
                      reg922 <= reg894;
                      reg923 <= reg861;
                      reg924 <= $unsigned(($unsigned($unsigned((8'hb5))) ?
                          {(wire834 ? reg914 : reg843)} : reg886));
                    end
                  else
                    begin
                      reg922 <= ({($signed(forvar887) ?
                              $signed(reg849) : reg902)} * $unsigned((8'ha0)));
                    end
                  for (forvar925 = (1'h0); (forvar925 < (1'h0)); forvar925 = (forvar925 + (1'h1)))
                    begin
                      reg926 <= ($signed((8'ha8)) <= $signed($signed(reg878)));
                      reg927 <= {(-reg919[(1'h1):(1'h0)])};
                      reg928 <= ((reg908[(1'h0):(1'h0)] * $unsigned(reg895)) >= {$unsigned($signed(reg872))});
                      reg929 <= (^~({(&reg891)} >= $unsigned((~forvar863))));
                    end
                  if (forvar888)
                    begin
                      reg930 <= reg893[(2'h2):(1'h1)];
                      reg931 <= (reg858[(2'h2):(1'h0)] ?
                          (^~(reg866[(1'h1):(1'h0)] >= ((8'hb2) ?
                              wire834 : (8'hae)))) : ($unsigned(forvar915) ?
                              reg848 : reg894[(3'h6):(2'h2)]));
                    end
                  else
                    begin
                      reg930 <= $unsigned(reg862);
                      reg931 <= reg840;
                      reg932 <= ((($unsigned(reg846) ?
                          $signed((8'hba)) : (reg896 ?
                              reg868 : reg898)) && (~|{reg889})) | reg898);
                    end
                  reg933 <= $unsigned($signed(($signed(reg852) && (~^forvar858))));
                end
              else
                begin
                  for (forvar922 = (1'h0); (forvar922 < (1'h1)); forvar922 = (forvar922 + (1'h1)))
                    begin
                      reg923 <= $signed(forvar917[(3'h6):(3'h6)]);
                      reg924 <= ((^reg922) ?
                          $unsigned(forvar908) : $signed(forvar858));
                      reg925 <= $unsigned($signed((|(&reg930))));
                      reg926 <= ($unsigned($unsigned(((8'hb9) - (8'hac)))) ?
                          forvar871 : $unsigned((^~wire3)));
                    end
                end
              for (forvar934 = (1'h0); (forvar934 < (1'h1)); forvar934 = (forvar934 + (1'h1)))
                begin
                  for (forvar935 = (1'h0); (forvar935 < (1'h0)); forvar935 = (forvar935 + (1'h1)))
                    begin
                      reg936 <= $unsigned($signed($signed($unsigned(reg884))));
                    end
                  for (forvar937 = (1'h0); (forvar937 < (2'h3)); forvar937 = (forvar937 + (1'h1)))
                    begin
                      reg938 <= ($signed($unsigned(reg840[(2'h2):(1'h0)])) || {(reg865 ?
                              $unsigned(wire834) : reg866)});
                    end
                  reg939 <= reg868[(4'he):(1'h0)];
                end
            end
          for (forvar940 = (1'h0); (forvar940 < (2'h2)); forvar940 = (forvar940 + (1'h1)))
            begin
              reg941 <= {(+($unsigned(reg897) & (reg884 | reg873)))};
              for (forvar942 = (1'h0); (forvar942 < (1'h1)); forvar942 = (forvar942 + (1'h1)))
                begin
                  for (forvar943 = (1'h0); (forvar943 < (2'h3)); forvar943 = (forvar943 + (1'h1)))
                    begin
                      reg944 <= forvar837;
                    end
                  if ((reg861[(1'h0):(1'h0)] ?
                      ({(forvar918 > reg928)} ?
                          ((8'had) && $unsigned((8'haf))) : $unsigned(reg928)) : $unsigned((^~$signed(forvar876)))))
                    begin
                      reg945 <= $unsigned(forvar937);
                    end
                  else
                    begin
                      reg945 <= reg903;
                      reg946 <= $signed($unsigned((~$unsigned(forvar935))));
                      reg947 <= reg924[(2'h2):(2'h2)];
                    end
                end
              if (($signed((^(reg927 < reg844))) > (-(forvar883 >= {reg898}))))
                begin
                  if (reg932)
                    begin
                      reg948 <= ({(^~(forvar888 << reg865))} ?
                          ($unsigned((-forvar887)) ?
                              (((8'had) >= reg916) & ((8'hb0) != forvar858)) : forvar937[(2'h2):(1'h1)]) : $unsigned(((reg865 ?
                              (8'hb1) : wire836) ^~ $unsigned(forvar863))));
                      reg949 <= ((^~forvar901[(1'h0):(1'h0)]) * $unsigned(((~|reg897) >> $signed(reg842))));
                    end
                  else
                    begin
                      reg948 <= {(8'hac)};
                    end
                  if ((|(^({(8'h9c)} ? (|wire3) : reg843[(3'h5):(2'h3)]))))
                    begin
                      reg950 <= ($unsigned((8'hb7)) > $unsigned($signed(reg947[(3'h4):(2'h3)])));
                      reg951 <= $signed(reg920);
                      reg952 <= {reg916};
                      reg953 <= (reg861[(2'h3):(2'h2)] ?
                          $signed(forvar907) : $unsigned((^~(reg886 ?
                              reg896 : reg941))));
                    end
                  else
                    begin
                      reg950 <= (reg900 + $signed($signed((8'ha8))));
                      reg951 <= {((8'ha8) >> $unsigned(reg921[(1'h1):(1'h1)]))};
                    end
                  for (forvar954 = (1'h0); (forvar954 < (1'h1)); forvar954 = (forvar954 + (1'h1)))
                    begin
                      reg955 <= reg905;
                      reg956 <= (+forvar915);
                    end
                end
              else
                begin
                  reg948 <= (reg839[(4'he):(3'h4)] <= (($signed(reg906) ~^ reg885) ?
                      $unsigned($unsigned(reg886)) : $unsigned((+reg884))));
                end
              for (forvar957 = (1'h0); (forvar957 < (2'h3)); forvar957 = (forvar957 + (1'h1)))
                begin
                  for (forvar958 = (1'h0); (forvar958 < (2'h3)); forvar958 = (forvar958 + (1'h1)))
                    begin
                      reg959 <= (|wire836);
                    end
                  if ($unsigned($unsigned($signed($unsigned(forvar925)))))
                    begin
                      reg960 <= $unsigned(reg855);
                      reg961 <= (8'hb0);
                      reg962 <= $unsigned(reg889);
                    end
                  else
                    begin
                      reg960 <= forvar925;
                    end
                  for (forvar963 = (1'h0); (forvar963 < (1'h0)); forvar963 = (forvar963 + (1'h1)))
                    begin
                      reg964 <= forvar871[(3'h6):(2'h2)];
                      reg965 <= reg870[(3'h7):(2'h2)];
                      reg966 <= $unsigned($unsigned(forvar917[(3'h4):(3'h4)]));
                      reg967 <= forvar900[(2'h3):(2'h3)];
                    end
                end
            end
        end
      else
        begin
          if ($signed(wire836[(3'h5):(2'h3)]))
            begin
              if (((reg960[(4'hc):(1'h0)] ?
                  reg922 : $unsigned((^~reg960))) <<< forvar871[(4'hb):(3'h5)]))
                begin
                  if ((forvar838[(2'h2):(2'h2)] ?
                      $signed(($signed(reg914) ?
                          (8'h9e) : (~&reg928))) : ((forvar851[(3'h4):(1'h1)] ?
                              reg967 : (reg947 <<< reg955)) ?
                          reg932[(4'ha):(2'h3)] : (reg899 ?
                              {reg922} : (&reg902)))))
                    begin
                      reg907 <= reg875;
                      reg908 <= $unsigned((reg947[(2'h2):(1'h0)] >> $unsigned($signed(reg886))));
                      reg909 <= forvar887;
                    end
                  else
                    begin
                      reg907 <= {(!{$signed(wire0)})};
                    end
                end
              else
                begin
                  for (forvar907 = (1'h0); (forvar907 < (2'h2)); forvar907 = (forvar907 + (1'h1)))
                    begin
                      reg908 <= (forvar871[(4'h8):(3'h7)] != reg936);
                      reg909 <= forvar942;
                      reg910 <= ((reg884 > ((reg932 ? reg841 : wire0) ?
                          forvar864[(2'h2):(2'h2)] : $unsigned(reg965))) == reg857[(3'h5):(1'h1)]);
                      reg911 <= (~^(reg931[(3'h5):(1'h0)] && (~&(reg838 ?
                          forvar863 : (8'ha4)))));
                    end
                end
              for (forvar912 = (1'h0); (forvar912 < (1'h0)); forvar912 = (forvar912 + (1'h1)))
                begin
                  if ((~(|reg924[(2'h3):(2'h3)])))
                    begin
                      reg913 <= {((reg845 >>> reg944[(5'h10):(4'he)]) ?
                              $signed((reg873 << wire836)) : $signed({reg953}))};
                    end
                  else
                    begin
                      reg913 <= $unsigned(reg860);
                      reg914 <= $unsigned($signed((^~(wire2 ?
                          reg919 : reg924))));
                      reg915 <= (((~&reg962) ?
                          {reg875[(3'h4):(1'h1)]} : ($unsigned(reg866) <= $unsigned(reg945))) || (wire3[(1'h1):(1'h1)] ?
                          reg930[(1'h1):(1'h1)] : (forvar954[(1'h1):(1'h0)] ^~ reg848)));
                    end
                  for (forvar916 = (1'h0); (forvar916 < (2'h2)); forvar916 = (forvar916 + (1'h1)))
                    begin
                      reg917 <= (forvar912 >= reg848);
                      reg918 <= $unsigned(reg950[(1'h0):(1'h0)]);
                    end
                end
              if (reg933[(1'h0):(1'h0)])
                begin
                  for (forvar919 = (1'h0); (forvar919 < (2'h3)); forvar919 = (forvar919 + (1'h1)))
                    begin
                      reg920 <= ($signed(reg926) ?
                          (^$signed((reg933 ? (8'hab) : forvar863))) : reg898);
                      reg921 <= (wire836[(3'h5):(1'h1)] <<< (|$unsigned($signed((8'hb6)))));
                    end
                  for (forvar922 = (1'h0); (forvar922 < (1'h0)); forvar922 = (forvar922 + (1'h1)))
                    begin
                      reg923 <= $signed(wire4);
                    end
                  for (forvar924 = (1'h0); (forvar924 < (2'h3)); forvar924 = (forvar924 + (1'h1)))
                    begin
                      reg925 <= (&((^wire3) << (((8'ha6) ?
                          reg904 : (8'hb4)) | forvar957)));
                      reg926 <= reg908;
                      reg927 <= ({reg884[(1'h0):(1'h0)]} > {$unsigned({reg899})});
                    end
                  for (forvar928 = (1'h0); (forvar928 < (1'h0)); forvar928 = (forvar928 + (1'h1)))
                    begin
                      reg929 <= forvar928;
                      reg930 <= $unsigned($unsigned($unsigned({reg854})));
                      reg931 <= reg930[(1'h1):(1'h1)];
                      reg932 <= ($signed(($unsigned((8'h9f)) ?
                          (8'hb8) : $signed(reg919))) >= ({(reg959 ?
                                  forvar892 : forvar880)} ?
                          (forvar871 ?
                              reg908[(3'h5):(2'h3)] : (-(8'hb4))) : forvar963));
                    end
                end
              else
                begin
                  reg919 <= {((8'ha2) ?
                          (reg902[(2'h3):(1'h0)] - $unsigned((8'hb2))) : $signed((forvar864 ?
                              (8'hb3) : wire0)))};
                  for (forvar920 = (1'h0); (forvar920 < (2'h2)); forvar920 = (forvar920 + (1'h1)))
                    begin
                      reg921 <= $unsigned(reg861[(3'h5):(3'h5)]);
                    end
                  if ((((-reg899) ?
                      (8'ha3) : reg847[(3'h7):(1'h1)]) < forvar901[(1'h1):(1'h0)]))
                    begin
                      reg922 <= $signed(reg953[(4'h9):(3'h5)]);
                    end
                  else
                    begin
                      reg922 <= (~^({{reg926}} ?
                          $signed($signed(reg965)) : {$signed(reg951)}));
                      reg923 <= ($signed((wire3[(1'h0):(1'h0)] & (forvar851 ?
                              forvar838 : reg933))) ?
                          (forvar918[(3'h5):(2'h3)] ?
                              $signed($signed(reg961)) : $signed($unsigned(reg903))) : $unsigned({(reg865 ?
                                  reg918 : forvar876)}));
                    end
                  if (reg924[(2'h3):(1'h1)])
                    begin
                      reg924 <= reg855;
                    end
                  else
                    begin
                      reg924 <= $signed((~^$unsigned((wire5 | (8'ha5)))));
                      reg925 <= $unsigned($unsigned($signed((+forvar907))));
                      reg926 <= (|((reg898 ?
                              (forvar851 < (8'hae)) : (reg884 ^~ reg843)) ?
                          $signed(reg920[(4'h8):(3'h4)]) : $signed((reg930 <<< forvar869))));
                    end
                end
              if (reg870)
                begin
                  for (forvar933 = (1'h0); (forvar933 < (1'h1)); forvar933 = (forvar933 + (1'h1)))
                    begin
                      reg934 <= ((~&reg879) * $signed((^~((8'hba) ?
                          reg925 : reg852))));
                    end
                  for (forvar935 = (1'h0); (forvar935 < (2'h2)); forvar935 = (forvar935 + (1'h1)))
                    begin
                      reg936 <= $signed(((&(~reg867)) >>> $unsigned((~|reg886))));
                      reg937 <= forvar858;
                    end
                  for (forvar938 = (1'h0); (forvar938 < (1'h1)); forvar938 = (forvar938 + (1'h1)))
                    begin
                      reg939 <= $signed((((reg889 ? (8'ha2) : forvar858) ?
                              {forvar838} : reg922) ?
                          (~^(reg857 ?
                              forvar901 : reg914)) : (~reg937[(2'h3):(1'h1)])));
                      reg940 <= $unsigned($signed($signed($signed(forvar915))));
                    end
                end
              else
                begin
                  if ($signed(reg885))
                    begin
                      reg933 <= ($signed((|(~^(8'ha7)))) - $unsigned(forvar954));
                      reg934 <= ((((^~(8'hae)) || $signed((8'hb1))) ?
                              reg933 : {(-reg929)}) ?
                          reg965[(4'h8):(2'h3)] : $signed((&(reg890 >> reg882))));
                      reg935 <= reg895;
                    end
                  else
                    begin
                      reg933 <= (+(+((^reg848) ?
                          $unsigned((8'hb9)) : {reg966})));
                      reg934 <= ($signed((~(reg908 ~^ reg964))) || ($signed(((8'had) ?
                          forvar837 : forvar864)) ^~ (8'hb2)));
                      reg935 <= (+($unsigned({(8'ha5)}) ?
                          (^((8'hb3) >> reg928)) : ({wire2} ^ $signed(forvar957))));
                    end
                  if ((reg856 == ($signed((~|reg956)) & ((8'ha5) ?
                      reg924 : reg874[(2'h2):(1'h0)]))))
                    begin
                      reg936 <= (~(((forvar863 ? reg924 : reg898) ?
                              $unsigned(reg903) : reg870) ?
                          ($signed(reg859) || $unsigned((8'hb5))) : ((reg949 <<< wire4) ?
                              (^forvar916) : forvar907)));
                      reg937 <= forvar922;
                      reg938 <= (forvar917 ?
                          wire1 : ($unsigned($signed(reg907)) <<< (|((8'hae) - reg848))));
                      reg939 <= reg941[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg936 <= (8'hb7);
                      reg937 <= ($unsigned({reg925[(3'h5):(1'h1)]}) ^~ $signed($signed($signed((8'hb8)))));
                      reg938 <= wire5[(4'h9):(4'h8)];
                    end
                  if ($signed((^~$unsigned((reg951 ? reg875 : forvar838)))))
                    begin
                      reg940 <= {$unsigned({(forvar869 ? reg917 : (8'hac))})};
                      reg941 <= forvar957;
                      reg942 <= $unsigned((^($unsigned(forvar837) ?
                          (!wire3) : reg924)));
                    end
                  else
                    begin
                      reg940 <= ($signed((^$signed(reg932))) == (8'hb3));
                    end
                end
            end
          else
            begin
              for (forvar907 = (1'h0); (forvar907 < (1'h0)); forvar907 = (forvar907 + (1'h1)))
                begin
                  for (forvar908 = (1'h0); (forvar908 < (2'h3)); forvar908 = (forvar908 + (1'h1)))
                    begin
                      reg909 <= $signed($unsigned({$signed((8'h9c))}));
                      reg910 <= $unsigned(reg845[(3'h4):(2'h3)]);
                    end
                  if (((~&(~|$unsigned(reg874))) - (((reg881 ?
                              (8'hb0) : reg891) ?
                          (^~reg956) : (forvar858 ? reg898 : reg853)) ?
                      (((8'ha4) ? reg883 : reg854) ?
                          forvar924[(2'h3):(1'h0)] : (forvar887 ?
                              reg911 : forvar851)) : $signed((forvar871 ?
                          forvar934 : reg960)))))
                    begin
                      reg911 <= (reg959[(3'h4):(2'h2)] ?
                          reg911[(3'h4):(2'h3)] : $unsigned((reg920[(1'h1):(1'h0)] + reg867)));
                    end
                  else
                    begin
                      reg911 <= (reg838[(3'h6):(2'h3)] ?
                          (($signed((8'h9e)) != {forvar915}) ?
                              (~(~^reg886)) : (!reg960)) : (~&$unsigned({forvar935})));
                    end
                  if ({($unsigned(reg964[(2'h2):(1'h0)]) - forvar922[(2'h2):(1'h1)])})
                    begin
                      reg912 <= $unsigned(reg962[(1'h0):(1'h0)]);
                      reg913 <= reg940[(3'h7):(3'h7)];
                      reg914 <= reg883;
                    end
                  else
                    begin
                      reg912 <= $signed(((!$signed((8'ha1))) <= {(reg946 ?
                              reg894 : (8'ha9))}));
                      reg913 <= forvar933;
                      reg914 <= (~|((reg933[(4'hf):(4'he)] >>> reg859[(1'h0):(1'h0)]) ?
                          $unsigned((reg916 >= reg868)) : {reg961}));
                      reg915 <= reg917;
                    end
                end
              if (forvar963[(4'hb):(3'h6)])
                begin
                  for (forvar916 = (1'h0); (forvar916 < (1'h0)); forvar916 = (forvar916 + (1'h1)))
                    begin
                      reg917 <= ((^$signed({forvar916})) ?
                          (-(8'hba)) : $unsigned((((8'ha2) ?
                              forvar957 : (8'ha3)) * $unsigned(reg895))));
                      reg918 <= forvar922[(3'h6):(3'h6)];
                      reg919 <= reg883;
                      reg920 <= $unsigned($signed((|$unsigned(forvar940))));
                    end
                  for (forvar921 = (1'h0); (forvar921 < (2'h2)); forvar921 = (forvar921 + (1'h1)))
                    begin
                      reg922 <= $signed((+(forvar938[(4'hd):(1'h1)] ?
                          {reg944} : (reg839 <= reg852))));
                    end
                  if ((~reg945[(4'h9):(2'h2)]))
                    begin
                      reg923 <= ($signed($signed(reg881)) ?
                          (^~forvar958[(3'h4):(2'h2)]) : $unsigned($signed((reg945 ?
                              reg884 : reg920))));
                    end
                  else
                    begin
                      reg923 <= ((((reg846 == wire2) * $signed(reg920)) - reg844[(3'h4):(2'h3)]) | {({reg879} & {forvar907})});
                      reg924 <= reg944;
                    end
                end
              else
                begin
                  if ($signed((reg845 ?
                      ({reg941} + $unsigned((8'hb3))) : $unsigned(forvar871))))
                    begin
                      reg916 <= ($unsigned($signed((8'ha9))) + $unsigned({(reg927 ?
                              wire3 : reg855)}));
                      reg917 <= $unsigned({reg895});
                      reg918 <= reg848[(3'h4):(2'h3)];
                      reg919 <= ($signed(((|reg904) ?
                          (!reg946) : $signed(wire2))) != $signed(reg843[(4'h9):(1'h0)]));
                    end
                  else
                    begin
                      reg916 <= ({$signed({reg848})} >>> $signed($signed(((8'hb3) ^ forvar954))));
                    end
                  if ($unsigned((-$signed(reg916[(2'h3):(1'h0)]))))
                    begin
                      reg920 <= ($unsigned((((8'ha7) == forvar887) ?
                              ((8'hba) ~^ reg941) : $unsigned(reg884))) ?
                          {(reg858 ?
                                  reg910[(3'h4):(1'h1)] : {forvar957})} : reg862);
                    end
                  else
                    begin
                      reg920 <= reg915[(2'h3):(2'h2)];
                      reg921 <= {forvar901};
                      reg922 <= {(~^forvar888[(1'h0):(1'h0)])};
                      reg923 <= {{(reg933 ? {forvar851} : forvar851)}};
                    end
                  if ((~^(~^$unsigned(((8'ha1) ? reg939 : (8'ha0))))))
                    begin
                      reg924 <= (8'ha1);
                      reg925 <= (8'hba);
                    end
                  else
                    begin
                      reg924 <= reg956;
                    end
                  reg926 <= (reg922[(3'h4):(1'h0)] ?
                      (reg886 | {$signed((8'h9e))}) : $unsigned(reg854));
                end
              for (forvar927 = (1'h0); (forvar927 < (1'h0)); forvar927 = (forvar927 + (1'h1)))
                begin
                  for (forvar928 = (1'h0); (forvar928 < (1'h0)); forvar928 = (forvar928 + (1'h1)))
                    begin
                      reg929 <= reg959[(3'h4):(1'h0)];
                      reg930 <= ($unsigned(reg844) > (8'hb6));
                    end
                  if ({($signed($unsigned(reg894)) ?
                          $unsigned($signed(reg900)) : (~&(~wire5)))})
                    begin
                      reg931 <= reg877[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg931 <= (!(+$unsigned((reg870 >>> reg895))));
                    end
                end
            end
          if (reg896)
            begin
              for (forvar943 = (1'h0); (forvar943 < (2'h2)); forvar943 = (forvar943 + (1'h1)))
                begin
                  for (forvar944 = (1'h0); (forvar944 < (1'h0)); forvar944 = (forvar944 + (1'h1)))
                    begin
                      reg945 <= ($signed(forvar921) ?
                          $unsigned(((reg912 ?
                              (8'hac) : forvar912) >>> wire836[(4'h8):(3'h7)])) : (($unsigned(reg846) == (|wire2)) >>> ((^~(8'hba)) ?
                              wire0[(4'h8):(3'h5)] : reg860)));
                    end
                  for (forvar946 = (1'h0); (forvar946 < (1'h1)); forvar946 = (forvar946 + (1'h1)))
                    begin
                      reg947 <= (reg895[(2'h2):(1'h1)] ?
                          forvar940[(1'h1):(1'h1)] : ($unsigned((~^reg952)) - (forvar883[(2'h3):(2'h3)] >>> (reg914 ^ reg940))));
                    end
                  reg948 <= $signed($signed($signed(wire5)));
                end
            end
          else
            begin
              if (reg841)
                begin
                  if (reg886[(2'h2):(2'h2)])
                    begin
                      reg943 <= forvar871[(2'h3):(2'h3)];
                      reg944 <= ($signed($unsigned($signed((8'h9c)))) ?
                          ({reg934} ?
                              $unsigned((reg936 ^~ reg904)) : $signed(forvar954[(2'h2):(2'h2)])) : reg899);
                      reg945 <= reg838;
                      reg946 <= $unsigned(reg945);
                    end
                  else
                    begin
                      reg943 <= reg854;
                      reg944 <= $signed((8'hba));
                      reg945 <= $signed({$unsigned($unsigned(reg923))});
                    end
                  for (forvar947 = (1'h0); (forvar947 < (2'h2)); forvar947 = (forvar947 + (1'h1)))
                    begin
                      reg948 <= (forvar880 ?
                          $signed(((~(8'hac)) || $unsigned(forvar915))) : (-(~|((8'ha5) ?
                              forvar954 : wire3))));
                      reg949 <= reg915[(3'h4):(3'h4)];
                      reg950 <= $unsigned({(forvar938 ?
                              (reg862 ? reg910 : reg895) : (~^reg933))});
                    end
                  reg951 <= (~^(reg878[(2'h2):(2'h2)] && forvar900[(1'h1):(1'h0)]));
                  if ($signed({({(8'hb0)} ? $unsigned(reg950) : reg898)}))
                    begin
                      reg952 <= forvar864[(4'h8):(3'h5)];
                      reg953 <= (&$unsigned((!$unsigned(forvar924))));
                      reg954 <= forvar842[(4'ha):(2'h3)];
                    end
                  else
                    begin
                      reg952 <= $unsigned(($unsigned({reg961}) - forvar847));
                      reg953 <= {reg908};
                      reg954 <= $unsigned($unsigned($signed(((8'hac) ^ reg929))));
                    end
                end
              else
                begin
                  reg943 <= reg870[(3'h4):(3'h4)];
                  for (forvar944 = (1'h0); (forvar944 < (1'h1)); forvar944 = (forvar944 + (1'h1)))
                    begin
                      reg945 <= $unsigned($signed((!(!reg865))));
                      reg946 <= (~|forvar943[(3'h5):(3'h5)]);
                      reg947 <= $signed(((reg889 & (^reg847)) ?
                          reg954[(4'h8):(2'h3)] : (^~$signed(reg896))));
                    end
                  for (forvar948 = (1'h0); (forvar948 < (2'h3)); forvar948 = (forvar948 + (1'h1)))
                    begin
                      reg949 <= reg896[(4'hb):(3'h6)];
                      reg950 <= {reg949[(2'h3):(1'h0)]};
                      reg951 <= $signed((reg927 ~^ $signed(forvar922)));
                    end
                  if (reg959[(2'h3):(1'h0)])
                    begin
                      reg952 <= $signed({{(reg902 ? (8'ha3) : (8'hb4))}});
                      reg953 <= wire5;
                    end
                  else
                    begin
                      reg952 <= (reg859[(2'h2):(1'h0)] | $signed(wire1));
                    end
                end
              for (forvar955 = (1'h0); (forvar955 < (2'h2)); forvar955 = (forvar955 + (1'h1)))
                begin
                  for (forvar956 = (1'h0); (forvar956 < (1'h1)); forvar956 = (forvar956 + (1'h1)))
                    begin
                      reg957 <= $unsigned(forvar963[(3'h7):(1'h0)]);
                      reg958 <= ({forvar938} > {reg945[(1'h0):(1'h0)]});
                    end
                  for (forvar959 = (1'h0); (forvar959 < (1'h0)); forvar959 = (forvar959 + (1'h1)))
                    begin
                      reg960 <= (($signed($signed(reg900)) || forvar888) ?
                          reg857 : reg883[(2'h3):(1'h0)]);
                    end
                  if ((~|(^~reg961[(4'h9):(3'h6)])))
                    begin
                      reg961 <= $unsigned((-forvar946));
                      reg962 <= wire0[(4'hc):(3'h6)];
                    end
                  else
                    begin
                      reg961 <= {(8'ha1)};
                      reg962 <= ((reg891[(2'h3):(2'h3)] ?
                              (8'h9f) : $unsigned($signed(forvar942))) ?
                          ($signed(((8'ha1) <<< forvar924)) << $signed(reg966)) : $unsigned(reg946[(1'h0):(1'h0)]));
                      reg963 <= (^~$signed($unsigned(reg946[(1'h0):(1'h0)])));
                      reg964 <= (((8'hb3) ?
                          reg943 : forvar869) >> reg938[(1'h1):(1'h1)]);
                    end
                end
            end
          for (forvar965 = (1'h0); (forvar965 < (1'h0)); forvar965 = (forvar965 + (1'h1)))
            begin
              for (forvar966 = (1'h0); (forvar966 < (1'h1)); forvar966 = (forvar966 + (1'h1)))
                begin
                  for (forvar967 = (1'h0); (forvar967 < (2'h3)); forvar967 = (forvar967 + (1'h1)))
                    begin
                      reg968 <= forvar915;
                    end
                end
            end
          for (forvar969 = (1'h0); (forvar969 < (2'h3)); forvar969 = (forvar969 + (1'h1)))
            begin
              if ((8'haf))
                begin
                  if ((8'h9e))
                    begin
                      reg970 <= $unsigned(reg950);
                      reg971 <= {forvar837[(4'ha):(3'h4)]};
                    end
                  else
                    begin
                      reg970 <= $unsigned($signed(forvar946[(2'h2):(1'h1)]));
                      reg971 <= $signed(forvar958);
                      reg972 <= ($signed(reg866) ?
                          $unsigned(forvar925[(4'h9):(3'h4)]) : (^(forvar948 >>> (+(8'had)))));
                      reg973 <= reg971;
                    end
                  reg974 <= reg854[(2'h2):(2'h2)];
                  for (forvar975 = (1'h0); (forvar975 < (2'h2)); forvar975 = (forvar975 + (1'h1)))
                    begin
                      reg976 <= forvar959[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  reg970 <= ((-($signed(forvar948) ?
                      reg976 : (forvar863 ?
                          (8'h9e) : reg870))) > (($unsigned(forvar917) ?
                      ((8'hb3) <= reg960) : reg954) >>> $signed((forvar916 ?
                      reg948 : forvar943))));
                  for (forvar971 = (1'h0); (forvar971 < (2'h3)); forvar971 = (forvar971 + (1'h1)))
                    begin
                      reg972 <= $unsigned($signed(((reg891 != forvar858) ?
                          (!(8'had)) : (|reg904))));
                      reg973 <= $unsigned(($signed($signed(wire1)) + $signed(reg914[(4'hb):(1'h1)])));
                      reg974 <= (~reg944);
                      reg975 <= $unsigned((~&((~|forvar920) << {reg939})));
                    end
                  reg976 <= (~^(&($unsigned((8'ha7)) ?
                      $signed(wire3) : (reg952 ? reg886 : (8'hb8)))));
                end
            end
        end
      if (($unsigned({(~(8'hb8))}) >>> (((forvar901 <<< forvar880) ?
          $unsigned(reg925) : forvar967[(1'h1):(1'h0)]) * forvar863[(4'ha):(2'h2)])))
        begin
          if ((-($unsigned((-reg905)) ?
              ((reg972 ^~ (8'ha8)) >= (forvar925 ?
                  forvar955 : reg955)) : $unsigned($signed(forvar933)))))
            begin
              if (((^($unsigned(forvar963) ?
                      $signed((8'ha2)) : (reg953 <<< wire4))) ?
                  (^~({reg972} - (reg919 ?
                      reg843 : reg844))) : $signed((((8'h9e) << reg874) ?
                      (reg973 ? reg841 : forvar928) : reg945[(3'h5):(1'h1)]))))
                begin
                  if (($unsigned(reg946) ?
                      $unsigned($signed((|reg973))) : $unsigned(reg944[(4'hf):(4'h8)])))
                    begin
                      reg977 <= forvar900[(2'h2):(1'h0)];
                      reg978 <= $unsigned({$unsigned({forvar954})});
                      reg979 <= (^~(forvar863[(3'h7):(2'h2)] >= $signed((reg865 && reg922))));
                    end
                  else
                    begin
                      reg977 <= (forvar958[(3'h4):(2'h2)] ?
                          (($unsigned(forvar922) ? {reg906} : forvar869) ?
                              (reg944[(4'hf):(2'h3)] ~^ (forvar888 * (8'haa))) : reg971) : $signed(((reg963 ?
                                  reg878 : reg940) ?
                              forvar858[(3'h5):(2'h3)] : reg861)));
                      reg978 <= $signed(reg900);
                      reg979 <= (forvar919[(1'h1):(1'h0)] ?
                          $signed($signed((forvar933 <<< reg912))) : $signed(forvar946));
                    end
                  reg980 <= (8'haf);
                end
              else
                begin
                  if (($signed(forvar869[(3'h7):(1'h1)]) ?
                      (reg841[(4'hb):(1'h1)] ?
                          reg955 : {(reg847 * reg877)}) : reg855[(3'h7):(1'h1)]))
                    begin
                      reg977 <= reg922;
                      reg978 <= wire0[(4'he):(4'hb)];
                      reg979 <= forvar871;
                      reg980 <= (~forvar946[(4'h8):(3'h7)]);
                    end
                  else
                    begin
                      reg977 <= $signed($unsigned((+$unsigned(reg949))));
                      reg978 <= $signed((reg879 ?
                          (reg894 || $signed(forvar965)) : $unsigned(reg870[(3'h4):(2'h2)])));
                      reg979 <= $signed({$signed(((8'hae) ?
                              (8'hae) : reg875))});
                      reg980 <= (^(^((reg956 ?
                          reg840 : (8'hb0)) - reg847[(4'ha):(4'h8)])));
                    end
                  for (forvar981 = (1'h0); (forvar981 < (2'h3)); forvar981 = (forvar981 + (1'h1)))
                    begin
                      reg982 <= ($unsigned($unsigned((reg944 ?
                          forvar956 : forvar927))) ^ ($signed((forvar958 ?
                              reg899 : (8'hab))) ?
                          forvar938[(5'h10):(4'hc)] : $unsigned($signed(reg970))));
                      reg983 <= ($signed((|reg902[(2'h2):(1'h1)])) || $signed(((reg967 ?
                              forvar954 : forvar957) ?
                          forvar933 : reg976[(1'h1):(1'h0)])));
                      reg984 <= $unsigned(reg857);
                      reg985 <= reg941;
                    end
                  for (forvar986 = (1'h0); (forvar986 < (1'h0)); forvar986 = (forvar986 + (1'h1)))
                    begin
                      reg987 <= reg966[(4'hc):(4'hb)];
                    end
                end
              if ((8'h9c))
                begin
                  if ({(((reg918 ? forvar863 : forvar924) ^~ (reg870 ?
                              forvar959 : reg937)) ?
                          (^~(-(8'hb8))) : reg843)})
                    begin
                      reg988 <= $signed((($signed(wire4) == reg915[(1'h0):(1'h0)]) ?
                          (reg926[(4'ha):(4'h9)] == $signed(reg838)) : forvar900[(2'h2):(1'h1)]));
                      reg989 <= (((8'ha4) <= $signed($signed(reg927))) ^~ reg974);
                      reg990 <= reg933[(3'h4):(2'h3)];
                      reg991 <= reg975[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg988 <= reg945;
                    end
                  for (forvar992 = (1'h0); (forvar992 < (2'h2)); forvar992 = (forvar992 + (1'h1)))
                    begin
                      reg993 <= reg922;
                      reg994 <= {reg845[(3'h4):(1'h1)]};
                    end
                  for (forvar995 = (1'h0); (forvar995 < (1'h0)); forvar995 = (forvar995 + (1'h1)))
                    begin
                      reg996 <= reg862;
                      reg997 <= reg916;
                      reg998 <= $signed(((reg951[(1'h0):(1'h0)] ?
                          (!reg854) : ((8'hb2) ?
                              (8'hb3) : forvar992)) == reg865[(1'h0):(1'h0)]));
                    end
                  for (forvar999 = (1'h0); (forvar999 < (1'h0)); forvar999 = (forvar999 + (1'h1)))
                    begin
                      reg1000 <= (!forvar947[(3'h4):(1'h1)]);
                      reg1001 <= $signed((~&reg938));
                    end
                end
              else
                begin
                  if (reg898[(1'h0):(1'h0)])
                    begin
                      reg988 <= $unsigned({reg940});
                      reg989 <= ((forvar847[(3'h7):(2'h2)] & $signed($unsigned(forvar958))) >> {((forvar901 > forvar943) == {reg940})});
                      reg990 <= $unsigned($unsigned(((~&forvar995) > ((8'ha7) && reg910))));
                    end
                  else
                    begin
                      reg988 <= ({$signed(((8'hb1) ? forvar966 : reg917))} ?
                          ($unsigned($signed((8'h9d))) == $unsigned($unsigned((8'h9d)))) : {reg842});
                      reg989 <= reg852;
                    end
                  if (((+$unsigned((reg936 ? reg840 : forvar999))) ?
                      reg908 : reg932))
                    begin
                      reg991 <= $unsigned((({forvar837} ^ reg968) - reg861[(3'h6):(3'h6)]));
                      reg992 <= {reg994};
                      reg993 <= $signed(((~&$unsigned((8'hb3))) ?
                          (-(reg907 && forvar883)) : reg890[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg991 <= (($signed({(8'ha7)}) ?
                          $unsigned(reg925) : reg961[(4'ha):(3'h6)]) & reg845);
                      reg992 <= forvar837;
                    end
                  for (forvar994 = (1'h0); (forvar994 < (1'h0)); forvar994 = (forvar994 + (1'h1)))
                    begin
                      reg995 <= (forvar948[(3'h4):(3'h4)] ?
                          forvar946[(4'hc):(4'h8)] : {{$unsigned(reg906)}});
                      reg996 <= $unsigned(($unsigned($signed(reg878)) ?
                          ($unsigned((8'haf)) ?
                              (reg872 - reg968) : (~|reg941)) : $signed(reg898[(1'h0):(1'h0)])));
                      reg997 <= ($unsigned(reg852[(4'h8):(3'h6)]) ?
                          $signed($signed($unsigned((8'ha1)))) : $signed((~|{forvar918})));
                    end
                  if ($signed(forvar933))
                    begin
                      reg998 <= $signed(($signed($signed(forvar999)) > (!((8'ha8) >> reg900))));
                      reg999 <= $unsigned(forvar851[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg998 <= (~^(reg938[(4'h9):(3'h6)] >>> $unsigned((reg939 ?
                          reg955 : reg855))));
                      reg999 <= ({reg997[(4'h9):(3'h4)]} ?
                          $signed(((&forvar922) ?
                              (forvar942 ^~ forvar999) : $signed(reg917))) : (~^((forvar943 ?
                                  (8'ha4) : reg872) ?
                              (^(8'hb2)) : reg849)));
                    end
                end
              if (reg938[(1'h1):(1'h1)])
                begin
                  for (forvar1002 = (1'h0); (forvar1002 < (2'h2)); forvar1002 = (forvar1002 + (1'h1)))
                    begin
                      reg1003 <= $unsigned((forvar994[(1'h0):(1'h0)] - $signed(reg935[(2'h2):(1'h1)])));
                    end
                  if (reg980)
                    begin
                      reg1004 <= $signed(($unsigned((|reg964)) || (|reg999[(2'h3):(2'h3)])));
                      reg1005 <= (reg891 ?
                          {((forvar954 <<< reg938) ?
                                  (reg992 & reg858) : reg988[(3'h7):(1'h0)])} : {(-reg913[(1'h1):(1'h0)])});
                      reg1006 <= reg935;
                    end
                  else
                    begin
                      reg1004 <= $unsigned((reg980 ?
                          (+$signed(reg904)) : ((forvar981 <<< forvar925) == reg870)));
                      reg1005 <= reg922;
                    end
                  for (forvar1007 = (1'h0); (forvar1007 < (2'h3)); forvar1007 = (forvar1007 + (1'h1)))
                    begin
                      reg1008 <= $signed(reg918);
                      reg1009 <= {$unsigned(reg848)};
                    end
                  for (forvar1010 = (1'h0); (forvar1010 < (1'h1)); forvar1010 = (forvar1010 + (1'h1)))
                    begin
                      reg1011 <= ((((-reg1004) ^ ((8'had) ?
                          reg996 : forvar957)) | (~|(reg846 ?
                          reg953 : forvar837))) << (((|forvar1002) ?
                          (reg1001 | reg911) : forvar869) || reg908[(3'h7):(2'h3)]));
                    end
                end
              else
                begin
                  for (forvar1002 = (1'h0); (forvar1002 < (2'h2)); forvar1002 = (forvar1002 + (1'h1)))
                    begin
                      reg1003 <= reg957;
                      reg1004 <= $unsigned((8'ha1));
                    end
                  for (forvar1005 = (1'h0); (forvar1005 < (2'h2)); forvar1005 = (forvar1005 + (1'h1)))
                    begin
                      reg1006 <= (8'h9f);
                      reg1007 <= (|$signed((~^((8'hb3) ? forvar924 : reg997))));
                      reg1008 <= $signed((reg940 <= forvar958));
                      reg1009 <= $signed((^(-reg995[(3'h4):(2'h3)])));
                    end
                  if (reg977[(1'h0):(1'h0)])
                    begin
                      reg1010 <= (reg877 ^~ (((reg900 ?
                          (8'ha2) : reg852) << $signed(reg838)) * $signed((forvar892 ?
                          reg889 : reg930))));
                      reg1011 <= {(($unsigned(reg857) ?
                                  reg948[(3'h4):(1'h1)] : (reg963 ?
                                      reg856 : (8'ha8))) ?
                              (+(reg991 ? reg953 : reg983)) : ((reg962 ?
                                  reg982 : reg1011) != reg939))};
                      reg1012 <= (((forvar927[(3'h6):(3'h5)] <= $unsigned(reg972)) ~^ reg949[(2'h3):(1'h0)]) ^ (+(forvar916[(1'h0):(1'h0)] < reg854)));
                      reg1013 <= $unsigned((^~{((8'hb1) ? reg980 : reg883)}));
                    end
                  else
                    begin
                      reg1010 <= reg890[(2'h2):(1'h0)];
                      reg1011 <= (+(~&{(reg896 == reg857)}));
                      reg1012 <= (forvar912 + (($signed(forvar869) ?
                          {reg865} : (reg881 ?
                              (8'ha9) : (8'ha9))) ^~ {forvar924}));
                    end
                  for (forvar1014 = (1'h0); (forvar1014 < (2'h2)); forvar1014 = (forvar1014 + (1'h1)))
                    begin
                      reg1015 <= reg953[(4'ha):(4'h8)];
                    end
                end
            end
          else
            begin
              for (forvar977 = (1'h0); (forvar977 < (2'h3)); forvar977 = (forvar977 + (1'h1)))
                begin
                  for (forvar978 = (1'h0); (forvar978 < (2'h3)); forvar978 = (forvar978 + (1'h1)))
                    begin
                      reg979 <= $signed(reg909[(4'hc):(4'h8)]);
                      reg980 <= {(reg961 ?
                              (reg964 ?
                                  reg970 : reg921) : reg984[(3'h7):(2'h3)])};
                    end
                end
            end
          reg1016 <= $unsigned((reg949[(1'h0):(1'h0)] <<< $unsigned($unsigned(reg995))));
          reg1017 <= forvar838;
        end
      else
        begin
          for (forvar977 = (1'h0); (forvar977 < (1'h0)); forvar977 = (forvar977 + (1'h1)))
            begin
              for (forvar978 = (1'h0); (forvar978 < (1'h0)); forvar978 = (forvar978 + (1'h1)))
                begin
                  for (forvar979 = (1'h0); (forvar979 < (2'h2)); forvar979 = (forvar979 + (1'h1)))
                    begin
                      reg980 <= $signed(((8'ha1) ^ $signed(reg919)));
                      reg981 <= ((reg996[(3'h5):(1'h1)] ?
                          (~^(~^forvar978)) : $unsigned((forvar901 + reg1011))) || reg867[(1'h1):(1'h1)]);
                      reg982 <= (8'hb4);
                      reg983 <= $signed($signed(({reg915} ?
                          (reg933 > (8'h9e)) : (reg952 ? reg944 : forvar978))));
                    end
                end
              if ((~^$unsigned((-(reg954 <= reg855)))))
                begin
                  for (forvar984 = (1'h0); (forvar984 < (1'h0)); forvar984 = (forvar984 + (1'h1)))
                    begin
                      reg985 <= ((+forvar880[(1'h1):(1'h0)]) ?
                          (reg862 ?
                              $signed($unsigned(reg1000)) : forvar946) : $unsigned($unsigned((reg1016 ?
                              forvar940 : reg922))));
                      reg986 <= ((forvar924 >>> $signed({forvar838})) ?
                          (((reg862 ? reg989 : reg843) ?
                                  $unsigned(forvar883) : (^~(8'h9e))) ?
                              $unsigned(reg939[(3'h6):(2'h3)]) : $unsigned($unsigned(forvar954))) : {forvar966[(3'h5):(2'h3)]});
                      reg987 <= reg988[(2'h3):(2'h3)];
                    end
                  reg988 <= {reg900};
                  reg989 <= $signed($unsigned($signed(((8'ha4) ?
                      (8'h9d) : reg1015))));
                  for (forvar990 = (1'h0); (forvar990 < (1'h0)); forvar990 = (forvar990 + (1'h1)))
                    begin
                      reg991 <= forvar955;
                    end
                end
              else
                begin
                  for (forvar984 = (1'h0); (forvar984 < (2'h2)); forvar984 = (forvar984 + (1'h1)))
                    begin
                      reg985 <= {((&(forvar942 & reg899)) || wire834)};
                    end
                end
            end
          for (forvar992 = (1'h0); (forvar992 < (2'h3)); forvar992 = (forvar992 + (1'h1)))
            begin
              for (forvar993 = (1'h0); (forvar993 < (2'h2)); forvar993 = (forvar993 + (1'h1)))
                begin
                  for (forvar994 = (1'h0); (forvar994 < (1'h1)); forvar994 = (forvar994 + (1'h1)))
                    begin
                      reg995 <= ($signed(reg900[(4'hf):(4'hd)]) ?
                          $unsigned($unsigned({(8'hb4)})) : $signed(forvar1014[(2'h2):(1'h0)]));
                      reg996 <= (wire4[(1'h0):(1'h0)] ?
                          reg983 : {(reg893 & forvar876)});
                      reg997 <= reg962;
                    end
                  for (forvar998 = (1'h0); (forvar998 < (2'h3)); forvar998 = (forvar998 + (1'h1)))
                    begin
                      reg999 <= $unsigned($unsigned($signed($unsigned((8'ha0)))));
                      reg1000 <= $unsigned((|$signed((reg987 ?
                          reg956 : reg859))));
                    end
                  if ((~|$unsigned(($unsigned(reg941) ?
                      (!reg854) : (^(8'ha5))))))
                    begin
                      reg1001 <= ((({reg839} ^~ reg850[(3'h4):(1'h0)]) ?
                              {(forvar921 ?
                                      reg932 : forvar933)} : $signed(((8'ha6) - reg883))) ?
                          (~^$signed(reg924)) : $signed($unsigned((&reg978))));
                      reg1002 <= {reg905[(3'h5):(2'h3)]};
                      reg1003 <= $signed(reg981);
                      reg1004 <= ((^reg1008) ?
                          ((~$signed(forvar984)) <<< reg1007) : $signed(($signed((8'hb8)) ?
                              $signed(wire3) : (8'ha8))));
                    end
                  else
                    begin
                      reg1001 <= $signed(reg991);
                      reg1002 <= reg988;
                      reg1003 <= forvar915;
                    end
                  reg1005 <= (($unsigned((forvar935 != reg915)) < forvar948) ?
                      $signed((~|forvar916)) : $unsigned(reg948));
                end
              if ((forvar863 == forvar883[(1'h1):(1'h1)]))
                begin
                  if ({(((~|reg972) ~^ (^~(8'ha1))) ?
                          ((~^forvar900) ?
                              reg1007 : (reg924 >>> reg914)) : reg998)})
                    begin
                      reg1006 <= (reg905 ?
                          forvar907[(2'h2):(2'h2)] : ({reg926} ?
                              $unsigned($signed(reg882)) : $unsigned($signed(forvar928))));
                      reg1007 <= $unsigned($signed(($unsigned(forvar921) == (~|reg947))));
                    end
                  else
                    begin
                      reg1006 <= $signed($unsigned(reg982[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  if ((((reg877[(2'h3):(2'h2)] ?
                          (|reg950) : (reg856 >= forvar851)) ?
                      $unsigned((reg954 > reg987)) : $signed(reg995[(1'h1):(1'h1)])) >= (($unsigned(reg950) << {reg860}) ?
                      $signed(forvar1007) : $unsigned(reg895[(2'h3):(2'h2)]))))
                    begin
                      reg1006 <= (~|(($signed(forvar956) >>> $unsigned(reg955)) ?
                          $unsigned((reg972 ?
                              reg1010 : reg874)) : (forvar942[(3'h7):(2'h2)] ?
                              $signed((8'hae)) : $signed((8'h9d)))));
                      reg1007 <= ({(~^reg904[(2'h3):(2'h2)])} ~^ $unsigned((^~$unsigned(reg998))));
                      reg1008 <= (wire0 ?
                          $unsigned(reg1011[(4'hf):(1'h0)]) : forvar838);
                      reg1009 <= reg1012;
                    end
                  else
                    begin
                      reg1006 <= (|$unsigned(((forvar883 ?
                              forvar958 : reg1006) ?
                          (~&(8'haa)) : (forvar864 ? reg975 : (8'hb5)))));
                      reg1007 <= ($signed(({forvar916} ?
                          (forvar943 && forvar938) : wire4[(2'h2):(1'h0)])) >= forvar986);
                      reg1008 <= ($unsigned(forvar887) ?
                          ($unsigned({reg928}) <<< $signed(forvar994[(4'h8):(2'h3)])) : (reg853[(1'h0):(1'h0)] <= $signed($unsigned(reg956))));
                    end
                  reg1010 <= (reg1000[(1'h1):(1'h1)] ?
                      (((forvar888 != forvar938) <<< $unsigned((8'ha2))) > $unsigned((reg989 == (8'hae)))) : forvar907[(2'h2):(1'h0)]);
                  for (forvar1011 = (1'h0); (forvar1011 < (1'h1)); forvar1011 = (forvar1011 + (1'h1)))
                    begin
                      reg1012 <= $unsigned($signed(forvar1007));
                    end
                  for (forvar1013 = (1'h0); (forvar1013 < (1'h0)); forvar1013 = (forvar1013 + (1'h1)))
                    begin
                      reg1014 <= $unsigned((-$unsigned(reg1015)));
                      reg1015 <= $unsigned((reg984[(3'h5):(2'h2)] | (+forvar917)));
                      reg1016 <= (reg873 ?
                          (!$unsigned((8'hb1))) : ((&(|(8'h9c))) & reg978[(1'h1):(1'h1)]));
                      reg1017 <= $unsigned({$unsigned($signed((8'ha2)))});
                    end
                end
              if ((reg856 ?
                  reg861[(1'h0):(1'h0)] : ($signed((forvar1007 * reg939)) <= $signed($unsigned(reg1005)))))
                begin
                  for (forvar1018 = (1'h0); (forvar1018 < (1'h0)); forvar1018 = (forvar1018 + (1'h1)))
                    begin
                      reg1019 <= (forvar901[(2'h2):(1'h0)] ?
                          (~|forvar907) : forvar1018);
                      reg1020 <= (&$unsigned((|{reg927})));
                      reg1021 <= (|(($signed(forvar858) ^~ (forvar880 ?
                              forvar971 : (8'ha2))) ?
                          $signed($signed(reg906)) : $unsigned((reg953 ?
                              reg897 : reg953))));
                    end
                  if ($unsigned((+($signed(forvar1010) ~^ (~|(8'ha8))))))
                    begin
                      reg1022 <= $signed({forvar851});
                      reg1023 <= reg915[(1'h0):(1'h0)];
                      reg1024 <= $signed(((^~$unsigned(reg918)) * ($unsigned(reg900) >= $unsigned(reg999))));
                      reg1025 <= $signed((+reg931));
                    end
                  else
                    begin
                      reg1022 <= (($unsigned(((8'h9e) == reg936)) ?
                              reg915 : ((~forvar869) ?
                                  $unsigned(forvar901) : forvar967[(2'h2):(1'h0)])) ?
                          forvar880 : ($unsigned((+reg1005)) ?
                              (8'hb1) : (!reg967[(3'h5):(1'h0)])));
                      reg1023 <= (reg900[(3'h4):(2'h3)] | (8'hb8));
                      reg1024 <= (^~$unsigned($signed((8'ha9))));
                      reg1025 <= ((|((8'h9d) ?
                              reg986[(2'h2):(1'h1)] : reg850[(3'h6):(3'h4)])) ?
                          ({$unsigned(reg981)} ?
                              ($signed(forvar925) ?
                                  $unsigned(reg995) : (~|reg1025)) : $unsigned($signed(forvar965))) : ((8'ha4) ?
                              reg953[(4'hb):(4'h9)] : (-forvar959[(2'h2):(1'h1)])));
                    end
                  if ((~&(^((8'ha2) <<< (reg1009 ? reg855 : forvar1018)))))
                    begin
                      reg1026 <= ($signed($signed($signed(reg909))) ?
                          reg968 : $unsigned($signed((reg936 ?
                              reg991 : reg873))));
                      reg1027 <= ($unsigned($signed($unsigned(reg954))) | $unsigned($unsigned(reg959[(4'hc):(4'hb)])));
                      reg1028 <= reg945;
                      reg1029 <= ($unsigned($unsigned({(8'hb8)})) - reg1011[(4'hf):(1'h1)]);
                    end
                  else
                    begin
                      reg1026 <= {(forvar920 ?
                              $signed((~^reg962)) : (reg914 >>> (~reg981)))};
                    end
                end
              else
                begin
                  for (forvar1018 = (1'h0); (forvar1018 < (1'h0)); forvar1018 = (forvar1018 + (1'h1)))
                    begin
                      reg1019 <= (reg1006[(4'h8):(3'h5)] + $signed(({reg907} - (~reg934))));
                      reg1020 <= $unsigned((forvar838[(1'h0):(1'h0)] != (~&reg945)));
                      reg1021 <= ($signed((reg896[(1'h1):(1'h1)] + (reg979 && forvar994))) ?
                          $signed((!(|(8'hb3)))) : $signed(reg996[(4'ha):(2'h3)]));
                    end
                  for (forvar1022 = (1'h0); (forvar1022 < (2'h3)); forvar1022 = (forvar1022 + (1'h1)))
                    begin
                      reg1023 <= (8'h9d);
                    end
                  for (forvar1024 = (1'h0); (forvar1024 < (2'h3)); forvar1024 = (forvar1024 + (1'h1)))
                    begin
                      reg1025 <= (8'haf);
                      reg1026 <= ({((~reg1000) >> {reg882})} <= reg1007[(3'h6):(1'h1)]);
                      reg1027 <= ((reg972[(2'h3):(2'h3)] & ((reg896 ?
                          reg936 : reg878) ~^ (~reg896))) ^~ (($signed(forvar959) ?
                          (reg938 ? reg986 : forvar880) : (forvar955 ?
                              reg872 : reg914)) >= $signed(forvar892)));
                    end
                  for (forvar1028 = (1'h0); (forvar1028 < (2'h2)); forvar1028 = (forvar1028 + (1'h1)))
                    begin
                      reg1029 <= $signed(reg1015[(4'h8):(1'h1)]);
                      reg1030 <= reg1020;
                      reg1031 <= {reg1023[(3'h7):(3'h5)]};
                    end
                end
              for (forvar1032 = (1'h0); (forvar1032 < (2'h2)); forvar1032 = (forvar1032 + (1'h1)))
                begin
                  for (forvar1033 = (1'h0); (forvar1033 < (2'h3)); forvar1033 = (forvar1033 + (1'h1)))
                    begin
                      reg1034 <= reg981;
                      reg1035 <= reg908[(3'h4):(2'h3)];
                      reg1036 <= ($unsigned(reg1012[(4'hf):(4'hd)]) == $unsigned($signed((reg991 ?
                          (8'had) : forvar925))));
                    end
                end
            end
          if (((&$signed($unsigned(reg916))) ?
              forvar975 : forvar993[(3'h6):(2'h3)]))
            begin
              for (forvar1037 = (1'h0); (forvar1037 < (2'h2)); forvar1037 = (forvar1037 + (1'h1)))
                begin
                  if (reg917)
                    begin
                      reg1038 <= (!($unsigned($unsigned(forvar946)) ?
                          ($unsigned(reg862) << $signed((8'hba))) : forvar918));
                      reg1039 <= (reg895 ?
                          (reg999[(3'h5):(1'h0)] ?
                              $signed(reg884[(3'h4):(2'h3)]) : ((reg1022 > forvar915) > {reg981})) : reg881[(3'h4):(2'h2)]);
                      reg1040 <= (8'h9d);
                      reg1041 <= $signed($unsigned(reg904));
                    end
                  else
                    begin
                      reg1038 <= ({reg985[(1'h0):(1'h0)]} < ($signed($unsigned((8'had))) << $unsigned(reg918)));
                      reg1039 <= reg956;
                      reg1040 <= ((!{$signed(forvar916)}) ^~ ({(reg845 ?
                                  reg853 : forvar842)} ?
                          ((^~reg924) + $signed(reg899)) : $signed((reg918 <= reg908))));
                    end
                  if ($signed(reg984[(1'h0):(1'h0)]))
                    begin
                      reg1042 <= $unsigned((^($unsigned(reg981) ?
                          $unsigned(reg1015) : (forvar844 ~^ (8'hb7)))));
                    end
                  else
                    begin
                      reg1042 <= {($unsigned({reg928}) ~^ $unsigned((reg943 ?
                              reg938 : reg983)))};
                      reg1043 <= ($signed(((reg943 | reg866) ?
                          reg861[(4'hb):(3'h6)] : (forvar892 && forvar977))) | ({(8'ha7)} ?
                          $signed((reg975 ?
                              reg1025 : reg999)) : $signed($unsigned(forvar938))));
                    end
                  for (forvar1044 = (1'h0); (forvar1044 < (2'h2)); forvar1044 = (forvar1044 + (1'h1)))
                    begin
                      reg1045 <= forvar1002;
                    end
                  for (forvar1046 = (1'h0); (forvar1046 < (2'h3)); forvar1046 = (forvar1046 + (1'h1)))
                    begin
                      reg1047 <= $signed($signed((+(reg1002 > reg920))));
                    end
                end
            end
          else
            begin
              reg1037 <= (reg1009[(3'h7):(3'h4)] < ({(forvar935 >> (8'ha4))} - {$signed(reg980)}));
              for (forvar1038 = (1'h0); (forvar1038 < (2'h2)); forvar1038 = (forvar1038 + (1'h1)))
                begin
                  if ($signed(reg857[(4'h9):(1'h0)]))
                    begin
                      reg1039 <= (8'ha6);
                      reg1040 <= forvar959;
                      reg1041 <= reg993[(4'hb):(4'hb)];
                      reg1042 <= ($unsigned((forvar892[(3'h5):(1'h1)] == reg962)) ?
                          reg930[(1'h0):(1'h0)] : forvar847[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg1039 <= (~^((+$signed(forvar918)) ?
                          (-reg932[(4'h9):(2'h2)]) : $unsigned((^~forvar871))));
                      reg1040 <= ($unsigned({(reg1026 ? reg1042 : reg886)}) ?
                          (~^forvar1010[(1'h1):(1'h1)]) : ((reg1027[(2'h3):(2'h3)] ?
                              (|forvar1010) : reg843[(4'hb):(4'hb)]) <= {{reg856}}));
                    end
                  for (forvar1043 = (1'h0); (forvar1043 < (2'h3)); forvar1043 = (forvar1043 + (1'h1)))
                    begin
                      reg1044 <= (!(({(8'hb6)} | (~|forvar934)) ?
                          $unsigned((reg920 ?
                              reg931 : forvar864)) : forvar901));
                      reg1045 <= (((reg895[(2'h3):(1'h1)] ?
                              {reg904} : forvar971[(2'h3):(1'h1)]) == (forvar925 ?
                              (reg971 > reg859) : (forvar921 >>> reg894))) ?
                          $signed((reg920 ?
                              reg1016[(3'h5):(1'h0)] : (forvar966 ?
                                  forvar876 : (8'ha5)))) : ($signed($unsigned(forvar871)) ?
                              (~&$signed(reg991)) : reg1023[(2'h3):(1'h1)]));
                      reg1046 <= forvar858[(3'h7):(3'h6)];
                      reg1047 <= {{$unsigned((~forvar924))}};
                    end
                  reg1048 <= $signed($unsigned({(reg928 ?
                          reg984 : forvar933)}));
                  if ($unsigned({$unsigned((reg1038 > forvar851))}))
                    begin
                      reg1049 <= {({(~|(8'hb6))} ~^ $unsigned((reg902 ?
                              forvar900 : forvar1022)))};
                    end
                  else
                    begin
                      reg1049 <= reg883[(2'h2):(1'h1)];
                      reg1050 <= (-forvar888);
                      reg1051 <= $unsigned(reg1004);
                    end
                end
              if (reg964[(2'h3):(1'h1)])
                begin
                  reg1052 <= $signed((~|(forvar924 < $signed(forvar838))));
                  if (($signed((8'ha8)) ^ ((forvar901[(3'h4):(3'h4)] <= $signed(reg907)) ?
                      wire4[(1'h0):(1'h0)] : (wire2 * $signed((8'ha5))))))
                    begin
                      reg1053 <= ($unsigned({$signed((8'hb5))}) ?
                          ((~^(!reg1015)) ?
                              ((reg1017 >>> reg950) ^ ((8'ha2) ?
                                  reg961 : (8'ha2))) : (((8'hb0) ?
                                      reg926 : reg981) ?
                                  reg932 : $unsigned(reg931))) : reg962);
                      reg1054 <= $unsigned(reg973);
                      reg1055 <= (~&forvar907[(1'h1):(1'h1)]);
                      reg1056 <= ($signed((~^$signed(forvar967))) ?
                          reg1004[(1'h0):(1'h0)] : $unsigned(reg931));
                    end
                  else
                    begin
                      reg1053 <= (^~(|(~(reg896 < reg845))));
                      reg1054 <= (forvar900 << (((^~(8'hb9)) ?
                          $signed(reg855) : (forvar1024 ?
                              reg872 : forvar1007)) >= ((reg987 && reg867) ?
                          $signed(forvar999) : forvar900)));
                      reg1055 <= ((~&(!(8'hac))) ?
                          (((reg998 | reg1035) ?
                              (|(8'hb6)) : $signed(reg958)) ^ reg915) : {(!(reg870 & reg889))});
                      reg1056 <= reg996;
                    end
                  for (forvar1057 = (1'h0); (forvar1057 < (2'h2)); forvar1057 = (forvar1057 + (1'h1)))
                    begin
                      reg1058 <= $signed((^$signed($signed(forvar992))));
                      reg1059 <= {(^~$signed((reg1014 | reg909)))};
                      reg1060 <= $signed(reg1023[(4'h9):(2'h3)]);
                      reg1061 <= $unsigned((reg918 >> {reg1038}));
                    end
                end
              else
                begin
                  for (forvar1052 = (1'h0); (forvar1052 < (1'h0)); forvar1052 = (forvar1052 + (1'h1)))
                    begin
                      reg1053 <= forvar871;
                    end
                  if ($signed((8'hac)))
                    begin
                      reg1054 <= (~|{reg1014[(2'h3):(2'h3)]});
                      reg1055 <= (~&$unsigned($unsigned(reg967[(4'h8):(2'h3)])));
                    end
                  else
                    begin
                      reg1054 <= $unsigned(($signed($unsigned((8'hb7))) ?
                          forvar995 : (^~(reg891 & forvar863))));
                    end
                  if (reg1056[(3'h4):(1'h1)])
                    begin
                      reg1056 <= (reg1050[(1'h0):(1'h0)] - ((&reg1003[(2'h3):(2'h2)]) >>> ((reg992 - reg913) ?
                          {reg875} : ((8'had) != forvar1002))));
                      reg1057 <= (~|$unsigned({$unsigned(reg903)}));
                      reg1058 <= ((|(^(~&reg971))) >= $signed({$signed((8'h9d))}));
                      reg1059 <= {reg1039[(3'h7):(1'h1)]};
                    end
                  else
                    begin
                      reg1056 <= reg954;
                      reg1057 <= (((8'hab) != (8'ha3)) ?
                          (+reg1013[(1'h1):(1'h1)]) : ($signed(forvar995) <= $signed(reg1023[(2'h3):(1'h1)])));
                    end
                end
            end
          reg1062 <= forvar887;
        end
      reg1063 <= reg924[(1'h0):(1'h0)];
    end
  assign wire1064 = reg920[(3'h6):(3'h5)];
  assign wire1065 = reg885;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module6  (y, clk, wire7, wire8, wire9, wire10, wire11);
  output wire [(32'h189d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire7;
  input wire signed [(2'h2):(1'h0)] wire8;
  input wire signed [(3'h5):(1'h0)] wire9;
  input wire signed [(4'he):(1'h0)] wire10;
  input wire [(4'hf):(1'h0)] wire11;
  wire [(4'hf):(1'h0)] wire833;
  wire signed [(4'hf):(1'h0)] wire832;
  wire signed [(3'h6):(1'h0)] wire831;
  wire signed [(2'h2):(1'h0)] wire12;
  wire [(4'hb):(1'h0)] wire13;
  wire signed [(4'hb):(1'h0)] wire155;
  wire [(4'h8):(1'h0)] wire156;
  wire [(4'ha):(1'h0)] wire171;
  wire [(4'hc):(1'h0)] wire173;
  wire [(4'hd):(1'h0)] wire174;
  wire [(4'h8):(1'h0)] wire447;
  wire signed [(2'h2):(1'h0)] wire609;
  wire [(4'h8):(1'h0)] wire610;
  wire signed [(4'hb):(1'h0)] wire829;
  reg signed [(3'h4):(1'h0)] reg608 = (1'h0);
  reg [(3'h5):(1'h0)] reg606 = (1'h0);
  reg [(2'h2):(1'h0)] reg605 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg603 = (1'h0);
  reg [(3'h5):(1'h0)] reg602 = (1'h0);
  reg [(4'hc):(1'h0)] reg600 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg599 = (1'h0);
  reg [(2'h2):(1'h0)] reg598 = (1'h0);
  reg [(4'h9):(1'h0)] reg586 = (1'h0);
  reg [(4'hb):(1'h0)] reg596 = (1'h0);
  reg [(2'h2):(1'h0)] reg595 = (1'h0);
  reg [(4'hc):(1'h0)] reg594 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg593 = (1'h0);
  reg [(3'h4):(1'h0)] reg592 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg591 = (1'h0);
  reg [(5'h10):(1'h0)] reg590 = (1'h0);
  reg signed [(4'he):(1'h0)] reg589 = (1'h0);
  reg [(3'h5):(1'h0)] reg588 = (1'h0);
  reg [(3'h7):(1'h0)] reg587 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg583 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg582 = (1'h0);
  reg [(4'hd):(1'h0)] reg581 = (1'h0);
  reg [(3'h6):(1'h0)] reg580 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg577 = (1'h0);
  reg [(3'h7):(1'h0)] reg579 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg578 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg576 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg575 = (1'h0);
  reg signed [(4'he):(1'h0)] reg574 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg573 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg572 = (1'h0);
  reg [(4'hd):(1'h0)] reg570 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg569 = (1'h0);
  reg signed [(4'he):(1'h0)] reg568 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg567 = (1'h0);
  reg [(4'hd):(1'h0)] reg565 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg564 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg563 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg562 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg561 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg560 = (1'h0);
  reg [(3'h7):(1'h0)] reg559 = (1'h0);
  reg [(3'h5):(1'h0)] reg558 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg557 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg556 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg554 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg552 = (1'h0);
  reg [(4'hc):(1'h0)] reg551 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg550 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg549 = (1'h0);
  reg [(3'h4):(1'h0)] reg547 = (1'h0);
  reg [(4'ha):(1'h0)] reg546 = (1'h0);
  reg [(4'hf):(1'h0)] reg545 = (1'h0);
  reg [(4'hd):(1'h0)] reg544 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg542 = (1'h0);
  reg signed [(4'he):(1'h0)] reg539 = (1'h0);
  reg [(3'h6):(1'h0)] reg528 = (1'h0);
  reg signed [(4'he):(1'h0)] reg538 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg537 = (1'h0);
  reg [(4'hf):(1'h0)] reg535 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg534 = (1'h0);
  reg [(2'h3):(1'h0)] reg533 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg531 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg530 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg529 = (1'h0);
  reg [(2'h2):(1'h0)] reg527 = (1'h0);
  reg [(3'h5):(1'h0)] reg526 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg525 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg524 = (1'h0);
  reg [(4'hb):(1'h0)] reg523 = (1'h0);
  reg [(3'h5):(1'h0)] reg520 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg519 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg517 = (1'h0);
  reg [(4'hd):(1'h0)] reg516 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg515 = (1'h0);
  reg signed [(4'he):(1'h0)] reg514 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg513 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg512 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg511 = (1'h0);
  reg [(2'h3):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg503 = (1'h0);
  reg [(3'h4):(1'h0)] reg508 = (1'h0);
  reg [(4'h8):(1'h0)] reg507 = (1'h0);
  reg signed [(4'he):(1'h0)] reg506 = (1'h0);
  reg [(4'h9):(1'h0)] reg505 = (1'h0);
  reg [(4'hc):(1'h0)] reg504 = (1'h0);
  reg [(4'hd):(1'h0)] reg502 = (1'h0);
  reg [(3'h5):(1'h0)] reg501 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg500 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg499 = (1'h0);
  reg [(2'h3):(1'h0)] reg498 = (1'h0);
  reg [(4'h9):(1'h0)] reg497 = (1'h0);
  reg signed [(4'he):(1'h0)] reg496 = (1'h0);
  reg [(2'h2):(1'h0)] reg495 = (1'h0);
  reg [(3'h7):(1'h0)] reg494 = (1'h0);
  reg [(4'ha):(1'h0)] reg493 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg491 = (1'h0);
  reg [(4'he):(1'h0)] reg481 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg490 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg489 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg488 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg487 = (1'h0);
  reg [(4'hb):(1'h0)] reg486 = (1'h0);
  reg [(4'ha):(1'h0)] reg485 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg484 = (1'h0);
  reg [(3'h6):(1'h0)] reg483 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg482 = (1'h0);
  reg [(4'he):(1'h0)] reg480 = (1'h0);
  reg [(2'h3):(1'h0)] reg479 = (1'h0);
  reg [(2'h2):(1'h0)] reg478 = (1'h0);
  reg [(4'h8):(1'h0)] reg477 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg473 = (1'h0);
  reg [(4'hf):(1'h0)] reg472 = (1'h0);
  reg [(2'h3):(1'h0)] reg470 = (1'h0);
  reg [(3'h4):(1'h0)] reg471 = (1'h0);
  reg [(4'he):(1'h0)] reg469 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg468 = (1'h0);
  reg [(4'hc):(1'h0)] reg467 = (1'h0);
  reg [(3'h5):(1'h0)] reg466 = (1'h0);
  reg [(5'h10):(1'h0)] reg465 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg464 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg463 = (1'h0);
  reg [(4'ha):(1'h0)] reg462 = (1'h0);
  reg [(3'h7):(1'h0)] reg461 = (1'h0);
  reg [(2'h2):(1'h0)] reg460 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg459 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg458 = (1'h0);
  reg [(3'h4):(1'h0)] reg457 = (1'h0);
  reg [(4'hf):(1'h0)] reg456 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg455 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg454 = (1'h0);
  reg [(4'hc):(1'h0)] reg453 = (1'h0);
  reg [(3'h6):(1'h0)] reg452 = (1'h0);
  reg [(4'he):(1'h0)] reg451 = (1'h0);
  reg [(4'he):(1'h0)] reg449 = (1'h0);
  reg [(4'hc):(1'h0)] reg450 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg446 = (1'h0);
  reg [(2'h2):(1'h0)] reg445 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg444 = (1'h0);
  reg [(2'h2):(1'h0)] reg442 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg440 = (1'h0);
  reg [(4'h8):(1'h0)] reg439 = (1'h0);
  reg [(5'h10):(1'h0)] reg438 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg437 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg436 = (1'h0);
  reg signed [(4'he):(1'h0)] reg409 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg400 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg395 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg431 = (1'h0);
  reg [(2'h3):(1'h0)] reg430 = (1'h0);
  reg [(4'he):(1'h0)] reg429 = (1'h0);
  reg [(3'h7):(1'h0)] reg428 = (1'h0);
  reg [(4'hb):(1'h0)] reg427 = (1'h0);
  reg [(3'h7):(1'h0)] reg426 = (1'h0);
  reg [(3'h6):(1'h0)] reg425 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg424 = (1'h0);
  reg [(4'hb):(1'h0)] reg423 = (1'h0);
  reg signed [(4'he):(1'h0)] reg422 = (1'h0);
  reg [(4'hd):(1'h0)] reg421 = (1'h0);
  reg [(2'h3):(1'h0)] reg420 = (1'h0);
  reg [(4'hd):(1'h0)] reg419 = (1'h0);
  reg [(4'h9):(1'h0)] reg417 = (1'h0);
  reg [(3'h4):(1'h0)] reg418 = (1'h0);
  reg [(4'h9):(1'h0)] reg416 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg415 = (1'h0);
  reg [(3'h6):(1'h0)] reg414 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg413 = (1'h0);
  reg [(4'hf):(1'h0)] reg412 = (1'h0);
  reg [(4'hc):(1'h0)] reg411 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg410 = (1'h0);
  reg [(3'h4):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg401 = (1'h0);
  reg [(4'he):(1'h0)] reg408 = (1'h0);
  reg signed [(4'he):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg405 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg404 = (1'h0);
  reg signed [(4'he):(1'h0)] reg403 = (1'h0);
  reg [(4'hd):(1'h0)] reg402 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg399 = (1'h0);
  reg [(3'h7):(1'h0)] reg398 = (1'h0);
  reg [(3'h6):(1'h0)] reg397 = (1'h0);
  reg [(3'h4):(1'h0)] reg396 = (1'h0);
  reg signed [(4'he):(1'h0)] reg394 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg393 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg391 = (1'h0);
  reg [(2'h3):(1'h0)] reg392 = (1'h0);
  reg signed [(4'he):(1'h0)] reg341 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg390 = (1'h0);
  reg [(3'h6):(1'h0)] reg389 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg388 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg386 = (1'h0);
  reg [(4'he):(1'h0)] reg385 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg383 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg382 = (1'h0);
  reg [(4'hb):(1'h0)] reg381 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg379 = (1'h0);
  reg [(4'ha):(1'h0)] reg378 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg377 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg367 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg376 = (1'h0);
  reg [(2'h3):(1'h0)] reg375 = (1'h0);
  reg [(4'ha):(1'h0)] reg374 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg373 = (1'h0);
  reg [(3'h5):(1'h0)] reg371 = (1'h0);
  reg [(5'h10):(1'h0)] reg370 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg369 = (1'h0);
  reg [(3'h5):(1'h0)] reg368 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg365 = (1'h0);
  reg [(4'hf):(1'h0)] reg364 = (1'h0);
  reg [(4'hb):(1'h0)] reg362 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg361 = (1'h0);
  reg [(5'h10):(1'h0)] reg360 = (1'h0);
  reg [(2'h2):(1'h0)] reg349 = (1'h0);
  reg [(4'hf):(1'h0)] reg345 = (1'h0);
  reg [(4'h8):(1'h0)] reg342 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg359 = (1'h0);
  reg [(4'hc):(1'h0)] reg358 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg357 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg356 = (1'h0);
  reg [(3'h5):(1'h0)] reg355 = (1'h0);
  reg [(4'hf):(1'h0)] reg354 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg353 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg352 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg351 = (1'h0);
  reg [(3'h5):(1'h0)] reg350 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg348 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg347 = (1'h0);
  reg [(3'h7):(1'h0)] reg346 = (1'h0);
  reg [(2'h2):(1'h0)] reg344 = (1'h0);
  reg [(2'h3):(1'h0)] reg343 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg340 = (1'h0);
  reg [(4'hf):(1'h0)] reg339 = (1'h0);
  reg [(4'he):(1'h0)] reg338 = (1'h0);
  reg [(4'hd):(1'h0)] reg337 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg336 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg335 = (1'h0);
  reg [(3'h7):(1'h0)] reg334 = (1'h0);
  reg signed [(4'he):(1'h0)] reg332 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg333 = (1'h0);
  reg [(3'h5):(1'h0)] reg331 = (1'h0);
  reg [(3'h5):(1'h0)] reg330 = (1'h0);
  reg [(3'h4):(1'h0)] reg329 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg325 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg318 = (1'h0);
  reg [(4'ha):(1'h0)] reg315 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg309 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg328 = (1'h0);
  reg [(5'h10):(1'h0)] reg327 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg326 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg324 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg323 = (1'h0);
  reg [(4'h8):(1'h0)] reg322 = (1'h0);
  reg [(4'hc):(1'h0)] reg321 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg320 = (1'h0);
  reg [(3'h6):(1'h0)] reg319 = (1'h0);
  reg [(4'ha):(1'h0)] reg305 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg317 = (1'h0);
  reg [(4'hf):(1'h0)] reg316 = (1'h0);
  reg [(5'h10):(1'h0)] reg314 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg313 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg312 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg311 = (1'h0);
  reg [(4'hf):(1'h0)] reg310 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg308 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg307 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg306 = (1'h0);
  reg [(4'hc):(1'h0)] reg304 = (1'h0);
  reg [(3'h5):(1'h0)] reg303 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg302 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg301 = (1'h0);
  reg [(3'h5):(1'h0)] reg300 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg299 = (1'h0);
  reg [(4'hf):(1'h0)] reg298 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg297 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg296 = (1'h0);
  reg [(4'hf):(1'h0)] reg294 = (1'h0);
  reg [(4'hb):(1'h0)] reg293 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg292 = (1'h0);
  reg [(3'h4):(1'h0)] reg290 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg288 = (1'h0);
  reg [(2'h3):(1'h0)] reg287 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg285 = (1'h0);
  reg [(4'h9):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg283 = (1'h0);
  reg [(3'h7):(1'h0)] reg281 = (1'h0);
  reg [(3'h7):(1'h0)] reg280 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg279 = (1'h0);
  reg [(2'h2):(1'h0)] reg278 = (1'h0);
  reg [(3'h6):(1'h0)] reg277 = (1'h0);
  reg [(3'h4):(1'h0)] reg276 = (1'h0);
  reg [(4'h8):(1'h0)] reg275 = (1'h0);
  reg [(4'he):(1'h0)] reg273 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg272 = (1'h0);
  reg [(4'hf):(1'h0)] reg271 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg270 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg266 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg227 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg248 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg244 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg243 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg234 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg231 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg226 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg263 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg256 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg249 = (1'h0);
  reg [(4'h9):(1'h0)] reg262 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg261 = (1'h0);
  reg [(4'h9):(1'h0)] reg260 = (1'h0);
  reg [(4'hf):(1'h0)] reg259 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg257 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg255 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg254 = (1'h0);
  reg [(4'ha):(1'h0)] reg253 = (1'h0);
  reg [(3'h4):(1'h0)] reg252 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg251 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg250 = (1'h0);
  reg [(5'h10):(1'h0)] reg247 = (1'h0);
  reg [(4'hf):(1'h0)] reg246 = (1'h0);
  reg [(4'h9):(1'h0)] reg245 = (1'h0);
  reg [(4'he):(1'h0)] reg242 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg241 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg240 = (1'h0);
  reg [(2'h2):(1'h0)] reg239 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg238 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg236 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg235 = (1'h0);
  reg [(4'he):(1'h0)] reg233 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg232 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg230 = (1'h0);
  reg [(3'h6):(1'h0)] reg229 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg228 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg224 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg223 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg222 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg221 = (1'h0);
  reg [(3'h4):(1'h0)] reg220 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg218 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg217 = (1'h0);
  reg [(3'h5):(1'h0)] reg216 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg214 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg213 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg212 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg211 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg210 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg209 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg208 = (1'h0);
  reg [(4'hc):(1'h0)] reg206 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg201 = (1'h0);
  reg [(4'hf):(1'h0)] reg199 = (1'h0);
  reg [(4'ha):(1'h0)] reg198 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg197 = (1'h0);
  reg [(4'h9):(1'h0)] reg195 = (1'h0);
  reg [(3'h4):(1'h0)] reg193 = (1'h0);
  reg [(2'h3):(1'h0)] reg192 = (1'h0);
  reg [(5'h10):(1'h0)] reg191 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg189 = (1'h0);
  reg [(2'h2):(1'h0)] reg188 = (1'h0);
  reg [(3'h7):(1'h0)] reg187 = (1'h0);
  reg [(2'h3):(1'h0)] reg185 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg183 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg182 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg180 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg178 = (1'h0);
  reg [(2'h2):(1'h0)] reg154 = (1'h0);
  reg [(5'h10):(1'h0)] reg153 = (1'h0);
  reg [(3'h4):(1'h0)] reg152 = (1'h0);
  reg [(4'hb):(1'h0)] reg150 = (1'h0);
  reg [(2'h2):(1'h0)] reg151 = (1'h0);
  reg [(2'h3):(1'h0)] reg149 = (1'h0);
  reg [(4'hf):(1'h0)] reg148 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg147 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg146 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg142 = (1'h0);
  reg [(3'h4):(1'h0)] reg138 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg144 = (1'h0);
  reg [(4'hd):(1'h0)] reg143 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg141 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg140 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg139 = (1'h0);
  reg [(4'h9):(1'h0)] reg137 = (1'h0);
  reg [(2'h2):(1'h0)] reg136 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg135 = (1'h0);
  reg [(4'ha):(1'h0)] reg134 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg133 = (1'h0);
  reg [(4'he):(1'h0)] reg130 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg129 = (1'h0);
  reg [(4'hf):(1'h0)] reg125 = (1'h0);
  reg [(4'h9):(1'h0)] reg124 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg123 = (1'h0);
  reg [(4'h8):(1'h0)] reg122 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg120 = (1'h0);
  reg [(4'hf):(1'h0)] reg119 = (1'h0);
  reg [(4'hc):(1'h0)] reg118 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg112 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg116 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg115 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg114 = (1'h0);
  reg [(4'he):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg111 = (1'h0);
  reg [(3'h5):(1'h0)] reg110 = (1'h0);
  reg [(4'hf):(1'h0)] reg109 = (1'h0);
  reg [(4'hb):(1'h0)] reg108 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg106 = (1'h0);
  reg [(4'he):(1'h0)] reg105 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg104 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg103 = (1'h0);
  reg [(4'hd):(1'h0)] reg102 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg101 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg100 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg99 = (1'h0);
  reg signed [(4'he):(1'h0)] reg98 = (1'h0);
  reg signed [(4'he):(1'h0)] reg97 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg95 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg94 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg93 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg91 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg88 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg87 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg86 = (1'h0);
  reg [(5'h10):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg84 = (1'h0);
  reg [(2'h3):(1'h0)] reg83 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg82 = (1'h0);
  reg [(4'hc):(1'h0)] reg81 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg80 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg78 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg77 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg75 = (1'h0);
  reg [(4'hc):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg73 = (1'h0);
  reg [(4'he):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg71 = (1'h0);
  reg [(2'h3):(1'h0)] reg70 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg65 = (1'h0);
  reg [(3'h7):(1'h0)] reg64 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg63 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg62 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg61 = (1'h0);
  reg [(2'h2):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg56 = (1'h0);
  reg [(4'ha):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg54 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg53 = (1'h0);
  reg [(4'hb):(1'h0)] reg52 = (1'h0);
  reg [(2'h2):(1'h0)] reg50 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg49 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg45 = (1'h0);
  reg [(4'hd):(1'h0)] reg43 = (1'h0);
  reg [(3'h4):(1'h0)] reg40 = (1'h0);
  reg [(3'h6):(1'h0)] reg36 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg48 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg47 = (1'h0);
  reg [(3'h4):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg44 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg42 = (1'h0);
  reg [(2'h3):(1'h0)] reg41 = (1'h0);
  reg [(2'h3):(1'h0)] reg39 = (1'h0);
  reg [(3'h7):(1'h0)] reg38 = (1'h0);
  reg [(4'hd):(1'h0)] reg37 = (1'h0);
  reg [(4'hf):(1'h0)] reg32 = (1'h0);
  reg [(4'h8):(1'h0)] reg35 = (1'h0);
  reg [(4'hc):(1'h0)] reg34 = (1'h0);
  reg [(3'h6):(1'h0)] reg33 = (1'h0);
  reg [(4'h8):(1'h0)] reg31 = (1'h0);
  reg [(4'hd):(1'h0)] reg30 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg29 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg28 = (1'h0);
  reg [(3'h5):(1'h0)] reg27 = (1'h0);
  reg [(4'ha):(1'h0)] reg15 = (1'h0);
  reg [(4'hc):(1'h0)] reg25 = (1'h0);
  reg [(2'h2):(1'h0)] reg24 = (1'h0);
  reg [(3'h5):(1'h0)] reg23 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg22 = (1'h0);
  reg [(3'h4):(1'h0)] reg21 = (1'h0);
  reg [(4'hc):(1'h0)] reg20 = (1'h0);
  reg [(3'h5):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg18 = (1'h0);
  reg [(3'h5):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg16 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar607 = (1'h0);
  reg [(4'h8):(1'h0)] forvar601 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar597 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar590 = (1'h0);
  reg [(4'h8):(1'h0)] forvar586 = (1'h0);
  reg [(4'hb):(1'h0)] forvar585 = (1'h0);
  reg [(3'h4):(1'h0)] forvar584 = (1'h0);
  reg [(4'hb):(1'h0)] forvar579 = (1'h0);
  reg [(3'h4):(1'h0)] forvar577 = (1'h0);
  reg [(3'h7):(1'h0)] forvar571 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar566 = (1'h0);
  reg [(4'hf):(1'h0)] forvar555 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar553 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar548 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar543 = (1'h0);
  reg [(4'h8):(1'h0)] forvar541 = (1'h0);
  reg [(4'hd):(1'h0)] forvar540 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar526 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar536 = (1'h0);
  reg [(3'h6):(1'h0)] forvar532 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar528 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar522 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar521 = (1'h0);
  reg [(4'h8):(1'h0)] forvar518 = (1'h0);
  reg [(3'h5):(1'h0)] forvar509 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar500 = (1'h0);
  reg [(3'h6):(1'h0)] forvar503 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar493 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar492 = (1'h0);
  reg [(5'h10):(1'h0)] forvar481 = (1'h0);
  reg [(3'h6):(1'h0)] forvar478 = (1'h0);
  reg [(5'h10):(1'h0)] forvar476 = (1'h0);
  reg [(2'h3):(1'h0)] forvar475 = (1'h0);
  reg [(3'h4):(1'h0)] forvar474 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar470 = (1'h0);
  reg [(4'hb):(1'h0)] forvar463 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar452 = (1'h0);
  reg [(3'h5):(1'h0)] forvar449 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar448 = (1'h0);
  reg [(4'h9):(1'h0)] forvar443 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar441 = (1'h0);
  reg [(2'h3):(1'h0)] forvar435 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar434 = (1'h0);
  reg [(4'h9):(1'h0)] forvar433 = (1'h0);
  reg [(4'hd):(1'h0)] forvar432 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar415 = (1'h0);
  reg [(3'h4):(1'h0)] forvar413 = (1'h0);
  reg [(4'he):(1'h0)] forvar410 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar407 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar394 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar397 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar393 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar424 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar428 = (1'h0);
  reg [(4'hc):(1'h0)] forvar422 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar418 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar417 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar409 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar402 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar406 = (1'h0);
  reg [(4'hb):(1'h0)] forvar401 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar400 = (1'h0);
  reg [(4'hf):(1'h0)] forvar395 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar391 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar339 = (1'h0);
  reg [(4'ha):(1'h0)] forvar338 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar335 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar330 = (1'h0);
  reg [(4'hb):(1'h0)] forvar321 = (1'h0);
  reg [(4'hc):(1'h0)] forvar311 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar307 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar308 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar387 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar384 = (1'h0);
  reg [(4'h8):(1'h0)] forvar380 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar368 = (1'h0);
  reg [(4'hc):(1'h0)] forvar372 = (1'h0);
  reg [(4'he):(1'h0)] forvar367 = (1'h0);
  reg [(4'hb):(1'h0)] forvar366 = (1'h0);
  reg [(4'hc):(1'h0)] forvar363 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar358 = (1'h0);
  reg [(4'h8):(1'h0)] forvar353 = (1'h0);
  reg [(3'h5):(1'h0)] forvar349 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar345 = (1'h0);
  reg [(3'h7):(1'h0)] forvar342 = (1'h0);
  reg [(4'h9):(1'h0)] forvar341 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar332 = (1'h0);
  reg [(3'h7):(1'h0)] forvar324 = (1'h0);
  reg [(3'h4):(1'h0)] forvar319 = (1'h0);
  reg [(4'hb):(1'h0)] forvar317 = (1'h0);
  reg [(3'h4):(1'h0)] forvar313 = (1'h0);
  reg [(4'hc):(1'h0)] forvar304 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar325 = (1'h0);
  reg [(4'ha):(1'h0)] forvar318 = (1'h0);
  reg [(3'h5):(1'h0)] forvar315 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar309 = (1'h0);
  reg [(3'h7):(1'h0)] forvar305 = (1'h0);
  reg [(4'h9):(1'h0)] forvar295 = (1'h0);
  reg [(5'h10):(1'h0)] forvar291 = (1'h0);
  reg [(4'he):(1'h0)] forvar286 = (1'h0);
  reg [(2'h2):(1'h0)] forvar282 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar274 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar269 = (1'h0);
  reg [(2'h3):(1'h0)] forvar268 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar267 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar265 = (1'h0);
  reg [(4'h9):(1'h0)] forvar261 = (1'h0);
  reg [(4'he):(1'h0)] forvar253 = (1'h0);
  reg [(5'h10):(1'h0)] forvar239 = (1'h0);
  reg [(3'h5):(1'h0)] forvar233 = (1'h0);
  reg [(4'h9):(1'h0)] forvar228 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar245 = (1'h0);
  reg [(4'hf):(1'h0)] forvar242 = (1'h0);
  reg [(4'hd):(1'h0)] forvar241 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar232 = (1'h0);
  reg [(2'h2):(1'h0)] forvar262 = (1'h0);
  reg [(4'hb):(1'h0)] forvar260 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar258 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar255 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar254 = (1'h0);
  reg [(4'ha):(1'h0)] forvar250 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar256 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar249 = (1'h0);
  reg [(4'hd):(1'h0)] forvar248 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar244 = (1'h0);
  reg [(4'hb):(1'h0)] forvar243 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar237 = (1'h0);
  reg [(2'h3):(1'h0)] forvar234 = (1'h0);
  reg [(3'h5):(1'h0)] forvar231 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar227 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar226 = (1'h0);
  reg [(4'hf):(1'h0)] forvar225 = (1'h0);
  reg [(4'hb):(1'h0)] forvar219 = (1'h0);
  reg [(3'h5):(1'h0)] forvar215 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar207 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar205 = (1'h0);
  reg [(4'hd):(1'h0)] forvar204 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar202 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar200 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar196 = (1'h0);
  reg [(4'hc):(1'h0)] forvar194 = (1'h0);
  reg [(4'hd):(1'h0)] forvar190 = (1'h0);
  reg [(5'h10):(1'h0)] forvar186 = (1'h0);
  reg [(4'he):(1'h0)] forvar184 = (1'h0);
  reg [(2'h3):(1'h0)] forvar181 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar179 = (1'h0);
  reg [(4'he):(1'h0)] forvar177 = (1'h0);
  reg [(3'h7):(1'h0)] forvar176 = (1'h0);
  reg [(4'h9):(1'h0)] forvar175 = (1'h0);
  reg [(4'hf):(1'h0)] forvar149 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar150 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar143 = (1'h0);
  reg [(4'hd):(1'h0)] forvar141 = (1'h0);
  reg [(2'h2):(1'h0)] forvar139 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar135 = (1'h0);
  reg [(4'h9):(1'h0)] forvar142 = (1'h0);
  reg [(4'hb):(1'h0)] forvar138 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar132 = (1'h0);
  reg [(4'h8):(1'h0)] forvar131 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar128 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar127 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar126 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar121 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar118 = (1'h0);
  reg [(4'hf):(1'h0)] forvar113 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar108 = (1'h0);
  reg [(4'hf):(1'h0)] forvar112 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar109 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar107 = (1'h0);
  reg [(4'he):(1'h0)] forvar96 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar90 = (1'h0);
  reg [(4'ha):(1'h0)] forvar89 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar81 = (1'h0);
  reg [(2'h2):(1'h0)] forvar79 = (1'h0);
  reg [(3'h5):(1'h0)] forvar76 = (1'h0);
  reg [(4'he):(1'h0)] forvar71 = (1'h0);
  reg [(4'hb):(1'h0)] forvar68 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar67 = (1'h0);
  reg [(3'h4):(1'h0)] forvar66 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar60 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar58 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar51 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar46 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar41 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar39 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar45 = (1'h0);
  reg [(4'h8):(1'h0)] forvar43 = (1'h0);
  reg [(3'h5):(1'h0)] forvar40 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar36 = (1'h0);
  reg [(4'h9):(1'h0)] forvar32 = (1'h0);
  reg [(2'h2):(1'h0)] forvar26 = (1'h0);
  reg [(2'h2):(1'h0)] forvar21 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar19 = (1'h0);
  reg [(4'h9):(1'h0)] forvar18 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar15 = (1'h0);
  reg [(2'h2):(1'h0)] forvar14 = (1'h0);
  assign y = {wire833,
                 wire832,
                 wire831,
                 wire12,
                 wire13,
                 wire155,
                 wire156,
                 wire171,
                 wire173,
                 wire174,
                 wire447,
                 wire609,
                 wire610,
                 wire829,
                 reg608,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg600,
                 reg599,
                 reg598,
                 reg586,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 reg577,
                 reg579,
                 reg578,
                 reg576,
                 reg575,
                 reg574,
                 reg573,
                 reg572,
                 reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg565,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 reg556,
                 reg554,
                 reg552,
                 reg551,
                 reg550,
                 reg549,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 reg542,
                 reg539,
                 reg528,
                 reg538,
                 reg537,
                 reg535,
                 reg534,
                 reg533,
                 reg531,
                 reg530,
                 reg529,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg520,
                 reg519,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg503,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg502,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg491,
                 reg481,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg480,
                 reg479,
                 reg478,
                 reg477,
                 reg473,
                 reg472,
                 reg470,
                 reg471,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg449,
                 reg450,
                 reg446,
                 reg445,
                 reg444,
                 reg442,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg409,
                 reg400,
                 reg395,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg417,
                 reg418,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 reg406,
                 reg401,
                 reg408,
                 reg407,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg394,
                 reg393,
                 reg391,
                 reg392,
                 reg341,
                 reg390,
                 reg389,
                 reg388,
                 reg386,
                 reg385,
                 reg383,
                 reg382,
                 reg381,
                 reg379,
                 reg378,
                 reg377,
                 reg367,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg365,
                 reg364,
                 reg362,
                 reg361,
                 reg360,
                 reg349,
                 reg345,
                 reg342,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg350,
                 reg348,
                 reg347,
                 reg346,
                 reg344,
                 reg343,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg332,
                 reg333,
                 reg331,
                 reg330,
                 reg329,
                 reg325,
                 reg318,
                 reg315,
                 reg309,
                 reg328,
                 reg327,
                 reg326,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 reg305,
                 reg317,
                 reg316,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg308,
                 reg307,
                 reg306,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg294,
                 reg293,
                 reg292,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg285,
                 reg284,
                 reg283,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg266,
                 reg227,
                 reg248,
                 reg244,
                 reg243,
                 reg234,
                 reg231,
                 reg226,
                 reg264,
                 reg263,
                 reg256,
                 reg249,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg247,
                 reg246,
                 reg245,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg236,
                 reg235,
                 reg233,
                 reg232,
                 reg230,
                 reg229,
                 reg228,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg218,
                 reg217,
                 reg216,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg206,
                 reg203,
                 reg201,
                 reg199,
                 reg198,
                 reg197,
                 reg195,
                 reg193,
                 reg192,
                 reg191,
                 reg189,
                 reg188,
                 reg187,
                 reg185,
                 reg183,
                 reg182,
                 reg180,
                 reg178,
                 reg154,
                 reg153,
                 reg152,
                 reg150,
                 reg151,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg142,
                 reg138,
                 reg145,
                 reg144,
                 reg143,
                 reg141,
                 reg140,
                 reg139,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg130,
                 reg129,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg112,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg78,
                 reg77,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg59,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg50,
                 reg49,
                 reg45,
                 reg43,
                 reg40,
                 reg36,
                 reg48,
                 reg47,
                 reg46,
                 reg44,
                 reg42,
                 reg41,
                 reg39,
                 reg38,
                 reg37,
                 reg32,
                 reg35,
                 reg34,
                 reg33,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg15,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 forvar607,
                 forvar601,
                 forvar597,
                 forvar590,
                 forvar586,
                 forvar585,
                 forvar584,
                 forvar579,
                 forvar577,
                 forvar571,
                 forvar566,
                 forvar555,
                 forvar553,
                 forvar548,
                 forvar543,
                 forvar541,
                 forvar540,
                 forvar526,
                 forvar536,
                 forvar532,
                 forvar528,
                 forvar522,
                 forvar521,
                 forvar518,
                 forvar509,
                 forvar500,
                 forvar503,
                 forvar493,
                 forvar492,
                 forvar481,
                 forvar478,
                 forvar476,
                 forvar475,
                 forvar474,
                 forvar470,
                 forvar463,
                 forvar452,
                 forvar449,
                 forvar448,
                 forvar443,
                 forvar441,
                 forvar435,
                 forvar434,
                 forvar433,
                 forvar432,
                 forvar415,
                 forvar413,
                 forvar410,
                 forvar407,
                 forvar394,
                 forvar397,
                 forvar393,
                 forvar424,
                 forvar428,
                 forvar422,
                 forvar418,
                 forvar417,
                 forvar409,
                 forvar402,
                 forvar406,
                 forvar401,
                 forvar400,
                 forvar395,
                 forvar391,
                 forvar339,
                 forvar338,
                 forvar335,
                 forvar330,
                 forvar321,
                 forvar311,
                 forvar307,
                 forvar308,
                 forvar387,
                 forvar384,
                 forvar380,
                 forvar368,
                 forvar372,
                 forvar367,
                 forvar366,
                 forvar363,
                 forvar358,
                 forvar353,
                 forvar349,
                 forvar345,
                 forvar342,
                 forvar341,
                 forvar332,
                 forvar324,
                 forvar319,
                 forvar317,
                 forvar313,
                 forvar304,
                 forvar325,
                 forvar318,
                 forvar315,
                 forvar309,
                 forvar305,
                 forvar295,
                 forvar291,
                 forvar286,
                 forvar282,
                 forvar274,
                 forvar269,
                 forvar268,
                 forvar267,
                 forvar265,
                 forvar261,
                 forvar253,
                 forvar239,
                 forvar233,
                 forvar228,
                 forvar245,
                 forvar242,
                 forvar241,
                 forvar232,
                 forvar262,
                 forvar260,
                 forvar258,
                 forvar255,
                 forvar254,
                 forvar250,
                 forvar256,
                 forvar249,
                 forvar248,
                 forvar244,
                 forvar243,
                 forvar237,
                 forvar234,
                 forvar231,
                 forvar227,
                 forvar226,
                 forvar225,
                 forvar219,
                 forvar215,
                 forvar207,
                 forvar205,
                 forvar204,
                 forvar202,
                 forvar200,
                 forvar196,
                 forvar194,
                 forvar190,
                 forvar186,
                 forvar184,
                 forvar181,
                 forvar179,
                 forvar177,
                 forvar176,
                 forvar175,
                 forvar149,
                 forvar150,
                 forvar143,
                 forvar141,
                 forvar139,
                 forvar135,
                 forvar142,
                 forvar138,
                 forvar132,
                 forvar131,
                 forvar128,
                 forvar127,
                 forvar126,
                 forvar121,
                 forvar118,
                 forvar113,
                 forvar108,
                 forvar112,
                 forvar109,
                 forvar107,
                 forvar96,
                 forvar90,
                 forvar89,
                 forvar81,
                 forvar79,
                 forvar76,
                 forvar71,
                 forvar68,
                 forvar67,
                 forvar66,
                 forvar60,
                 forvar58,
                 forvar51,
                 forvar46,
                 forvar41,
                 forvar39,
                 forvar45,
                 forvar43,
                 forvar40,
                 forvar36,
                 forvar32,
                 forvar26,
                 forvar21,
                 forvar19,
                 forvar18,
                 forvar15,
                 forvar14,
                 (1'h0)};
  assign wire12 = (8'ha3);
  assign wire13 = (wire8 >= wire8[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      if (wire13)
        begin
          if ($signed(($signed(wire9) ?
              $signed($unsigned(wire12)) : wire12[(1'h1):(1'h0)])))
            begin
              for (forvar14 = (1'h0); (forvar14 < (1'h0)); forvar14 = (forvar14 + (1'h1)))
                begin
                  for (forvar15 = (1'h0); (forvar15 < (1'h1)); forvar15 = (forvar15 + (1'h1)))
                    begin
                      reg16 <= wire8[(1'h0):(1'h0)];
                      reg17 <= $signed((^~((wire10 ? wire10 : (8'hb4)) ?
                          wire8[(1'h1):(1'h1)] : wire11[(2'h2):(1'h1)])));
                      reg18 <= wire8[(1'h1):(1'h0)];
                      reg19 <= ($signed((8'h9d)) ?
                          forvar15 : (-{reg17[(1'h0):(1'h0)]}));
                    end
                  if ($signed((wire13[(4'hb):(2'h2)] ? reg17 : wire7)))
                    begin
                      reg20 <= (wire12 ?
                          {$signed(forvar15[(2'h2):(1'h0)])} : reg17);
                      reg21 <= $unsigned($signed(((wire11 ?
                          reg18 : reg20) ~^ $signed(forvar14))));
                      reg22 <= wire9;
                    end
                  else
                    begin
                      reg20 <= $signed(({wire13[(3'h6):(3'h5)]} ?
                          $unsigned(reg22[(3'h6):(2'h2)]) : (wire11 ?
                              (-wire12) : (wire8 >= wire13))));
                      reg21 <= wire7;
                    end
                  if ($unsigned(((^~(wire13 >> wire10)) >>> $signed((forvar14 ^~ (8'ha9))))))
                    begin
                      reg23 <= $unsigned($signed((wire13 ?
                          $signed(wire7) : reg18)));
                      reg24 <= $signed($signed($unsigned(reg18)));
                      reg25 <= (8'haf);
                    end
                  else
                    begin
                      reg23 <= forvar15[(4'hb):(3'h6)];
                      reg24 <= (wire9 ?
                          $signed((reg18 | $signed(wire13))) : $signed((+(-wire8))));
                      reg25 <= $unsigned((((8'hb4) >>> forvar15[(4'h9):(4'h9)]) ?
                          reg17 : $signed((|reg18))));
                    end
                end
            end
          else
            begin
              for (forvar14 = (1'h0); (forvar14 < (1'h1)); forvar14 = (forvar14 + (1'h1)))
                begin
                  reg15 <= ($signed((~|reg20[(1'h0):(1'h0)])) ?
                      $unsigned((8'ha8)) : reg22[(1'h0):(1'h0)]);
                  if (((-wire8[(2'h2):(2'h2)]) ?
                      {reg21} : {$unsigned($signed(wire8))}))
                    begin
                      reg16 <= $signed($unsigned(reg15));
                      reg17 <= (wire11[(4'hb):(2'h3)] ?
                          ($unsigned((&wire8)) ?
                              wire13 : ($unsigned(wire13) ?
                                  wire12 : (reg15 ?
                                      (8'hb7) : (8'h9e)))) : $unsigned((!(reg18 ?
                              (8'hb1) : reg24))));
                    end
                  else
                    begin
                      reg16 <= wire8[(1'h1):(1'h1)];
                    end
                end
              for (forvar18 = (1'h0); (forvar18 < (1'h0)); forvar18 = (forvar18 + (1'h1)))
                begin
                  for (forvar19 = (1'h0); (forvar19 < (1'h1)); forvar19 = (forvar19 + (1'h1)))
                    begin
                      reg20 <= $signed($unsigned((^~(reg20 ?
                          forvar15 : wire8))));
                    end
                  for (forvar21 = (1'h0); (forvar21 < (2'h2)); forvar21 = (forvar21 + (1'h1)))
                    begin
                      reg22 <= (~$signed((8'hb4)));
                      reg23 <= (wire13 ~^ $signed((wire10 ?
                          (~^reg19) : (8'hb2))));
                      reg24 <= $unsigned((+(forvar15[(4'h8):(3'h7)] <= (reg23 < reg16))));
                      reg25 <= {($unsigned(reg17) ?
                              ((reg22 || (8'ha2)) ?
                                  (!(8'ha3)) : (reg23 ?
                                      reg15 : reg24)) : {$unsigned(reg23)})};
                    end
                  for (forvar26 = (1'h0); (forvar26 < (2'h3)); forvar26 = (forvar26 + (1'h1)))
                    begin
                      reg27 <= {reg24[(1'h1):(1'h0)]};
                      reg28 <= {wire10[(4'ha):(3'h6)]};
                      reg29 <= $signed({(|forvar26)});
                      reg30 <= (~&$signed($unsigned(wire13[(4'ha):(3'h7)])));
                    end
                end
              reg31 <= reg17;
            end
          if ($signed(forvar26))
            begin
              if ($signed($unsigned({$signed(reg16)})))
                begin
                  for (forvar32 = (1'h0); (forvar32 < (2'h2)); forvar32 = (forvar32 + (1'h1)))
                    begin
                      reg33 <= forvar14;
                      reg34 <= ((forvar19[(4'h9):(3'h7)] ?
                          reg17[(2'h2):(2'h2)] : (reg31[(2'h3):(2'h3)] ^~ $signed(wire10))) * $unsigned($signed($unsigned(wire9))));
                      reg35 <= $signed((^~$signed($signed(reg15))));
                    end
                end
              else
                begin
                  if ((^~$unsigned($unsigned((reg24 ? (8'hb2) : reg23)))))
                    begin
                      reg32 <= {((|forvar32[(4'h8):(4'h8)]) ?
                              $unsigned((~&forvar18)) : ((reg30 ?
                                  reg19 : (8'had)) == forvar26))};
                      reg33 <= $signed($signed((~|(~|forvar15))));
                    end
                  else
                    begin
                      reg32 <= $signed($unsigned(reg21));
                    end
                end
              for (forvar36 = (1'h0); (forvar36 < (1'h1)); forvar36 = (forvar36 + (1'h1)))
                begin
                  if (forvar26[(2'h2):(1'h1)])
                    begin
                      reg37 <= (~&((~&{reg28}) ?
                          reg15[(4'ha):(3'h7)] : forvar36[(4'hc):(4'h9)]));
                      reg38 <= (+(8'h9f));
                    end
                  else
                    begin
                      reg37 <= (~&((((8'had) ? forvar26 : reg37) != {wire7}) ?
                          (|$unsigned(forvar26)) : {((8'hac) ?
                                  (8'hba) : wire11)}));
                      reg38 <= reg29;
                      reg39 <= {(&reg22[(2'h3):(2'h3)])};
                    end
                  for (forvar40 = (1'h0); (forvar40 < (1'h0)); forvar40 = (forvar40 + (1'h1)))
                    begin
                      reg41 <= wire9[(2'h2):(1'h0)];
                      reg42 <= $unsigned((forvar32[(2'h3):(1'h0)] ?
                          $signed(reg24) : $unsigned(forvar15[(2'h2):(2'h2)])));
                    end
                end
              for (forvar43 = (1'h0); (forvar43 < (2'h2)); forvar43 = (forvar43 + (1'h1)))
                begin
                  reg44 <= $unsigned({$signed(reg23)});
                  for (forvar45 = (1'h0); (forvar45 < (2'h2)); forvar45 = (forvar45 + (1'h1)))
                    begin
                      reg46 <= reg28[(4'h9):(1'h0)];
                      reg47 <= ({((reg41 <<< reg18) > $signed(reg27))} ?
                          $unsigned($unsigned(forvar15[(3'h7):(2'h3)])) : $signed(forvar26[(1'h1):(1'h1)]));
                      reg48 <= (~|$unsigned($unsigned((forvar32 << reg30))));
                    end
                end
            end
          else
            begin
              if ($unsigned($signed($signed((forvar40 + forvar21)))))
                begin
                  if ({$unsigned(reg31)})
                    begin
                      reg32 <= ({((reg35 ? wire13 : wire9) >= $signed(reg39))} ?
                          $signed((forvar40 | $signed(reg34))) : (wire12 ?
                              (&wire11[(3'h5):(1'h1)]) : reg25[(3'h5):(2'h3)]));
                      reg33 <= reg16;
                      reg34 <= $unsigned($signed($signed($signed(wire13))));
                    end
                  else
                    begin
                      reg32 <= $signed((reg21[(2'h3):(2'h3)] ?
                          (&(~&reg33)) : reg24[(2'h2):(1'h0)]));
                      reg33 <= (!($unsigned({reg38}) <<< $signed((reg42 ^~ forvar32))));
                      reg34 <= $signed($unsigned({(forvar26 ?
                              forvar43 : (8'hb1))}));
                      reg35 <= ((($unsigned(wire8) ?
                              forvar45 : (~^reg30)) <= $signed(reg34[(3'h7):(3'h7)])) ?
                          forvar40 : reg41);
                    end
                  if ({({$unsigned((8'ha1))} >>> $signed((reg48 <<< reg32)))})
                    begin
                      reg36 <= $unsigned(({reg18[(1'h0):(1'h0)]} & reg30[(1'h1):(1'h0)]));
                      reg37 <= ((({reg35} & reg28[(3'h4):(3'h4)]) ?
                          $signed((!forvar15)) : (reg35 > reg36[(3'h6):(1'h1)])) >> forvar26[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg36 <= ({(~$unsigned(forvar21))} ?
                          (reg22 == forvar40) : $signed($unsigned(((8'hb0) <= wire8))));
                      reg37 <= (8'h9c);
                    end
                  reg38 <= (~&(~|forvar14[(1'h1):(1'h1)]));
                  for (forvar39 = (1'h0); (forvar39 < (1'h1)); forvar39 = (forvar39 + (1'h1)))
                    begin
                      reg40 <= forvar14[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar32 = (1'h0); (forvar32 < (2'h2)); forvar32 = (forvar32 + (1'h1)))
                    begin
                      reg33 <= ($signed({$signed((8'ha1))}) ?
                          ((forvar14[(1'h0):(1'h0)] >>> reg24[(1'h1):(1'h1)]) ?
                              {$unsigned(reg25)} : (~reg30)) : ((8'hac) ?
                              reg28 : $signed((reg16 ? forvar15 : (8'ha1)))));
                      reg34 <= (reg16 ?
                          ($signed(reg28[(4'h9):(3'h4)]) || {(reg28 ?
                                  wire7 : reg46)}) : ($signed((^reg46)) * $unsigned(reg48[(1'h0):(1'h0)])));
                      reg35 <= (~|(($signed(reg47) >= (^~reg39)) ?
                          (|{reg19}) : $signed($unsigned(reg41))));
                    end
                  if ((^~((~&$unsigned(forvar18)) > reg24)))
                    begin
                      reg36 <= {{$unsigned(forvar39[(4'hd):(1'h0)])}};
                      reg37 <= wire10;
                      reg38 <= ((&((~^(8'h9d)) ?
                              reg21[(3'h4):(1'h0)] : (8'ha0))) ?
                          forvar15 : (+{{forvar26}}));
                      reg39 <= wire10;
                    end
                  else
                    begin
                      reg36 <= {forvar26};
                      reg37 <= reg29[(4'h9):(3'h5)];
                      reg38 <= $unsigned((-$unsigned(reg32[(1'h0):(1'h0)])));
                      reg39 <= $unsigned({$signed($signed(reg22))});
                    end
                  reg40 <= ($unsigned(forvar39) << {$signed($unsigned((8'hae)))});
                  for (forvar41 = (1'h0); (forvar41 < (1'h0)); forvar41 = (forvar41 + (1'h1)))
                    begin
                      reg42 <= (8'h9c);
                      reg43 <= {(^~reg30[(3'h4):(3'h4)])};
                      reg44 <= (reg15 != $unsigned(reg43));
                      reg45 <= reg41;
                    end
                end
              for (forvar46 = (1'h0); (forvar46 < (1'h1)); forvar46 = (forvar46 + (1'h1)))
                begin
                  if (((forvar26 ?
                      $unsigned($unsigned(forvar32)) : ($unsigned(reg44) ?
                          $unsigned(wire8) : (!(8'h9d)))) - (~&{(reg29 ?
                          (8'ha9) : wire13)})))
                    begin
                      reg47 <= (^~((reg47[(3'h6):(3'h5)] >= reg45) - $signed(reg44)));
                      reg48 <= (+$signed(((~forvar45) ?
                          wire7[(1'h0):(1'h0)] : wire11)));
                      reg49 <= reg36;
                      reg50 <= ($signed((forvar32 ^ $unsigned(wire12))) != {(^reg28)});
                    end
                  else
                    begin
                      reg47 <= reg24[(1'h0):(1'h0)];
                      reg48 <= ((~&forvar36[(2'h3):(1'h0)]) ^ reg45);
                    end
                  for (forvar51 = (1'h0); (forvar51 < (1'h1)); forvar51 = (forvar51 + (1'h1)))
                    begin
                      reg52 <= wire12;
                      reg53 <= $signed(($unsigned({reg31}) ^~ ({reg39} && {reg18})));
                    end
                  if ((^~(~|($signed(reg44) - (reg49 ? (8'ha9) : (8'hab))))))
                    begin
                      reg54 <= (~|{forvar39[(4'hf):(2'h3)]});
                    end
                  else
                    begin
                      reg54 <= (~|reg21);
                    end
                  if ((forvar39[(5'h10):(1'h1)] != $unsigned(forvar40[(2'h2):(1'h0)])))
                    begin
                      reg55 <= (|reg36[(3'h5):(2'h3)]);
                      reg56 <= $unsigned($unsigned($signed($unsigned(forvar51))));
                      reg57 <= $signed((8'hae));
                    end
                  else
                    begin
                      reg55 <= $signed((8'h9c));
                    end
                end
              for (forvar58 = (1'h0); (forvar58 < (2'h2)); forvar58 = (forvar58 + (1'h1)))
                begin
                  if ($unsigned({$signed(((8'haa) <<< (8'h9e)))}))
                    begin
                      reg59 <= {(((reg15 & reg28) ?
                                  forvar39[(3'h7):(1'h1)] : reg22[(3'h4):(2'h2)]) ?
                              $unsigned(reg40[(3'h4):(1'h1)]) : (+{reg44}))};
                    end
                  else
                    begin
                      reg59 <= ((((reg37 >= reg37) ? reg28 : $signed(reg49)) ?
                              (&$unsigned(forvar40)) : forvar40) ?
                          reg44[(2'h3):(2'h3)] : (($unsigned((8'hb4)) ?
                              (reg59 ?
                                  reg48 : reg28) : $unsigned(reg23)) << ((reg15 > reg39) * (forvar36 ?
                              (8'ha3) : wire9))));
                    end
                  for (forvar60 = (1'h0); (forvar60 < (1'h1)); forvar60 = (forvar60 + (1'h1)))
                    begin
                      reg61 <= $unsigned($signed(((forvar15 ?
                              reg42 : forvar39) ?
                          (reg41 ? reg44 : (8'hb5)) : $signed(wire7))));
                      reg62 <= (~^{$signed(reg31)});
                      reg63 <= reg44[(3'h4):(2'h3)];
                    end
                  reg64 <= reg17;
                  reg65 <= (reg63 ?
                      $signed($unsigned(reg33)) : $signed(((8'ha1) <= $unsigned(reg45))));
                end
            end
        end
      else
        begin
          for (forvar14 = (1'h0); (forvar14 < (2'h2)); forvar14 = (forvar14 + (1'h1)))
            begin
              reg15 <= (reg59[(1'h0):(1'h0)] < forvar58);
              reg16 <= $signed(($unsigned($unsigned(reg28)) ?
                  ({(8'ha4)} + (8'ha5)) : $unsigned($signed(reg17))));
            end
          reg17 <= (^reg53);
        end
      for (forvar66 = (1'h0); (forvar66 < (2'h2)); forvar66 = (forvar66 + (1'h1)))
        begin
          for (forvar67 = (1'h0); (forvar67 < (2'h2)); forvar67 = (forvar67 + (1'h1)))
            begin
              if (forvar18)
                begin
                  for (forvar68 = (1'h0); (forvar68 < (2'h2)); forvar68 = (forvar68 + (1'h1)))
                    begin
                      reg69 <= ((8'hb8) * $signed($signed($unsigned(reg21))));
                      reg70 <= $unsigned(($unsigned($signed(reg42)) >>> forvar14[(1'h0):(1'h0)]));
                      reg71 <= (reg31 && (~&(reg55[(3'h4):(3'h4)] != $unsigned(reg47))));
                      reg72 <= (-reg33[(1'h1):(1'h0)]);
                    end
                  reg73 <= (forvar15[(4'hc):(3'h4)] <<< (+(-$unsigned(reg49))));
                end
              else
                begin
                  for (forvar68 = (1'h0); (forvar68 < (1'h1)); forvar68 = (forvar68 + (1'h1)))
                    begin
                      reg69 <= (8'haf);
                      reg70 <= {($signed(forvar18[(1'h1):(1'h1)]) ?
                              (reg73 ?
                                  reg36 : (reg20 ?
                                      forvar51 : reg41)) : $unsigned((&(8'ha6))))};
                    end
                  for (forvar71 = (1'h0); (forvar71 < (1'h1)); forvar71 = (forvar71 + (1'h1)))
                    begin
                      reg72 <= reg45;
                      reg73 <= ((((~&reg44) || (reg43 ? reg69 : forvar60)) ?
                          (^~forvar15) : (^$unsigned(forvar36))) != {$unsigned(reg34)});
                      reg74 <= forvar32[(4'h9):(4'h9)];
                      reg75 <= reg22;
                    end
                  for (forvar76 = (1'h0); (forvar76 < (1'h1)); forvar76 = (forvar76 + (1'h1)))
                    begin
                      reg77 <= (reg21 >> ((forvar41 > (reg20 * reg16)) >> (+reg49)));
                      reg78 <= reg55[(2'h3):(1'h0)];
                    end
                  for (forvar79 = (1'h0); (forvar79 < (1'h0)); forvar79 = (forvar79 + (1'h1)))
                    begin
                      reg80 <= (~{(reg69[(2'h2):(1'h1)] >>> (reg15 > forvar18))});
                    end
                end
              if ($signed({{(reg72 || reg52)}}))
                begin
                  if (reg16[(4'he):(1'h1)])
                    begin
                      reg81 <= reg64;
                      reg82 <= (($unsigned(wire7[(1'h1):(1'h0)]) ?
                              reg81 : (^(8'ha6))) ?
                          reg33[(3'h4):(3'h4)] : $signed(($signed(reg71) ?
                              $signed((8'ha0)) : $signed(reg34))));
                      reg83 <= reg33;
                      reg84 <= reg80[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg81 <= $unsigned($unsigned(reg59[(2'h2):(2'h2)]));
                    end
                  if ({({(forvar41 < forvar32)} ?
                          ($unsigned(reg82) < forvar58[(3'h7):(3'h7)]) : $signed((reg69 ?
                              reg83 : forvar26)))})
                    begin
                      reg85 <= $unsigned(((^reg19) ?
                          $unsigned({reg73}) : (+{reg52})));
                      reg86 <= (8'ha4);
                      reg87 <= forvar26;
                      reg88 <= reg44[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg85 <= $unsigned($signed((reg18 ^~ {reg29})));
                    end
                end
              else
                begin
                  for (forvar81 = (1'h0); (forvar81 < (2'h3)); forvar81 = (forvar81 + (1'h1)))
                    begin
                      reg82 <= (forvar51[(4'h8):(3'h6)] < reg33[(1'h1):(1'h1)]);
                    end
                  if ((~|(~(~(&(8'ha9))))))
                    begin
                      reg83 <= (reg50[(1'h1):(1'h1)] <= (8'hb7));
                    end
                  else
                    begin
                      reg83 <= {reg37[(4'hc):(4'hc)]};
                      reg84 <= reg24;
                    end
                end
              for (forvar89 = (1'h0); (forvar89 < (1'h1)); forvar89 = (forvar89 + (1'h1)))
                begin
                  for (forvar90 = (1'h0); (forvar90 < (2'h2)); forvar90 = (forvar90 + (1'h1)))
                    begin
                      reg91 <= $signed($signed((reg17[(2'h3):(1'h0)] - forvar79)));
                      reg92 <= forvar41;
                    end
                  if ($unsigned((8'ha3)))
                    begin
                      reg93 <= reg86[(2'h3):(1'h1)];
                      reg94 <= $signed(($signed((&reg93)) ?
                          $signed((~|reg59)) : {(~^(8'hab))}));
                    end
                  else
                    begin
                      reg93 <= ((^~((^reg18) ?
                              $unsigned(forvar18) : $unsigned(forvar14))) ?
                          (({(8'hb0)} >> (reg19 ? forvar45 : (8'ha7))) ?
                              $signed($signed(reg64)) : {{reg46}}) : $unsigned($signed($unsigned(reg32))));
                      reg94 <= $signed($unsigned({forvar51[(4'h9):(4'h9)]}));
                      reg95 <= (~&{{$unsigned((8'ha1))}});
                    end
                  for (forvar96 = (1'h0); (forvar96 < (1'h0)); forvar96 = (forvar96 + (1'h1)))
                    begin
                      reg97 <= ((^reg40) ?
                          (((reg62 ?
                              reg91 : reg56) >>> reg62[(2'h3):(2'h2)]) <= $signed((!forvar90))) : (~&(|(8'hb6))));
                      reg98 <= ($signed(($unsigned(reg85) ?
                              (~reg61) : (reg78 >= reg25))) ?
                          wire9[(3'h4):(3'h4)] : (!(((8'ha2) > (8'h9c)) ?
                              (forvar51 ?
                                  forvar51 : wire13) : reg71[(3'h5):(2'h2)])));
                      reg99 <= $unsigned($signed({(reg17 ? reg34 : forvar43)}));
                    end
                  if ($unsigned(((((8'h9e) >>> forvar46) ?
                          ((8'hab) ? reg93 : reg80) : (-reg37)) ?
                      ({wire13} - forvar39[(1'h1):(1'h0)]) : $unsigned((reg39 >>> (8'hb9))))))
                    begin
                      reg100 <= reg43[(4'hb):(3'h5)];
                      reg101 <= ((reg87 ?
                              (8'ha2) : $signed($unsigned((8'hb9)))) ?
                          $signed({wire11[(3'h5):(2'h2)]}) : (reg64 - $unsigned((reg82 >> forvar60))));
                      reg102 <= $signed(forvar58[(3'h6):(1'h0)]);
                      reg103 <= ((((reg40 ^~ reg78) << reg34) + $signed($unsigned(reg42))) ?
                          ($signed((~&wire10)) < $unsigned(forvar96)) : wire8);
                    end
                  else
                    begin
                      reg100 <= $signed($unsigned(reg19[(2'h3):(1'h0)]));
                      reg101 <= $signed($unsigned(($signed(reg63) ?
                          reg24[(2'h2):(1'h0)] : (+wire12))));
                      reg102 <= (-(((~&reg31) ? forvar18 : (~|reg41)) ?
                          $unsigned((reg61 ? reg59 : (8'hb2))) : forvar79));
                      reg103 <= reg47;
                    end
                end
              reg104 <= (!reg69[(4'h8):(1'h0)]);
            end
          reg105 <= $signed(reg95[(2'h2):(1'h1)]);
          reg106 <= (+(^~$unsigned($unsigned((8'had)))));
        end
      if ((reg91 <= {(~reg30)}))
        begin
          for (forvar107 = (1'h0); (forvar107 < (2'h2)); forvar107 = (forvar107 + (1'h1)))
            begin
              if (({reg21[(1'h1):(1'h1)]} ?
                  (reg95 ?
                      {(reg48 ? reg75 : reg17)} : ((reg57 ? reg70 : forvar51) ?
                          reg55 : reg15)) : (+{forvar90})))
                begin
                  reg108 <= (((8'h9c) - (((8'hae) ?
                      reg92 : reg23) + $unsigned(reg49))) + (reg35 ?
                      $unsigned(((8'hab) ?
                          reg71 : (8'ha1))) : reg55[(2'h3):(1'h0)]));
                  if (((!$signed((reg78 | reg71))) ?
                      {(~|(reg45 <<< (8'ha3)))} : (reg92 & reg18[(3'h4):(2'h2)])))
                    begin
                      reg109 <= {{(8'ha9)}};
                      reg110 <= ((($unsigned(forvar19) ?
                                  ((8'ha3) >= reg88) : (wire9 ?
                                      (8'hb4) : reg63)) ?
                              $unsigned({(8'hab)}) : $unsigned($unsigned(reg85))) ?
                          $unsigned((reg30[(4'ha):(2'h2)] == reg93[(3'h4):(3'h4)])) : $unsigned(wire8[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg109 <= (8'ha8);
                    end
                end
              else
                begin
                  reg108 <= $unsigned($signed((~^reg85)));
                  for (forvar109 = (1'h0); (forvar109 < (1'h0)); forvar109 = (forvar109 + (1'h1)))
                    begin
                      reg110 <= forvar14;
                      reg111 <= (+$signed({$signed(forvar58)}));
                    end
                end
            end
        end
      else
        begin
          for (forvar107 = (1'h0); (forvar107 < (2'h3)); forvar107 = (forvar107 + (1'h1)))
            begin
              if ((|$signed($signed(((8'ha2) ? reg111 : reg54)))))
                begin
                  if (($signed((reg53[(4'h9):(4'h8)] ?
                      (reg93 >>> reg43) : forvar21)) - $unsigned($unsigned(reg42[(4'hd):(4'hb)]))))
                    begin
                      reg108 <= (~&$unsigned($signed(forvar79[(1'h0):(1'h0)])));
                      reg109 <= $signed($signed((~$unsigned(forvar51))));
                    end
                  else
                    begin
                      reg108 <= (~reg99);
                      reg109 <= (^(({reg29} >> (~reg57)) == $signed(forvar19[(4'ha):(3'h4)])));
                      reg110 <= {forvar60};
                    end
                  reg111 <= $unsigned($unsigned((!((8'ha9) ?
                      reg34 : forvar19))));
                  for (forvar112 = (1'h0); (forvar112 < (2'h3)); forvar112 = (forvar112 + (1'h1)))
                    begin
                      reg113 <= ($signed(((forvar14 ? reg99 : reg80) ?
                          {reg87} : $signed(reg44))) >= {reg54});
                      reg114 <= ((^reg56) <= (reg111[(3'h4):(1'h0)] ?
                          ($signed(forvar39) & reg53[(3'h4):(1'h1)]) : reg42));
                      reg115 <= (^{(8'haa)});
                      reg116 <= (~&$signed((|reg77[(2'h3):(2'h3)])));
                    end
                end
              else
                begin
                  for (forvar108 = (1'h0); (forvar108 < (2'h2)); forvar108 = (forvar108 + (1'h1)))
                    begin
                      reg109 <= ((8'ha0) ?
                          reg46[(2'h2):(1'h1)] : $signed($unsigned($unsigned(reg16))));
                      reg110 <= {reg85};
                      reg111 <= $signed(((!$unsigned(reg81)) ^ $signed(((8'ha0) == reg101))));
                      reg112 <= (|(reg49[(2'h2):(2'h2)] ?
                          ($unsigned(reg55) >> (forvar79 ?
                              reg109 : (8'h9e))) : (^~forvar26)));
                    end
                  for (forvar113 = (1'h0); (forvar113 < (2'h2)); forvar113 = (forvar113 + (1'h1)))
                    begin
                      reg114 <= $signed((($unsigned((8'ha3)) ?
                          $signed(reg78) : (forvar113 ?
                              forvar15 : forvar26)) != (~&reg25[(3'h4):(1'h0)])));
                      reg115 <= reg27;
                      reg116 <= ((!$signed($unsigned(reg72))) ? reg42 : reg23);
                    end
                end
              if (forvar89[(3'h5):(2'h2)])
                begin
                  if (reg69[(3'h4):(2'h3)])
                    begin
                      reg117 <= $unsigned(reg28[(3'h5):(2'h2)]);
                      reg118 <= ({{(reg18 ? (8'h9e) : reg44)}} ?
                          {$unsigned((8'ha3))} : {(8'ha5)});
                    end
                  else
                    begin
                      reg117 <= ($unsigned(wire10) <<< $unsigned(reg42[(1'h0):(1'h0)]));
                      reg118 <= {forvar81[(3'h5):(2'h2)]};
                      reg119 <= $signed($unsigned((-{forvar32})));
                      reg120 <= {(reg94 ?
                              (8'hb5) : $unsigned($signed(forvar36)))};
                    end
                end
              else
                begin
                  reg117 <= $unsigned((~forvar81[(3'h5):(2'h2)]));
                  for (forvar118 = (1'h0); (forvar118 < (1'h0)); forvar118 = (forvar118 + (1'h1)))
                    begin
                      reg119 <= (^~(+reg46[(1'h0):(1'h0)]));
                      reg120 <= (^~($signed(((8'hb1) ? forvar60 : reg91)) ?
                          forvar113 : $signed((reg119 * (8'hab)))));
                    end
                end
              if ((~^$unsigned($signed($signed(reg49)))))
                begin
                  for (forvar121 = (1'h0); (forvar121 < (2'h2)); forvar121 = (forvar121 + (1'h1)))
                    begin
                      reg122 <= reg65[(4'hd):(4'h9)];
                      reg123 <= $unsigned((reg93 ?
                          (~&reg19[(3'h4):(2'h2)]) : ($unsigned((8'ha8)) ?
                              $unsigned(reg41) : (reg47 ? forvar40 : reg112))));
                      reg124 <= reg97;
                      reg125 <= ((((forvar19 >>> forvar58) ?
                                  forvar39 : $signed(reg97)) ?
                              $unsigned($signed(reg43)) : ($unsigned(forvar40) ?
                                  $signed((8'hb4)) : {reg120})) ?
                          forvar51 : $unsigned((~(8'ha7))));
                    end
                end
              else
                begin
                  for (forvar121 = (1'h0); (forvar121 < (1'h0)); forvar121 = (forvar121 + (1'h1)))
                    begin
                      reg122 <= reg77[(2'h2):(1'h0)];
                      reg123 <= $signed(forvar26);
                    end
                end
            end
          for (forvar126 = (1'h0); (forvar126 < (1'h1)); forvar126 = (forvar126 + (1'h1)))
            begin
              for (forvar127 = (1'h0); (forvar127 < (2'h3)); forvar127 = (forvar127 + (1'h1)))
                begin
                  for (forvar128 = (1'h0); (forvar128 < (1'h1)); forvar128 = (forvar128 + (1'h1)))
                    begin
                      reg129 <= (|$signed(($signed(reg115) ?
                          forvar68 : (forvar26 ? (8'hab) : reg125))));
                      reg130 <= {$unsigned(($unsigned(reg97) ?
                              {reg44} : ((8'ha7) ^ reg108)))};
                    end
                end
              for (forvar131 = (1'h0); (forvar131 < (1'h1)); forvar131 = (forvar131 + (1'h1)))
                begin
                  for (forvar132 = (1'h0); (forvar132 < (2'h2)); forvar132 = (forvar132 + (1'h1)))
                    begin
                      reg133 <= $unsigned(reg54);
                      reg134 <= $unsigned($signed(($unsigned(reg46) ?
                          (reg39 ? (8'h9c) : reg28) : wire10[(4'hd):(3'h6)])));
                    end
                end
            end
          if (forvar71[(4'hc):(3'h7)])
            begin
              if ((($signed($unsigned((8'hb3))) ?
                  $signed((^~reg78)) : reg106[(1'h0):(1'h0)]) << $signed(forvar19)))
                begin
                  if ((reg32 ?
                      forvar14 : $unsigned((reg81[(4'hb):(3'h5)] ?
                          (forvar58 ^ reg81) : (reg87 ? reg65 : reg31)))))
                    begin
                      reg135 <= (forvar76 != {((reg38 + (8'ha8)) ?
                              (reg61 || reg32) : {forvar107})});
                    end
                  else
                    begin
                      reg135 <= $unsigned(forvar81);
                      reg136 <= $unsigned($signed($unsigned((reg64 ?
                          reg21 : reg23))));
                      reg137 <= $signed($signed((reg87[(2'h2):(2'h2)] > (forvar43 ?
                          wire7 : forvar58))));
                    end
                  for (forvar138 = (1'h0); (forvar138 < (2'h2)); forvar138 = (forvar138 + (1'h1)))
                    begin
                      reg139 <= ($signed(($unsigned(reg22) ?
                              (8'ha3) : $signed(wire13))) ?
                          ($signed({reg102}) ?
                              $signed($unsigned(reg118)) : reg62) : forvar46[(3'h6):(3'h4)]);
                      reg140 <= {$signed((+reg35[(4'h8):(1'h1)]))};
                      reg141 <= ((-((forvar127 ? reg99 : reg87) ?
                          reg28[(4'h9):(1'h1)] : $signed(reg122))) - ((~|reg87) >>> (+$unsigned(reg65))));
                    end
                  for (forvar142 = (1'h0); (forvar142 < (2'h2)); forvar142 = (forvar142 + (1'h1)))
                    begin
                      reg143 <= ({$signed(forvar46[(4'h8):(3'h5)])} ?
                          (-((|reg92) ?
                              (reg64 ?
                                  reg52 : forvar58) : (~|(8'h9c)))) : {$signed((+forvar112))});
                      reg144 <= (|forvar108[(2'h2):(1'h0)]);
                      reg145 <= (reg33[(1'h1):(1'h1)] ?
                          (reg122[(3'h6):(1'h1)] >>> $unsigned($unsigned((8'hba)))) : $signed(((reg111 ~^ reg101) ?
                              reg124[(2'h3):(1'h1)] : (reg125 >>> reg63))));
                    end
                end
              else
                begin
                  for (forvar135 = (1'h0); (forvar135 < (1'h0)); forvar135 = (forvar135 + (1'h1)))
                    begin
                      reg136 <= $signed((~&((forvar107 != forvar71) ?
                          forvar40[(3'h4):(3'h4)] : $signed(reg139))));
                      reg137 <= (~|(($unsigned(reg44) ?
                          (forvar108 ?
                              reg100 : reg72) : $unsigned(reg50)) ^ reg70[(1'h0):(1'h0)]));
                      reg138 <= (reg35[(3'h5):(2'h2)] * $signed(reg112[(1'h1):(1'h0)]));
                    end
                  for (forvar139 = (1'h0); (forvar139 < (2'h2)); forvar139 = (forvar139 + (1'h1)))
                    begin
                      reg140 <= reg46;
                    end
                  for (forvar141 = (1'h0); (forvar141 < (2'h3)); forvar141 = (forvar141 + (1'h1)))
                    begin
                      reg142 <= $unsigned((((reg74 ?
                              reg21 : reg103) >= ((8'ha3) >> reg37)) ?
                          ((forvar39 ? reg135 : forvar71) ?
                              forvar39[(3'h7):(3'h4)] : reg30) : ({reg73} - forvar128)));
                    end
                  for (forvar143 = (1'h0); (forvar143 < (1'h0)); forvar143 = (forvar143 + (1'h1)))
                    begin
                      reg144 <= (reg124 ?
                          $signed((forvar18[(4'h9):(4'h9)] - reg73[(3'h4):(1'h0)])) : reg55);
                      reg145 <= reg105;
                      reg146 <= $unsigned((((reg39 ? reg28 : reg118) ?
                          (forvar46 ?
                              reg140 : reg73) : reg45[(2'h3):(1'h0)]) ^ ({reg46} ^ $unsigned((8'hba)))));
                      reg147 <= $unsigned({(8'ha1)});
                    end
                end
              if ($signed(reg87[(1'h0):(1'h0)]))
                begin
                  if ((reg137[(1'h1):(1'h0)] ~^ forvar14))
                    begin
                      reg148 <= reg45;
                      reg149 <= (+(reg38 ?
                          {(reg34 ?
                                  (8'ha0) : reg97)} : $unsigned($unsigned(reg147))));
                    end
                  else
                    begin
                      reg148 <= $signed($unsigned(reg141[(3'h4):(2'h3)]));
                    end
                  for (forvar150 = (1'h0); (forvar150 < (1'h0)); forvar150 = (forvar150 + (1'h1)))
                    begin
                      reg151 <= {{(forvar18[(1'h1):(1'h0)] ?
                                  reg55 : (reg35 <<< reg28))}};
                    end
                end
              else
                begin
                  reg148 <= {($unsigned($unsigned(forvar138)) >>> reg103[(1'h1):(1'h1)])};
                  for (forvar149 = (1'h0); (forvar149 < (2'h2)); forvar149 = (forvar149 + (1'h1)))
                    begin
                      reg150 <= $signed(reg40[(1'h0):(1'h0)]);
                      reg151 <= {$signed((reg44[(1'h1):(1'h0)] ?
                              reg18[(1'h1):(1'h1)] : (^reg137)))};
                      reg152 <= reg122[(4'h8):(1'h0)];
                      reg153 <= $signed((((+forvar18) ?
                          (8'hba) : $signed(reg77)) < $signed($signed(reg15))));
                    end
                end
            end
          else
            begin
              if ({reg63[(2'h3):(2'h3)]})
                begin
                  reg135 <= (~&(^~reg130[(3'h4):(1'h1)]));
                  reg136 <= ($unsigned(reg17[(1'h1):(1'h0)]) && (^$signed(forvar118)));
                  reg137 <= reg130;
                end
              else
                begin
                  if ((^$unsigned((&(reg29 ? forvar127 : reg50)))))
                    begin
                      reg135 <= (reg18 ?
                          $unsigned(reg29[(4'h8):(3'h6)]) : $signed($signed((reg57 ?
                              reg83 : reg98))));
                      reg136 <= $unsigned((&$signed({reg15})));
                      reg137 <= reg52;
                      reg138 <= (~^(8'hb1));
                    end
                  else
                    begin
                      reg135 <= $signed(reg152);
                    end
                end
            end
          reg154 <= ({reg21[(2'h2):(1'h1)]} ? wire11[(2'h3):(2'h3)] : forvar90);
        end
    end
  assign wire155 = (&reg85);
  assign wire156 = (~|$unsigned($signed(reg97)));
  module157 #() modinst172 (wire171, clk, reg113, reg82, reg142, reg104);
  assign wire173 = reg103[(4'hb):(4'ha)];
  assign wire174 = reg37[(2'h3):(2'h3)];
  always
    @(posedge clk) begin
      for (forvar175 = (1'h0); (forvar175 < (2'h3)); forvar175 = (forvar175 + (1'h1)))
        begin
          for (forvar176 = (1'h0); (forvar176 < (1'h1)); forvar176 = (forvar176 + (1'h1)))
            begin
              for (forvar177 = (1'h0); (forvar177 < (1'h1)); forvar177 = (forvar177 + (1'h1)))
                begin
                  reg178 <= reg108[(4'ha):(3'h5)];
                  for (forvar179 = (1'h0); (forvar179 < (2'h3)); forvar179 = (forvar179 + (1'h1)))
                    begin
                      reg180 <= $signed({reg130});
                    end
                  for (forvar181 = (1'h0); (forvar181 < (1'h1)); forvar181 = (forvar181 + (1'h1)))
                    begin
                      reg182 <= $signed((~$unsigned((reg34 + reg152))));
                      reg183 <= reg152;
                    end
                end
              for (forvar184 = (1'h0); (forvar184 < (2'h2)); forvar184 = (forvar184 + (1'h1)))
                begin
                  reg185 <= reg153[(4'h8):(1'h0)];
                  for (forvar186 = (1'h0); (forvar186 < (2'h2)); forvar186 = (forvar186 + (1'h1)))
                    begin
                      reg187 <= $signed((+(~^(reg17 || reg137))));
                      reg188 <= reg43[(4'hd):(1'h0)];
                      reg189 <= reg19[(1'h0):(1'h0)];
                    end
                  for (forvar190 = (1'h0); (forvar190 < (1'h1)); forvar190 = (forvar190 + (1'h1)))
                    begin
                      reg191 <= (8'hb3);
                      reg192 <= forvar181[(2'h3):(1'h1)];
                      reg193 <= (~&$unsigned($signed((&reg25))));
                    end
                end
            end
          for (forvar194 = (1'h0); (forvar194 < (1'h0)); forvar194 = (forvar194 + (1'h1)))
            begin
              reg195 <= reg152;
              for (forvar196 = (1'h0); (forvar196 < (2'h2)); forvar196 = (forvar196 + (1'h1)))
                begin
                  if ($unsigned($signed(reg189[(1'h0):(1'h0)])))
                    begin
                      reg197 <= $signed({({reg42} && (~reg140))});
                    end
                  else
                    begin
                      reg197 <= ($unsigned((^~(reg185 ^ wire8))) ?
                          (&{$signed(reg92)}) : reg105);
                      reg198 <= wire156[(4'h8):(1'h0)];
                      reg199 <= (&reg139);
                    end
                  for (forvar200 = (1'h0); (forvar200 < (2'h2)); forvar200 = (forvar200 + (1'h1)))
                    begin
                      reg201 <= (+(((~^reg61) >> {reg24}) ?
                          $signed($signed(reg119)) : reg182));
                    end
                  for (forvar202 = (1'h0); (forvar202 < (2'h3)); forvar202 = (forvar202 + (1'h1)))
                    begin
                      reg203 <= $signed($signed(reg41));
                    end
                end
              for (forvar204 = (1'h0); (forvar204 < (2'h2)); forvar204 = (forvar204 + (1'h1)))
                begin
                  for (forvar205 = (1'h0); (forvar205 < (1'h0)); forvar205 = (forvar205 + (1'h1)))
                    begin
                      reg206 <= ((($signed(reg46) ?
                          (~^reg197) : wire171) + $signed(reg197)) < $signed($signed(reg40[(1'h1):(1'h0)])));
                    end
                  for (forvar207 = (1'h0); (forvar207 < (1'h0)); forvar207 = (forvar207 + (1'h1)))
                    begin
                      reg208 <= $signed(reg19[(2'h3):(2'h2)]);
                      reg209 <= $unsigned(reg38[(2'h3):(2'h2)]);
                      reg210 <= {(^~reg103)};
                    end
                  if (($unsigned(({reg46} << reg95[(2'h2):(2'h2)])) > {forvar176[(3'h6):(1'h0)]}))
                    begin
                      reg211 <= $unsigned({((reg150 ? (8'hba) : wire8) ?
                              reg133[(3'h5):(3'h5)] : $unsigned(reg178))});
                      reg212 <= ($signed(reg49) - (($unsigned(reg130) ?
                              $unsigned(forvar175) : (&reg82)) ?
                          {{reg112}} : (((8'h9d) ? forvar177 : reg137) ?
                              reg102[(1'h0):(1'h0)] : (reg134 ?
                                  reg30 : reg24))));
                      reg213 <= {(~|(+(!reg211)))};
                      reg214 <= (|reg86[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg211 <= ($unsigned($unsigned({reg116})) == {(~&reg85)});
                      reg212 <= reg146[(1'h0):(1'h0)];
                    end
                  for (forvar215 = (1'h0); (forvar215 < (2'h2)); forvar215 = (forvar215 + (1'h1)))
                    begin
                      reg216 <= {(((reg117 ? reg80 : (8'ha1)) ^~ {reg69}) ?
                              (!reg143) : reg62)};
                      reg217 <= $unsigned(($signed(reg134) >>> {$unsigned(reg50)}));
                      reg218 <= ((~^$signed(reg143[(4'hb):(2'h2)])) ?
                          forvar215[(3'h4):(1'h0)] : ((reg136 * (forvar184 ^~ reg80)) ~^ $unsigned(((8'hba) < (8'hb0)))));
                    end
                end
              for (forvar219 = (1'h0); (forvar219 < (1'h1)); forvar219 = (forvar219 + (1'h1)))
                begin
                  if ($signed((((forvar175 ? (8'ha4) : (8'h9e)) & ((8'hb3) ?
                          reg98 : reg84)) ?
                      $unsigned((&reg94)) : $signed($unsigned(reg15)))))
                    begin
                      reg220 <= reg217;
                      reg221 <= (($unsigned(reg178[(2'h2):(1'h1)]) ?
                          forvar194 : $signed(reg116[(1'h1):(1'h1)])) > ($signed(reg119[(1'h1):(1'h1)]) ~^ ((|reg75) ?
                          (reg133 ? reg144 : reg195) : (&reg61))));
                      reg222 <= $unsigned((~forvar205));
                    end
                  else
                    begin
                      reg220 <= $unsigned(reg183);
                      reg221 <= forvar186[(3'h7):(2'h2)];
                      reg222 <= {(reg98 ?
                              (reg213[(2'h3):(1'h1)] >> $signed(reg109)) : $unsigned(reg98))};
                    end
                  if ((&reg134))
                    begin
                      reg223 <= reg138[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg223 <= $unsigned(reg43[(4'hb):(4'h9)]);
                      reg224 <= $unsigned(($signed($signed((8'ha2))) ?
                          (+reg18[(3'h4):(2'h2)]) : ((reg135 * reg185) >= (reg44 ^~ (8'ha1)))));
                    end
                end
            end
        end
      if ((~(8'hb9)))
        begin
          for (forvar225 = (1'h0); (forvar225 < (2'h2)); forvar225 = (forvar225 + (1'h1)))
            begin
              for (forvar226 = (1'h0); (forvar226 < (1'h1)); forvar226 = (forvar226 + (1'h1)))
                begin
                  for (forvar227 = (1'h0); (forvar227 < (2'h2)); forvar227 = (forvar227 + (1'h1)))
                    begin
                      reg228 <= (~&$unsigned((^(8'ha3))));
                      reg229 <= $unsigned((-(forvar181[(1'h0):(1'h0)] ?
                          $signed(reg214) : {wire9})));
                      reg230 <= ($signed(reg150) || reg42);
                    end
                  for (forvar231 = (1'h0); (forvar231 < (1'h0)); forvar231 = (forvar231 + (1'h1)))
                    begin
                      reg232 <= reg137;
                      reg233 <= reg101[(1'h0):(1'h0)];
                    end
                end
              if ((^reg115))
                begin
                  for (forvar234 = (1'h0); (forvar234 < (1'h1)); forvar234 = (forvar234 + (1'h1)))
                    begin
                      reg235 <= (!reg62);
                      reg236 <= (~&((reg84[(3'h7):(3'h6)] ? {(8'h9f)} : reg42) ?
                          reg84[(4'ha):(2'h3)] : reg198));
                    end
                  for (forvar237 = (1'h0); (forvar237 < (1'h1)); forvar237 = (forvar237 + (1'h1)))
                    begin
                      reg238 <= reg145[(1'h0):(1'h0)];
                      reg239 <= {((reg80 | (~|(8'haf))) >= $unsigned((8'ha5)))};
                      reg240 <= (reg195[(3'h4):(3'h4)] + ({(reg40 ?
                                  reg147 : wire11)} ?
                          $unsigned((reg95 ? reg113 : forvar181)) : reg236));
                      reg241 <= $unsigned($signed(reg229[(3'h5):(3'h4)]));
                    end
                end
              else
                begin
                  for (forvar234 = (1'h0); (forvar234 < (2'h3)); forvar234 = (forvar234 + (1'h1)))
                    begin
                      reg235 <= reg211;
                    end
                  if ((forvar176[(1'h0):(1'h0)] ?
                      $signed((~|(~&reg210))) : $signed($signed(reg24[(1'h1):(1'h0)]))))
                    begin
                      reg236 <= reg45;
                    end
                  else
                    begin
                      reg236 <= reg141[(3'h6):(1'h1)];
                    end
                end
              reg242 <= $unsigned(reg123);
              for (forvar243 = (1'h0); (forvar243 < (1'h0)); forvar243 = (forvar243 + (1'h1)))
                begin
                  for (forvar244 = (1'h0); (forvar244 < (1'h1)); forvar244 = (forvar244 + (1'h1)))
                    begin
                      reg245 <= reg47;
                      reg246 <= reg199[(2'h2):(2'h2)];
                    end
                end
            end
          reg247 <= (-$signed({reg29[(2'h2):(2'h2)]}));
          if (($signed(reg115[(1'h1):(1'h1)]) ?
              reg125[(4'hf):(4'hb)] : $signed(reg41[(1'h0):(1'h0)])))
            begin
              for (forvar248 = (1'h0); (forvar248 < (1'h0)); forvar248 = (forvar248 + (1'h1)))
                begin
                  for (forvar249 = (1'h0); (forvar249 < (1'h1)); forvar249 = (forvar249 + (1'h1)))
                    begin
                      reg250 <= {$unsigned($unsigned($signed(reg151)))};
                      reg251 <= {($unsigned((reg199 ?
                              reg37 : reg103)) || ((reg105 ?
                                  forvar234 : reg88) ?
                              $unsigned(reg144) : (reg180 ? reg29 : reg154)))};
                    end
                  if (((forvar190 ^ {(8'hae)}) > reg116[(2'h2):(2'h2)]))
                    begin
                      reg252 <= reg34[(3'h5):(3'h4)];
                      reg253 <= ((($unsigned(wire171) ?
                          $unsigned(reg104) : {(8'hba)}) ~^ {{reg30}}) >= reg25);
                      reg254 <= {forvar184};
                      reg255 <= $unsigned((((^(8'ha3)) <<< (8'hb4)) ?
                          (~|reg209[(3'h5):(3'h4)]) : {(+forvar205)}));
                    end
                  else
                    begin
                      reg252 <= reg147;
                    end
                  for (forvar256 = (1'h0); (forvar256 < (1'h0)); forvar256 = (forvar256 + (1'h1)))
                    begin
                      reg257 <= reg64;
                      reg258 <= {((~{forvar256}) ?
                              (~&(reg45 != reg59)) : $unsigned((~^reg102)))};
                    end
                  if (reg16[(4'hb):(1'h0)])
                    begin
                      reg259 <= $signed({reg25[(1'h1):(1'h1)]});
                      reg260 <= reg119[(3'h4):(2'h3)];
                      reg261 <= {{(reg191 ? (8'ha9) : reg99)}};
                      reg262 <= reg228[(4'ha):(4'h9)];
                    end
                  else
                    begin
                      reg259 <= ($signed(forvar234[(1'h0):(1'h0)]) ^~ {$unsigned((^~reg149))});
                      reg260 <= (reg212 < ($signed(reg141) || reg210));
                    end
                end
            end
          else
            begin
              for (forvar248 = (1'h0); (forvar248 < (2'h3)); forvar248 = (forvar248 + (1'h1)))
                begin
                  reg249 <= ($signed(wire12) >= reg88);
                  for (forvar250 = (1'h0); (forvar250 < (2'h3)); forvar250 = (forvar250 + (1'h1)))
                    begin
                      reg251 <= ((~(reg142 ?
                          reg235[(1'h1):(1'h0)] : $unsigned(reg191))) >= (((reg130 ?
                          forvar231 : (8'hb0)) > (^wire12)) - reg213));
                      reg252 <= $unsigned((((reg54 ?
                          reg82 : (8'ha0)) <= (&forvar244)) <<< $signed({reg101})));
                      reg253 <= $unsigned((({(8'ha2)} >>> $signed(reg105)) > (reg201 >>> (forvar215 <= reg139))));
                    end
                end
              for (forvar254 = (1'h0); (forvar254 < (1'h1)); forvar254 = (forvar254 + (1'h1)))
                begin
                  for (forvar255 = (1'h0); (forvar255 < (2'h2)); forvar255 = (forvar255 + (1'h1)))
                    begin
                      reg256 <= reg141[(2'h2):(1'h1)];
                      reg257 <= $signed(reg145[(2'h2):(2'h2)]);
                    end
                  for (forvar258 = (1'h0); (forvar258 < (1'h1)); forvar258 = (forvar258 + (1'h1)))
                    begin
                      reg259 <= reg148;
                    end
                  for (forvar260 = (1'h0); (forvar260 < (2'h2)); forvar260 = (forvar260 + (1'h1)))
                    begin
                      reg261 <= reg85[(4'hc):(4'hb)];
                    end
                  for (forvar262 = (1'h0); (forvar262 < (2'h2)); forvar262 = (forvar262 + (1'h1)))
                    begin
                      reg263 <= ($signed((+(forvar184 + (8'hb2)))) || $signed(reg247));
                    end
                end
              reg264 <= $signed({($unsigned(reg29) + reg106)});
            end
        end
      else
        begin
          for (forvar225 = (1'h0); (forvar225 < (1'h0)); forvar225 = (forvar225 + (1'h1)))
            begin
              reg226 <= (reg235[(2'h2):(1'h0)] << (^~reg114[(4'hb):(3'h5)]));
            end
          if ((({$signed(forvar207)} && $unsigned(reg25[(4'h9):(2'h3)])) ?
              reg83[(1'h1):(1'h0)] : (~|($signed((8'hab)) >= reg21[(1'h1):(1'h0)]))))
            begin
              for (forvar227 = (1'h0); (forvar227 < (2'h2)); forvar227 = (forvar227 + (1'h1)))
                begin
                  if (reg241)
                    begin
                      reg228 <= (^~$unsigned((reg214[(3'h5):(3'h4)] ?
                          (forvar176 + reg45) : (~|reg110))));
                      reg229 <= $signed(((~|((8'h9f) ? reg106 : reg250)) ?
                          (8'hb5) : ((!reg83) >>> (reg108 ? reg224 : reg143))));
                      reg230 <= ($unsigned(reg87) - (((wire155 ?
                                  reg212 : wire171) ?
                              $unsigned((8'hab)) : reg77) ?
                          ($signed(reg212) & {reg101}) : $signed(reg137[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg228 <= reg15[(1'h1):(1'h0)];
                      reg229 <= forvar258[(4'hb):(3'h6)];
                      reg230 <= (~|$unsigned($unsigned((8'ha8))));
                    end
                end
              if (((reg217[(1'h0):(1'h0)] ?
                  (reg189 <= (forvar215 ^ reg125)) : wire171) << ((reg37 >= $unsigned(forvar254)) + (+reg45[(4'h8):(3'h4)]))))
                begin
                  reg231 <= (forvar255[(4'h9):(4'h8)] ?
                      ($unsigned((|reg108)) ?
                          ((+(8'h9f)) ?
                              reg144 : (reg21 <= reg222)) : $unsigned((^reg83))) : wire174);
                  for (forvar232 = (1'h0); (forvar232 < (1'h0)); forvar232 = (forvar232 + (1'h1)))
                    begin
                      reg233 <= forvar262;
                      reg234 <= (reg250[(2'h3):(2'h3)] >= (reg54 >= (-$signed(reg185))));
                      reg235 <= (reg43 ?
                          (reg92 ?
                              reg91 : $unsigned((-reg220))) : ((-{reg180}) ^~ {{reg45}}));
                      reg236 <= $unsigned(($signed((reg119 & (8'hb3))) != $signed(((8'hac) - reg125))));
                    end
                  for (forvar237 = (1'h0); (forvar237 < (2'h3)); forvar237 = (forvar237 + (1'h1)))
                    begin
                      reg238 <= (8'ha1);
                      reg239 <= (~&forvar175);
                    end
                end
              else
                begin
                  if (($unsigned($signed((reg69 ?
                      (8'h9e) : reg218))) == (((reg221 ?
                          reg48 : reg29) * (forvar219 ? reg31 : wire11)) ?
                      (^$unsigned(reg153)) : ($signed(reg206) ?
                          (8'hb7) : reg29[(4'hd):(4'hb)]))))
                    begin
                      reg231 <= (({(8'ha5)} == $signed((wire7 && reg253))) ?
                          (+$signed({reg115})) : $unsigned((+(wire155 ?
                              reg95 : forvar204))));
                      reg232 <= (&reg251);
                      reg233 <= ($signed($unsigned((~^forvar260))) ?
                          {($signed(reg234) >= $unsigned((8'h9d)))} : forvar196);
                    end
                  else
                    begin
                      reg231 <= (~^reg208);
                      reg232 <= reg82;
                      reg233 <= reg193[(2'h2):(1'h1)];
                    end
                  for (forvar234 = (1'h0); (forvar234 < (2'h2)); forvar234 = (forvar234 + (1'h1)))
                    begin
                      reg235 <= ({$signed((forvar244 ? reg42 : reg41))} ?
                          reg125 : reg235);
                      reg236 <= ((reg101[(4'h8):(3'h7)] | $unsigned((reg142 >>> (8'hac)))) ?
                          wire174[(4'h9):(3'h7)] : $unsigned((-(~^reg233))));
                    end
                end
              reg240 <= reg61[(3'h5):(2'h3)];
              for (forvar241 = (1'h0); (forvar241 < (1'h0)); forvar241 = (forvar241 + (1'h1)))
                begin
                  for (forvar242 = (1'h0); (forvar242 < (1'h0)); forvar242 = (forvar242 + (1'h1)))
                    begin
                      reg243 <= $unsigned($unsigned((-reg92[(1'h0):(1'h0)])));
                      reg244 <= {(forvar196[(2'h3):(2'h3)] != $signed((reg214 >>> reg48)))};
                    end
                  for (forvar245 = (1'h0); (forvar245 < (2'h2)); forvar245 = (forvar245 + (1'h1)))
                    begin
                      reg246 <= $signed(reg52[(2'h3):(2'h2)]);
                      reg247 <= (^~(-((8'hb7) ?
                          $unsigned((8'ha4)) : (~|reg25))));
                      reg248 <= (&{$unsigned((reg48 ? reg211 : forvar260))});
                    end
                  for (forvar249 = (1'h0); (forvar249 < (2'h2)); forvar249 = (forvar249 + (1'h1)))
                    begin
                      reg250 <= $signed((&{(+reg50)}));
                      reg251 <= reg36;
                    end
                end
            end
          else
            begin
              if ((^~((8'hae) >> (reg120[(2'h3):(1'h1)] ?
                  $signed(reg23) : (&wire7)))))
                begin
                  for (forvar227 = (1'h0); (forvar227 < (2'h3)); forvar227 = (forvar227 + (1'h1)))
                    begin
                      reg228 <= $unsigned(((+(reg148 & reg151)) ?
                          forvar243[(2'h3):(2'h2)] : (|$unsigned(reg260))));
                      reg229 <= reg150[(3'h5):(2'h3)];
                      reg230 <= (forvar248 ?
                          ($signed((reg34 >>> wire9)) ?
                              reg28 : {reg233[(1'h1):(1'h1)]}) : $signed($signed(reg114[(3'h5):(2'h2)])));
                    end
                  reg231 <= reg92[(2'h2):(2'h2)];
                  if (((((reg154 ~^ (8'hb8)) >= $signed(reg206)) ?
                      ($unsigned(reg47) || {reg72}) : reg221[(3'h4):(1'h1)]) <<< (^($unsigned((8'ha0)) ?
                      reg223[(3'h5):(2'h3)] : $unsigned(reg40)))))
                    begin
                      reg232 <= reg31[(3'h5):(2'h2)];
                      reg233 <= reg130[(4'he):(3'h4)];
                      reg234 <= ($unsigned($signed($unsigned(reg198))) ^ ($signed((reg63 >> wire173)) == ((8'hb5) ?
                          $unsigned(reg38) : (reg73 ? forvar176 : reg77))));
                    end
                  else
                    begin
                      reg232 <= $signed({reg46});
                      reg233 <= $unsigned($signed((&reg235)));
                      reg234 <= (reg141[(4'hb):(4'hb)] + reg61[(4'h9):(3'h4)]);
                      reg235 <= forvar262[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  reg227 <= reg129;
                  for (forvar228 = (1'h0); (forvar228 < (2'h2)); forvar228 = (forvar228 + (1'h1)))
                    begin
                      reg229 <= ({($unsigned(reg52) ?
                                  wire171[(1'h0):(1'h0)] : (wire155 ?
                                      reg212 : reg212))} ?
                          reg144[(1'h0):(1'h0)] : $signed((|(!forvar181))));
                      reg230 <= (((((8'ha7) != forvar181) >= $signed(wire174)) << $unsigned($signed((8'h9f)))) == ($unsigned(reg252) && reg64[(3'h5):(3'h5)]));
                      reg231 <= $unsigned(({(reg261 ? reg234 : reg21)} ?
                          $signed($unsigned(reg21)) : (reg97 ?
                              reg32[(4'h8):(3'h6)] : (8'ha9))));
                      reg232 <= $signed(($signed(reg137[(1'h0):(1'h0)]) ?
                          $unsigned(reg123[(1'h1):(1'h1)]) : reg144[(4'h9):(3'h6)]));
                    end
                  for (forvar233 = (1'h0); (forvar233 < (1'h1)); forvar233 = (forvar233 + (1'h1)))
                    begin
                      reg234 <= $signed((reg62[(2'h2):(1'h1)] << $unsigned(reg27[(3'h4):(2'h3)])));
                      reg235 <= reg254[(1'h0):(1'h0)];
                      reg236 <= reg102;
                    end
                  for (forvar237 = (1'h0); (forvar237 < (2'h2)); forvar237 = (forvar237 + (1'h1)))
                    begin
                      reg238 <= $unsigned($unsigned(((^~reg135) <= (+(8'ha6)))));
                    end
                end
              for (forvar239 = (1'h0); (forvar239 < (1'h1)); forvar239 = (forvar239 + (1'h1)))
                begin
                  if ($unsigned((^~(forvar248[(2'h2):(1'h0)] != (~forvar228)))))
                    begin
                      reg240 <= (8'ha1);
                      reg241 <= $unsigned(reg49);
                      reg242 <= {reg52[(3'h7):(2'h2)]};
                    end
                  else
                    begin
                      reg240 <= (^(forvar176[(2'h2):(1'h1)] != ((~|(8'ha1)) >= (|(8'hb5)))));
                      reg241 <= $unsigned(((~|(&reg116)) ?
                          (^~reg230[(2'h2):(1'h0)]) : $unsigned($unsigned(reg203))));
                    end
                  for (forvar243 = (1'h0); (forvar243 < (2'h2)); forvar243 = (forvar243 + (1'h1)))
                    begin
                      reg244 <= ({reg189} - ($signed(reg41) ?
                          $unsigned((reg148 ? (8'hb7) : (8'hb5))) : forvar255));
                    end
                  for (forvar245 = (1'h0); (forvar245 < (2'h2)); forvar245 = (forvar245 + (1'h1)))
                    begin
                      reg246 <= ((forvar258 ?
                          (forvar260[(2'h2):(1'h1)] ?
                              (reg24 ?
                                  (8'ha8) : (8'ha7)) : reg231[(3'h6):(1'h0)]) : reg36) - $signed({(&forvar243)}));
                      reg247 <= (^(~|$unsigned((reg59 * forvar255))));
                      reg248 <= $signed((^~reg150[(3'h5):(3'h4)]));
                    end
                  for (forvar249 = (1'h0); (forvar249 < (1'h0)); forvar249 = (forvar249 + (1'h1)))
                    begin
                      reg250 <= $unsigned((reg77 | $unsigned({reg223})));
                      reg251 <= (8'hab);
                    end
                end
            end
          reg252 <= {((8'hb5) ? $signed(reg113) : {reg98})};
          for (forvar253 = (1'h0); (forvar253 < (2'h3)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 <= $unsigned({(((8'hb9) <<< (8'ha2)) * reg149)});
              for (forvar255 = (1'h0); (forvar255 < (1'h0)); forvar255 = (forvar255 + (1'h1)))
                begin
                  for (forvar256 = (1'h0); (forvar256 < (2'h2)); forvar256 = (forvar256 + (1'h1)))
                    begin
                      reg257 <= $unsigned(reg73[(1'h1):(1'h1)]);
                      reg258 <= $unsigned((((reg25 ? (8'ha9) : reg21) ?
                              (~(8'haa)) : {reg213}) ?
                          reg208[(1'h0):(1'h0)] : ((reg42 ? reg112 : reg235) ?
                              (reg111 < wire9) : $signed((8'h9e)))));
                      reg259 <= ($signed((&{forvar242})) ?
                          $signed(wire11) : (reg192 ?
                              forvar231 : ((8'ha7) ? forvar204 : wire13)));
                    end
                end
              for (forvar260 = (1'h0); (forvar260 < (1'h1)); forvar260 = (forvar260 + (1'h1)))
                begin
                  for (forvar261 = (1'h0); (forvar261 < (1'h0)); forvar261 = (forvar261 + (1'h1)))
                    begin
                      reg262 <= reg191[(4'hd):(2'h2)];
                      reg263 <= $signed((8'ha2));
                      reg264 <= ((+forvar181[(2'h2):(1'h0)]) | (({forvar234} * {reg242}) ?
                          (~(reg123 ?
                              reg140 : reg144)) : $unsigned($unsigned(reg153))));
                    end
                end
            end
        end
      for (forvar265 = (1'h0); (forvar265 < (1'h0)); forvar265 = (forvar265 + (1'h1)))
        begin
          reg266 <= ($unsigned(reg111) ?
              (forvar228 <<< ($signed(wire9) ~^ $signed(reg63))) : {(reg101[(3'h4):(1'h1)] <<< (&(8'hae)))});
          for (forvar267 = (1'h0); (forvar267 < (2'h2)); forvar267 = (forvar267 + (1'h1)))
            begin
              for (forvar268 = (1'h0); (forvar268 < (2'h3)); forvar268 = (forvar268 + (1'h1)))
                begin
                  for (forvar269 = (1'h0); (forvar269 < (2'h2)); forvar269 = (forvar269 + (1'h1)))
                    begin
                      reg270 <= forvar175[(3'h5):(2'h2)];
                      reg271 <= $signed((!forvar250));
                      reg272 <= ({$signed($signed(reg118))} << {((reg80 && (8'hb7)) - $unsigned((8'hab)))});
                      reg273 <= ($unsigned({reg226[(3'h4):(2'h3)]}) ?
                          (&reg240[(3'h6):(2'h2)]) : forvar256[(2'h3):(1'h0)]);
                    end
                  for (forvar274 = (1'h0); (forvar274 < (2'h2)); forvar274 = (forvar274 + (1'h1)))
                    begin
                      reg275 <= reg148;
                      reg276 <= reg24;
                      reg277 <= (((-$unsigned(reg104)) >>> (forvar190 | (reg271 ?
                              reg40 : reg16))) ?
                          ({(~reg45)} ?
                              (~|(forvar202 || reg110)) : ($unsigned(reg47) ?
                                  (reg130 <<< forvar231) : {(8'hb2)})) : ({(reg224 >> reg257)} ?
                              $signed((8'h9f)) : (reg47[(3'h5):(2'h2)] ?
                                  $unsigned(forvar253) : $unsigned((8'hab)))));
                    end
                  if ((reg45[(1'h0):(1'h0)] ?
                      reg212[(1'h0):(1'h0)] : forvar255[(3'h7):(3'h7)]))
                    begin
                      reg278 <= reg188[(2'h2):(2'h2)];
                      reg279 <= {($unsigned($unsigned(reg65)) ~^ $unsigned((reg55 ?
                              (8'hac) : forvar204)))};
                      reg280 <= reg118[(3'h7):(1'h0)];
                    end
                  else
                    begin
                      reg278 <= $signed((~&$unsigned(forvar258[(3'h5):(1'h1)])));
                      reg279 <= $unsigned($signed({$unsigned(reg36)}));
                    end
                  reg281 <= (|$unsigned($signed((reg41 + reg23))));
                end
              for (forvar282 = (1'h0); (forvar282 < (2'h2)); forvar282 = (forvar282 + (1'h1)))
                begin
                  if ((~^(reg25 & reg262)))
                    begin
                      reg283 <= $unsigned((-{wire8}));
                      reg284 <= forvar245;
                      reg285 <= reg236;
                    end
                  else
                    begin
                      reg283 <= $unsigned($signed(((forvar239 ?
                          (8'ha7) : (8'hb6)) ^ (reg57 ? wire12 : reg53))));
                    end
                  for (forvar286 = (1'h0); (forvar286 < (1'h0)); forvar286 = (forvar286 + (1'h1)))
                    begin
                      reg287 <= $unsigned((|{(8'hac)}));
                      reg288 <= (^~$signed((8'hba)));
                      reg289 <= reg95;
                      reg290 <= ((wire10 ?
                          (+(~&reg246)) : ((~^reg36) >> reg230[(1'h1):(1'h0)])) != $signed($unsigned({reg82})));
                    end
                  for (forvar291 = (1'h0); (forvar291 < (1'h0)); forvar291 = (forvar291 + (1'h1)))
                    begin
                      reg292 <= $unsigned(reg20);
                      reg293 <= ((reg208[(2'h3):(1'h1)] ?
                              (~|reg33[(2'h2):(1'h0)]) : {(-forvar243)}) ?
                          $unsigned($unsigned($unsigned((8'ha8)))) : $signed($signed((reg227 ?
                              reg92 : reg84))));
                    end
                end
              reg294 <= (((reg235 ?
                  $unsigned(reg187) : forvar261[(3'h4):(2'h2)]) << $unsigned($unsigned(reg20))) ~^ {$unsigned((reg122 ?
                      wire174 : reg218))});
              if ((~&reg72))
                begin
                  for (forvar295 = (1'h0); (forvar295 < (1'h0)); forvar295 = (forvar295 + (1'h1)))
                    begin
                      reg296 <= $unsigned($unsigned($unsigned((forvar261 - reg101))));
                    end
                end
              else
                begin
                  for (forvar295 = (1'h0); (forvar295 < (1'h1)); forvar295 = (forvar295 + (1'h1)))
                    begin
                      reg296 <= reg258;
                      reg297 <= reg139[(3'h6):(1'h0)];
                      reg298 <= {reg71[(1'h0):(1'h0)]};
                      reg299 <= $signed(reg272);
                    end
                  if ((^~($signed((reg110 == reg124)) ?
                      ({reg234} ? wire174[(4'hc):(4'h9)] : {reg97}) : reg36)))
                    begin
                      reg300 <= (reg224 < ((8'ha0) ~^ {(8'ha5)}));
                      reg301 <= $signed($signed($unsigned(reg288)));
                      reg302 <= reg120[(3'h6):(1'h1)];
                      reg303 <= $unsigned($signed($signed(reg75)));
                    end
                  else
                    begin
                      reg300 <= $signed($unsigned(reg297[(3'h7):(1'h1)]));
                      reg301 <= $signed($unsigned((|reg209)));
                      reg302 <= (~&(~(reg86 ?
                          reg42[(3'h7):(3'h6)] : (forvar184 ?
                              reg27 : reg199))));
                      reg303 <= ((^~(reg250[(2'h2):(2'h2)] ?
                              forvar207 : $signed(reg303))) ?
                          (~^((reg48 ?
                              reg29 : forvar256) != reg278)) : reg80[(2'h3):(1'h1)]);
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned((reg78 > ($signed(reg252) ? reg135 : {(8'hb3)}))))
        begin
          if ({((&(^~(8'hb4))) <= (8'h9d))})
            begin
              reg304 <= $signed({$signed($unsigned((8'hab)))});
              if (($signed($unsigned($unsigned((8'hb4)))) ^~ ((|reg289[(2'h3):(1'h0)]) && reg28[(4'h9):(3'h5)])))
                begin
                  for (forvar305 = (1'h0); (forvar305 < (1'h1)); forvar305 = (forvar305 + (1'h1)))
                    begin
                      reg306 <= ((reg100[(4'h8):(3'h4)] ?
                          $unsigned(reg57) : ({reg146} ?
                              reg122[(3'h6):(3'h4)] : (reg246 ?
                                  wire171 : reg111))) + $signed((|(^~reg36))));
                      reg307 <= (reg103 && reg83);
                      reg308 <= (8'h9c);
                    end
                  for (forvar309 = (1'h0); (forvar309 < (2'h2)); forvar309 = (forvar309 + (1'h1)))
                    begin
                      reg310 <= reg188[(2'h2):(1'h0)];
                      reg311 <= reg246[(3'h7):(3'h7)];
                      reg312 <= $unsigned(reg183);
                      reg313 <= {reg29[(4'hb):(4'hb)]};
                    end
                  reg314 <= reg101;
                  for (forvar315 = (1'h0); (forvar315 < (1'h1)); forvar315 = (forvar315 + (1'h1)))
                    begin
                      reg316 <= (~^reg85[(1'h1):(1'h1)]);
                      reg317 <= reg44;
                    end
                end
              else
                begin
                  reg305 <= reg33[(1'h1):(1'h1)];
                end
              for (forvar318 = (1'h0); (forvar318 < (1'h0)); forvar318 = (forvar318 + (1'h1)))
                begin
                  if ((-$signed(($unsigned(reg272) != (~|(8'hb9))))))
                    begin
                      reg319 <= ((({reg236} || $unsigned(reg260)) ?
                              $signed($signed(reg201)) : (&(reg229 ?
                                  reg42 : (8'h9f)))) ?
                          reg195 : reg306[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg319 <= ($signed(reg281) * ($signed($signed(reg307)) ?
                          (reg18 ?
                              (reg73 << reg142) : (&(8'ha0))) : $unsigned($signed((8'hab)))));
                      reg320 <= {(+{$unsigned(reg259)})};
                      reg321 <= {$unsigned((~^reg255[(3'h5):(3'h4)]))};
                      reg322 <= (~^(($signed(reg146) ~^ ((8'hb1) ?
                              reg33 : (8'hab))) ?
                          $unsigned((8'ha5)) : {(8'ha9)}));
                    end
                  reg323 <= reg308;
                  reg324 <= ((~&reg260[(3'h5):(1'h0)]) == reg144[(2'h2):(1'h0)]);
                  for (forvar325 = (1'h0); (forvar325 < (2'h2)); forvar325 = (forvar325 + (1'h1)))
                    begin
                      reg326 <= {{reg251}};
                      reg327 <= (&(~&wire173[(3'h4):(2'h3)]));
                      reg328 <= ((+reg275[(3'h7):(1'h0)]) & (-($unsigned((8'ha4)) <<< (8'h9c))));
                    end
                end
            end
          else
            begin
              for (forvar304 = (1'h0); (forvar304 < (1'h1)); forvar304 = (forvar304 + (1'h1)))
                begin
                  for (forvar305 = (1'h0); (forvar305 < (1'h0)); forvar305 = (forvar305 + (1'h1)))
                    begin
                      reg306 <= reg238[(1'h0):(1'h0)];
                      reg307 <= (reg143[(3'h4):(1'h1)] == reg37[(3'h6):(1'h1)]);
                      reg308 <= (8'hb5);
                    end
                  if (reg183)
                    begin
                      reg309 <= ($unsigned(reg64[(3'h6):(2'h3)]) ?
                          $signed($unsigned({reg224})) : (&$unsigned($unsigned((8'haa)))));
                      reg310 <= (|($unsigned($unsigned(reg38)) + {$unsigned(reg61)}));
                      reg311 <= (~$unsigned(((reg78 << reg210) ?
                          (reg312 > reg48) : $signed(reg141))));
                      reg312 <= ($unsigned(reg61[(2'h2):(2'h2)]) ?
                          ({$unsigned(reg313)} ?
                              (reg210[(2'h2):(1'h1)] ?
                                  reg149[(2'h2):(1'h1)] : reg238[(3'h5):(2'h3)]) : (&reg254)) : (8'hab));
                    end
                  else
                    begin
                      reg309 <= wire7;
                    end
                  for (forvar313 = (1'h0); (forvar313 < (1'h0)); forvar313 = (forvar313 + (1'h1)))
                    begin
                      reg314 <= $signed($signed((reg275 > (reg233 << reg105))));
                      reg315 <= $signed((($signed((8'hb0)) == $unsigned(wire13)) << $unsigned(reg203[(4'hd):(4'hb)])));
                    end
                end
              reg316 <= ($signed(reg130) == reg28);
              if ($unsigned((~^(8'hb4))))
                begin
                  for (forvar317 = (1'h0); (forvar317 < (2'h3)); forvar317 = (forvar317 + (1'h1)))
                    begin
                      reg318 <= $unsigned({reg21[(1'h0):(1'h0)]});
                    end
                  for (forvar319 = (1'h0); (forvar319 < (1'h1)); forvar319 = (forvar319 + (1'h1)))
                    begin
                      reg320 <= (^~$unsigned($signed($unsigned((8'ha5)))));
                      reg321 <= reg266;
                      reg322 <= {$unsigned((8'ha4))};
                      reg323 <= (($unsigned(reg281[(3'h6):(2'h3)]) ?
                              $signed({reg213}) : (~&wire173)) ?
                          (($unsigned((8'ha5)) - $unsigned(reg63)) > $signed($signed(reg84))) : {(reg52 ^~ $unsigned((8'hb5)))});
                    end
                  for (forvar324 = (1'h0); (forvar324 < (1'h0)); forvar324 = (forvar324 + (1'h1)))
                    begin
                      reg325 <= reg53[(3'h5):(3'h4)];
                      reg326 <= $unsigned({reg199});
                      reg327 <= ((((reg145 ? (8'hba) : reg252) ?
                                  reg216 : (reg239 ? reg64 : reg236)) ?
                              $signed($signed(reg261)) : $signed($unsigned(reg65))) ?
                          ($signed(((8'hb2) << reg298)) ?
                              (&$unsigned(reg150)) : (reg32 >> $unsigned(reg234))) : {reg145});
                      reg328 <= ($signed($signed({reg104})) ?
                          $signed(((reg188 ? reg189 : reg233) ?
                              reg135 : reg43)) : reg307[(1'h0):(1'h0)]);
                    end
                  if ($signed({((-reg296) && {(8'hb4)})}))
                    begin
                      reg329 <= (+(reg242[(4'hc):(4'h9)] ?
                          $unsigned($unsigned(reg139)) : reg154));
                    end
                  else
                    begin
                      reg329 <= $signed(forvar304);
                      reg330 <= wire156;
                      reg331 <= reg95[(2'h2):(1'h1)];
                    end
                end
              else
                begin
                  if ($unsigned(({(+reg185)} ?
                      (~^$unsigned(reg277)) : (&{reg301}))))
                    begin
                      reg317 <= ((($unsigned(reg38) && (~^reg185)) ?
                              ($unsigned((8'hb4)) || $unsigned(reg240)) : ((reg302 ?
                                      reg258 : (8'ha0)) ?
                                  ((8'ha1) ?
                                      reg301 : reg293) : $unsigned(reg130))) ?
                          ((reg154[(1'h1):(1'h0)] >>> reg257[(3'h5):(3'h5)]) ?
                              (reg249[(3'h5):(2'h3)] ?
                                  {reg153} : $unsigned(forvar325)) : $signed(reg244[(2'h3):(1'h1)])) : (reg119 ~^ $unsigned($signed(reg147))));
                      reg318 <= reg91;
                      reg319 <= ($unsigned({{reg182}}) && $unsigned(($unsigned(reg24) ?
                          (reg46 ? reg130 : reg302) : (reg259 & reg257))));
                    end
                  else
                    begin
                      reg317 <= (reg303[(2'h2):(1'h1)] ?
                          ((~(reg15 << reg323)) && reg187) : $signed(reg330[(1'h0):(1'h0)]));
                    end
                  if (reg221)
                    begin
                      reg320 <= reg308;
                    end
                  else
                    begin
                      reg320 <= reg23;
                      reg321 <= reg221;
                      reg322 <= (((+$signed(reg122)) || $signed(((8'hb4) ^~ reg299))) | {$unsigned((|reg110))});
                      reg323 <= {($signed(((8'hb1) ? reg305 : (8'ha5))) ?
                              reg206[(3'h4):(1'h1)] : $unsigned((^reg249)))};
                    end
                end
              if ($signed($signed($signed({(8'had)}))))
                begin
                  for (forvar332 = (1'h0); (forvar332 < (1'h1)); forvar332 = (forvar332 + (1'h1)))
                    begin
                      reg333 <= $signed($unsigned(reg80[(2'h3):(1'h1)]));
                    end
                end
              else
                begin
                  reg332 <= (~^reg43[(3'h5):(1'h1)]);
                  if (((!reg314) ?
                      $signed($unsigned({(8'ha0)})) : $signed((reg130[(1'h1):(1'h1)] || (-reg16)))))
                    begin
                      reg333 <= ((+(|{(8'hb9)})) <= $signed($unsigned($unsigned(reg329))));
                      reg334 <= $signed(reg144[(1'h0):(1'h0)]);
                      reg335 <= reg258[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg333 <= $signed((|$signed((reg35 * reg224))));
                      reg334 <= reg271;
                    end
                  if ($unsigned(reg325[(4'h8):(1'h0)]))
                    begin
                      reg336 <= {{((reg314 & reg214) ?
                                  {reg201} : (reg78 != (8'hb0)))}};
                      reg337 <= (&(reg246[(4'hb):(4'hb)] ?
                          $unsigned((reg258 + reg240)) : (-(8'ha5))));
                    end
                  else
                    begin
                      reg336 <= $unsigned(({reg78[(3'h5):(3'h5)]} ?
                          $signed((^~reg92)) : (~^(^~reg119))));
                      reg337 <= (~|reg322);
                    end
                  if ({wire155})
                    begin
                      reg338 <= ($unsigned((~^(^reg153))) ^ (!$signed((reg301 ?
                          reg34 : reg146))));
                    end
                  else
                    begin
                      reg338 <= $unsigned($signed(($signed(reg100) != (reg30 >> (8'hac)))));
                      reg339 <= reg333[(2'h3):(2'h2)];
                      reg340 <= reg232[(4'hc):(1'h0)];
                    end
                end
            end
          if ({(+($signed(reg241) ? reg338 : $unsigned((8'ha0))))})
            begin
              for (forvar341 = (1'h0); (forvar341 < (2'h2)); forvar341 = (forvar341 + (1'h1)))
                begin
                  for (forvar342 = (1'h0); (forvar342 < (1'h1)); forvar342 = (forvar342 + (1'h1)))
                    begin
                      reg343 <= (reg113[(2'h3):(2'h3)] ~^ ((reg257 >>> (~&forvar324)) ?
                          $unsigned(forvar325[(1'h0):(1'h0)]) : $signed((reg86 > reg35))));
                      reg344 <= reg246;
                    end
                end
              for (forvar345 = (1'h0); (forvar345 < (1'h0)); forvar345 = (forvar345 + (1'h1)))
                begin
                  if ((($signed(reg214) <<< $signed((reg198 ?
                          reg44 : (8'ha2)))) ?
                      (reg48[(1'h1):(1'h0)] << $unsigned($unsigned(reg102))) : (|forvar315)))
                    begin
                      reg346 <= (^~$signed(($unsigned((8'hac)) ?
                          $unsigned(reg143) : (reg124 || forvar309))));
                      reg347 <= ($signed({$signed(reg19)}) ?
                          (^~(^~(reg139 ?
                              reg153 : (8'ha5)))) : ((~&reg289[(3'h6):(2'h3)]) ?
                              $unsigned(((8'hb0) & wire11)) : wire13));
                    end
                  else
                    begin
                      reg346 <= $signed((($unsigned(reg148) << reg324) ?
                          (|(forvar315 ? reg278 : reg294)) : $signed((reg43 ?
                              reg134 : reg195))));
                      reg347 <= {reg315[(3'h7):(2'h3)]};
                      reg348 <= (((~^reg285) == {reg135}) ~^ (((-wire8) * reg104) && (|$signed(reg319))));
                    end
                  for (forvar349 = (1'h0); (forvar349 < (2'h2)); forvar349 = (forvar349 + (1'h1)))
                    begin
                      reg350 <= (~|(wire174[(4'ha):(4'ha)] - reg28));
                      reg351 <= reg328;
                    end
                end
              reg352 <= ({$unsigned((&reg212))} ?
                  $signed(reg182) : ((&(~^(8'ha7))) + {reg302}));
              if ($signed((~reg141[(1'h1):(1'h1)])))
                begin
                  reg353 <= reg302[(1'h1):(1'h0)];
                  if ($unsigned(((8'ha4) ?
                      forvar341 : ($signed(reg182) ?
                          reg81 : reg105[(3'h5):(3'h5)]))))
                    begin
                      reg354 <= $signed(reg135);
                      reg355 <= $signed((((reg154 > (8'ha2)) ?
                          reg317[(1'h1):(1'h0)] : {reg264}) && (reg312 * reg180[(1'h1):(1'h1)])));
                      reg356 <= reg318;
                    end
                  else
                    begin
                      reg354 <= reg260;
                    end
                  if (reg18)
                    begin
                      reg357 <= $signed((~|(reg309[(1'h0):(1'h0)] ?
                          (forvar341 ?
                              (8'hae) : reg300) : reg86[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg357 <= ($unsigned(reg292) > reg17);
                      reg358 <= $unsigned({((^~reg86) ? (!reg354) : {reg344})});
                    end
                  reg359 <= reg35[(1'h1):(1'h1)];
                end
              else
                begin
                  for (forvar353 = (1'h0); (forvar353 < (1'h0)); forvar353 = (forvar353 + (1'h1)))
                    begin
                      reg354 <= $signed(((~^reg54) ?
                          $unsigned(wire155[(2'h3):(1'h1)]) : $signed($signed(reg236))));
                    end
                end
            end
          else
            begin
              if ($signed((^~reg189)))
                begin
                  for (forvar341 = (1'h0); (forvar341 < (2'h2)); forvar341 = (forvar341 + (1'h1)))
                    begin
                      reg342 <= {((!(reg152 ?
                              reg301 : reg108)) ^~ {reg151[(1'h1):(1'h1)]})};
                      reg343 <= reg199[(4'hd):(1'h1)];
                      reg344 <= ((reg182[(2'h2):(1'h1)] | $unsigned((reg340 ?
                              (8'hb1) : (8'ha1)))) ?
                          (forvar318[(4'ha):(4'h9)] * reg262[(3'h5):(3'h4)]) : ((^{reg122}) ?
                              ($signed(reg23) ~^ {reg262}) : (reg139[(1'h1):(1'h0)] ?
                                  (8'ha1) : (reg140 - reg235))));
                      reg345 <= reg33[(2'h3):(1'h1)];
                    end
                  if (reg347)
                    begin
                      reg346 <= $signed((-(+(8'hb8))));
                      reg347 <= reg287;
                      reg348 <= $signed(reg238);
                      reg349 <= $unsigned($unsigned((~^reg115[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg346 <= {($signed(reg236) <= ($signed(reg303) ?
                              $unsigned((8'ha0)) : (reg232 || reg100)))};
                      reg347 <= ($signed(reg106[(2'h3):(2'h3)]) <= reg32);
                    end
                  reg350 <= (8'hb0);
                  if (reg235)
                    begin
                      reg351 <= reg137;
                    end
                  else
                    begin
                      reg351 <= (reg302[(2'h3):(1'h1)] & reg146[(2'h2):(2'h2)]);
                      reg352 <= $signed(reg84);
                    end
                end
              else
                begin
                  for (forvar341 = (1'h0); (forvar341 < (1'h1)); forvar341 = (forvar341 + (1'h1)))
                    begin
                      reg342 <= ((($signed((8'hb5)) ?
                              reg37 : $unsigned(reg276)) + ((reg328 ?
                                  reg333 : reg236) ?
                              $signed(reg249) : reg198[(4'h8):(3'h5)])) ?
                          reg41 : (((reg118 ? forvar319 : reg50) ?
                                  reg98 : $signed(reg272)) ?
                              {(reg43 ? reg101 : reg78)} : ((reg247 ?
                                  reg201 : (8'hae)) >= reg85[(2'h3):(2'h2)])));
                      reg343 <= (!$signed($signed((~&reg307))));
                    end
                  reg344 <= {$unsigned((~^(wire12 ? (8'hb8) : (8'h9e))))};
                  if (((!$unsigned((reg82 ~^ (8'h9c)))) == ({((8'hb0) ?
                          reg130 : reg180)} <= {reg272})))
                    begin
                      reg345 <= (8'ha0);
                    end
                  else
                    begin
                      reg345 <= $unsigned(($signed((reg283 - reg193)) ?
                          (|$signed(reg52)) : (8'hac)));
                      reg346 <= ((|(~|$signed(reg234))) ?
                          $signed({(&reg48)}) : reg319[(3'h5):(2'h2)]);
                      reg347 <= $unsigned($unsigned(((^reg34) << $unsigned(reg246))));
                      reg348 <= (reg213 * ((&(-reg324)) ?
                          (~(|(8'ha7))) : (~&(reg62 ? reg220 : reg34))));
                    end
                end
              for (forvar353 = (1'h0); (forvar353 < (2'h3)); forvar353 = (forvar353 + (1'h1)))
                begin
                  if (reg314[(4'hc):(2'h2)])
                    begin
                      reg354 <= $signed($unsigned($signed((-reg129))));
                      reg355 <= ($signed((~|reg25[(2'h2):(1'h0)])) ?
                          $signed({reg210[(4'h8):(3'h4)]}) : $signed({(reg357 ?
                                  reg259 : reg249)}));
                      reg356 <= (((~&$signed((8'hb7))) ?
                          $unsigned(reg296) : reg99) >= reg335);
                    end
                  else
                    begin
                      reg354 <= reg275;
                      reg355 <= $signed($signed({(reg218 ? reg45 : reg189)}));
                      reg356 <= ($signed($unsigned(((8'haa) ?
                              reg335 : reg284))) ?
                          reg278[(1'h0):(1'h0)] : reg224);
                      reg357 <= (8'hae);
                    end
                  for (forvar358 = (1'h0); (forvar358 < (2'h3)); forvar358 = (forvar358 + (1'h1)))
                    begin
                      reg359 <= {reg261[(2'h3):(1'h0)]};
                      reg360 <= (!(^((reg358 ? reg111 : reg21) ?
                          reg216[(1'h1):(1'h0)] : $signed(reg18))));
                      reg361 <= $unsigned($signed($unsigned((+(8'hb6)))));
                    end
                  reg362 <= (+(($unsigned(reg297) ?
                      (^reg259) : {reg15}) - reg54));
                  for (forvar363 = (1'h0); (forvar363 < (2'h2)); forvar363 = (forvar363 + (1'h1)))
                    begin
                      reg364 <= (&$signed((~|reg105[(1'h1):(1'h0)])));
                      reg365 <= (8'ha9);
                    end
                end
            end
          if (((8'hb6) - (~^forvar349)))
            begin
              for (forvar366 = (1'h0); (forvar366 < (2'h3)); forvar366 = (forvar366 + (1'h1)))
                begin
                  for (forvar367 = (1'h0); (forvar367 < (1'h0)); forvar367 = (forvar367 + (1'h1)))
                    begin
                      reg368 <= reg62;
                      reg369 <= ((^~(reg115 ? (|reg183) : $unsigned(reg193))) ?
                          $signed((reg249 != (reg82 != reg125))) : (|$unsigned(forvar366[(3'h4):(1'h1)])));
                      reg370 <= (!({reg40[(2'h3):(1'h1)]} ?
                          reg78[(3'h6):(1'h0)] : reg91));
                      reg371 <= reg104;
                    end
                  for (forvar372 = (1'h0); (forvar372 < (2'h3)); forvar372 = (forvar372 + (1'h1)))
                    begin
                      reg373 <= reg285;
                      reg374 <= ($unsigned($signed($signed(reg148))) == reg49);
                      reg375 <= {(((reg346 + reg192) ?
                                  (reg347 ?
                                      reg136 : reg299) : reg143[(4'hb):(4'ha)]) ?
                              (8'hb3) : ((reg34 >> (8'hac)) ?
                                  {reg333} : reg317))};
                    end
                  reg376 <= (&$unsigned(reg206));
                end
            end
          else
            begin
              for (forvar366 = (1'h0); (forvar366 < (2'h2)); forvar366 = (forvar366 + (1'h1)))
                begin
                  reg367 <= $unsigned((~^reg118[(3'h4):(3'h4)]));
                  for (forvar368 = (1'h0); (forvar368 < (2'h3)); forvar368 = (forvar368 + (1'h1)))
                    begin
                      reg369 <= $signed($signed($signed(reg271)));
                      reg370 <= reg45[(2'h2):(1'h1)];
                      reg371 <= $signed(($signed(((8'hb6) ?
                          reg254 : reg78)) <= (^~(^reg31))));
                    end
                  for (forvar372 = (1'h0); (forvar372 < (2'h2)); forvar372 = (forvar372 + (1'h1)))
                    begin
                      reg373 <= ({(reg361[(3'h6):(3'h6)] ?
                              (reg144 && reg21) : $unsigned((8'hb2)))} | {$unsigned(reg280[(3'h7):(2'h2)])});
                      reg374 <= (~^((reg94 ?
                          $unsigned(reg328) : ((8'h9c) ?
                              (8'hb6) : reg264)) != $unsigned((reg191 ?
                          reg135 : reg260))));
                    end
                end
              if ($signed(reg253[(4'h8):(3'h5)]))
                begin
                  if ((8'hb4))
                    begin
                      reg375 <= (reg328[(3'h5):(3'h5)] > $signed($signed(reg110)));
                      reg376 <= reg104;
                      reg377 <= $unsigned(($signed($signed(reg290)) && $unsigned($signed(reg373))));
                      reg378 <= $unsigned($signed({$signed(forvar315)}));
                    end
                  else
                    begin
                      reg375 <= $signed(wire174[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  if ((8'ha9))
                    begin
                      reg375 <= (wire10[(1'h0):(1'h0)] > $signed(($signed(reg276) ~^ (8'hb9))));
                      reg376 <= ($unsigned(reg97) ?
                          $unsigned($unsigned(reg113[(4'h9):(4'h8)])) : $unsigned((reg149[(1'h1):(1'h0)] ?
                              $signed(wire7) : {reg257})));
                      reg377 <= $signed({((8'ha0) < reg50)});
                      reg378 <= ({reg250[(2'h2):(1'h0)]} || ($signed((&(8'ha1))) ?
                          {reg208} : reg111[(3'h4):(1'h0)]));
                    end
                  else
                    begin
                      reg375 <= ($unsigned($signed((reg57 ?
                              reg75 : forvar368))) ?
                          reg259[(4'ha):(2'h2)] : reg77[(2'h2):(1'h0)]);
                      reg376 <= ((reg330[(2'h3):(2'h3)] ?
                          {$unsigned(reg261)} : (^(~&reg277))) & {reg42[(4'hb):(4'hb)]});
                      reg377 <= wire171;
                      reg378 <= ((~|$signed($unsigned(reg64))) ?
                          (&reg359[(2'h2):(1'h1)]) : $unsigned($signed({reg180})));
                    end
                  reg379 <= (^$unsigned((reg328 && $unsigned(reg193))));
                  for (forvar380 = (1'h0); (forvar380 < (1'h0)); forvar380 = (forvar380 + (1'h1)))
                    begin
                      reg381 <= ($signed(reg28[(2'h2):(1'h0)]) ?
                          (^~(reg83[(2'h2):(2'h2)] ?
                              (reg151 ?
                                  reg241 : reg294) : $signed(reg257))) : (|(8'ha9)));
                      reg382 <= reg245;
                      reg383 <= ($signed(((reg250 <= reg347) & (forvar325 ?
                              reg227 : reg19))) ?
                          ((((8'ha6) & reg314) + $signed(reg133)) ?
                              $unsigned(reg367[(1'h0):(1'h0)]) : {((8'ha8) << (8'hb8))}) : {reg264[(2'h2):(1'h1)]});
                    end
                end
              for (forvar384 = (1'h0); (forvar384 < (1'h1)); forvar384 = (forvar384 + (1'h1)))
                begin
                  reg385 <= (-$unsigned(({(8'ha8)} >>> (|reg310))));
                  reg386 <= (reg25 < (($signed(reg87) ?
                      (~^reg303) : reg377) || reg63));
                  for (forvar387 = (1'h0); (forvar387 < (2'h2)); forvar387 = (forvar387 + (1'h1)))
                    begin
                      reg388 <= $unsigned((~&{(&reg103)}));
                      reg389 <= ((~^reg364) >>> $unsigned({{reg321}}));
                      reg390 <= $unsigned(reg119[(3'h4):(3'h4)]);
                    end
                end
            end
        end
      else
        begin
          if (reg53)
            begin
              if (($signed(forvar304) ?
                  $signed(reg262[(3'h4):(2'h3)]) : ($unsigned({(8'haa)}) < reg382[(3'h7):(1'h0)])))
                begin
                  if ($signed((((~|reg367) ?
                      (&reg61) : reg116) << $signed($signed(reg272)))))
                    begin
                      reg304 <= ((^reg65) ?
                          {{{reg236}}} : ($signed(reg28) ?
                              reg299 : ($unsigned(reg374) || (reg240 ^~ reg313))));
                      reg305 <= $unsigned((~&reg95[(2'h3):(1'h0)]));
                      reg306 <= ((-$signed((forvar332 ? reg115 : reg21))) ?
                          $unsigned($unsigned((!forvar363))) : $unsigned(reg228[(4'h8):(2'h3)]));
                      reg307 <= $unsigned((reg302 ^ ((8'ha8) ?
                          reg369 : reg297)));
                    end
                  else
                    begin
                      reg304 <= forvar319;
                      reg305 <= (-(&$signed(reg206[(4'h9):(4'h8)])));
                      reg306 <= reg293;
                      reg307 <= $unsigned((~&reg85));
                    end
                  for (forvar308 = (1'h0); (forvar308 < (2'h2)); forvar308 = (forvar308 + (1'h1)))
                    begin
                      reg309 <= reg217;
                      reg310 <= reg285;
                    end
                  reg311 <= (($signed($signed((8'h9e))) == ((-reg337) <<< reg57)) ?
                      (($unsigned(reg122) ?
                          $unsigned(reg324) : $unsigned(reg85)) & $signed({(8'hb1)})) : (reg332[(4'hc):(3'h6)] ?
                          $signed(((8'hb5) || reg248)) : reg209));
                end
              else
                begin
                  for (forvar304 = (1'h0); (forvar304 < (2'h2)); forvar304 = (forvar304 + (1'h1)))
                    begin
                      reg305 <= {reg223};
                      reg306 <= $unsigned(((8'hb2) ?
                          (8'hae) : ((wire8 ? reg283 : reg150) < (reg336 ?
                              (8'hb9) : (8'hab)))));
                      reg307 <= $signed($signed((~^$unsigned(reg149))));
                    end
                end
              if ($unsigned((reg46[(2'h3):(1'h1)] ?
                  reg314 : $unsigned((^~reg61)))))
                begin
                  if (reg99)
                    begin
                      reg312 <= reg153;
                      reg313 <= reg303[(2'h2):(2'h2)];
                      reg314 <= $unsigned(reg356);
                    end
                  else
                    begin
                      reg312 <= $unsigned($unsigned(((!reg348) ?
                          (reg139 ^~ forvar345) : (reg129 ?
                              forvar325 : reg74))));
                      reg313 <= wire156[(3'h4):(2'h2)];
                    end
                  for (forvar315 = (1'h0); (forvar315 < (1'h1)); forvar315 = (forvar315 + (1'h1)))
                    begin
                      reg316 <= ($unsigned(($signed(reg306) ?
                              (reg206 ? reg20 : reg152) : $signed(reg220))) ?
                          $signed($signed(reg191)) : $signed(reg55));
                    end
                end
              else
                begin
                  if ((reg300 == reg95[(1'h0):(1'h0)]))
                    begin
                      reg312 <= $signed(forvar304);
                      reg313 <= (reg223[(1'h1):(1'h0)] ^~ (^$unsigned(((8'ha2) ^ reg75))));
                      reg314 <= $signed($unsigned(((reg276 ?
                          reg378 : reg98) <= {(8'had)})));
                    end
                  else
                    begin
                      reg312 <= (8'ha6);
                      reg313 <= ({(|$unsigned(forvar308))} * {reg106[(1'h1):(1'h0)]});
                      reg314 <= (wire8 - (~$signed((forvar345 < reg203))));
                    end
                  if (reg123[(3'h5):(2'h3)])
                    begin
                      reg315 <= {reg54};
                      reg316 <= ((reg264 ?
                              $unsigned($signed(reg212)) : $signed(forvar305[(2'h3):(2'h3)])) ?
                          reg152[(2'h3):(1'h0)] : ((&{reg334}) ?
                              reg21[(2'h3):(2'h2)] : {(reg290 != reg285)}));
                    end
                  else
                    begin
                      reg315 <= (^$signed((~^reg301)));
                      reg316 <= $unsigned(forvar305[(3'h7):(3'h4)]);
                      reg317 <= ((~&$signed(reg145)) ?
                          forvar308[(3'h5):(2'h3)] : $signed(($signed(reg123) ?
                              ((8'ha8) & wire11) : (reg276 < reg151))));
                    end
                  reg318 <= $signed(reg304);
                  if (reg251)
                    begin
                      reg319 <= $unsigned((8'ha4));
                      reg320 <= (~^(8'haf));
                      reg321 <= $signed((|forvar368[(3'h6):(1'h1)]));
                    end
                  else
                    begin
                      reg319 <= ($unsigned(reg319) ?
                          reg109 : (~|$unsigned(reg224[(2'h3):(1'h1)])));
                      reg320 <= ((8'h9c) >> (-((~|reg129) ?
                          (~&reg361) : $signed(reg284))));
                      reg321 <= ($signed((|$unsigned(reg213))) * reg302);
                    end
                end
            end
          else
            begin
              if (((+$signed($signed(reg34))) != $unsigned(reg334)))
                begin
                  if ({((|$unsigned((8'hb9))) ?
                          (reg124 ? (^reg266) : (~reg201)) : (8'had))})
                    begin
                      reg304 <= $unsigned(reg236[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg304 <= reg74;
                      reg305 <= ($unsigned((reg61[(3'h7):(2'h3)] ~^ (reg143 >= reg279))) >> (reg354 ?
                          (~|$unsigned(reg83)) : $signed((^~reg138))));
                      reg306 <= {({forvar368[(1'h0):(1'h0)]} & (reg114[(3'h5):(1'h0)] <= $unsigned(reg248)))};
                    end
                  for (forvar307 = (1'h0); (forvar307 < (2'h3)); forvar307 = (forvar307 + (1'h1)))
                    begin
                      reg308 <= $signed(reg353[(2'h2):(2'h2)]);
                      reg309 <= $unsigned(reg208[(3'h7):(3'h4)]);
                      reg310 <= ($unsigned(reg31[(4'h8):(1'h0)]) ?
                          reg284 : reg213);
                    end
                  for (forvar311 = (1'h0); (forvar311 < (1'h0)); forvar311 = (forvar311 + (1'h1)))
                    begin
                      reg312 <= ((reg65 != $unsigned((reg63 * forvar319))) ?
                          {$unsigned((+reg78))} : reg27[(3'h4):(1'h0)]);
                    end
                end
              else
                begin
                  if (reg266)
                    begin
                      reg304 <= (($signed({reg284}) > $unsigned($signed(reg145))) ~^ $signed((~^(~^(8'hb0)))));
                    end
                  else
                    begin
                      reg304 <= (|$unsigned((reg95 ^~ {reg316})));
                      reg305 <= reg81[(4'hb):(1'h1)];
                      reg306 <= $signed(($signed(reg328[(3'h7):(1'h1)]) ?
                          ((wire173 ? reg56 : reg284) ?
                              reg84 : (~|(8'hac))) : ((~^(8'hb9)) <<< $unsigned(reg146))));
                    end
                  reg307 <= (((~(8'hb9)) >> reg338) > reg256[(4'h8):(2'h3)]);
                  for (forvar308 = (1'h0); (forvar308 < (1'h1)); forvar308 = (forvar308 + (1'h1)))
                    begin
                      reg309 <= reg319[(1'h1):(1'h1)];
                    end
                end
              if (({$signed(reg106[(2'h2):(1'h1)])} << $unsigned(reg106[(1'h1):(1'h0)])))
                begin
                  for (forvar313 = (1'h0); (forvar313 < (2'h3)); forvar313 = (forvar313 + (1'h1)))
                    begin
                      reg314 <= {{((reg57 ^ reg371) ?
                                  reg197 : ((8'hb3) ~^ reg358))}};
                      reg315 <= (^~$signed((~^(8'hac))));
                      reg316 <= {reg112[(1'h0):(1'h0)]};
                    end
                  if ((~(+(!(!reg44)))))
                    begin
                      reg317 <= wire12[(1'h1):(1'h1)];
                      reg318 <= reg43;
                    end
                  else
                    begin
                      reg317 <= $signed(reg235[(1'h1):(1'h0)]);
                      reg318 <= $unsigned(reg369);
                      reg319 <= ((({reg24} ? (reg34 || (8'hba)) : (+reg371)) ?
                              reg309[(1'h1):(1'h0)] : $unsigned(reg123[(3'h5):(3'h4)])) ?
                          reg70[(1'h1):(1'h0)] : ($unsigned((^reg373)) ~^ ($signed(reg340) ?
                              $signed(reg310) : reg296[(3'h6):(2'h2)])));
                      reg320 <= reg98[(4'ha):(3'h7)];
                    end
                end
              else
                begin
                  if (((|reg17[(1'h1):(1'h0)]) | {{{reg82}}}))
                    begin
                      reg313 <= {reg182[(2'h3):(2'h2)]};
                      reg314 <= ((+(reg250[(1'h1):(1'h1)] ?
                              (reg292 ? forvar368 : reg340) : (^~reg316))) ?
                          (~&{{reg102}}) : ({reg195} ?
                              (reg19[(1'h0):(1'h0)] - $signed((8'hb1))) : reg55[(4'h9):(2'h3)]));
                    end
                  else
                    begin
                      reg313 <= (~&(^reg358[(4'hc):(4'ha)]));
                      reg314 <= ({$unsigned({reg276})} ?
                          reg99 : {(+(reg35 >> reg386))});
                    end
                  reg315 <= reg17[(2'h2):(1'h1)];
                  if ($unsigned(((^~(+(8'hb9))) | $signed(((8'h9d) ?
                      (8'had) : reg227)))))
                    begin
                      reg316 <= (~|(((reg206 ? reg314 : reg234) ?
                          ((8'ha0) ?
                              reg222 : (8'ha0)) : reg351[(1'h1):(1'h0)]) ^~ reg343[(2'h3):(1'h1)]));
                      reg317 <= ((reg34 ?
                          reg63[(1'h1):(1'h0)] : $unsigned(reg129)) == (((|(8'ha4)) ?
                              (reg53 ? reg338 : (8'hb8)) : (wire12 * wire173)) ?
                          $unsigned({reg316}) : $unsigned($signed((8'had)))));
                    end
                  else
                    begin
                      reg316 <= (((|(forvar380 ?
                              reg15 : forvar384)) ^~ reg317[(3'h4):(2'h2)]) ?
                          $signed((reg228[(4'h9):(3'h7)] ?
                              (~forvar368) : $unsigned(reg151))) : (^~reg75[(3'h6):(1'h1)]));
                      reg317 <= $unsigned(reg25[(2'h3):(2'h2)]);
                      reg318 <= (&(+reg386));
                      reg319 <= (|(|reg91[(1'h0):(1'h0)]));
                    end
                end
              for (forvar321 = (1'h0); (forvar321 < (1'h1)); forvar321 = (forvar321 + (1'h1)))
                begin
                  if ((reg56 + ((reg235[(2'h2):(2'h2)] ?
                          (|reg238) : $unsigned(reg300)) ?
                      $unsigned((~&(8'h9e))) : $unsigned(forvar324[(2'h3):(1'h1)]))))
                    begin
                      reg322 <= ($unsigned(((reg140 >= (8'hb9)) ?
                              (~reg62) : {reg374})) ?
                          (|$unsigned({reg82})) : (8'hba));
                      reg323 <= (reg136[(1'h1):(1'h1)] ?
                          reg273 : (reg25 && reg147));
                      reg324 <= reg309[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg322 <= (~$signed($unsigned(reg330)));
                      reg323 <= {(!$signed($unsigned((8'hae))))};
                      reg324 <= reg317;
                    end
                  for (forvar325 = (1'h0); (forvar325 < (1'h1)); forvar325 = (forvar325 + (1'h1)))
                    begin
                      reg326 <= reg342;
                      reg327 <= $signed(reg111[(2'h3):(2'h2)]);
                      reg328 <= ((~&$unsigned($signed(reg331))) ^ (reg30 == ($unsigned(reg243) + (forvar332 ?
                          reg311 : (8'ha9)))));
                      reg329 <= (-reg189[(2'h2):(2'h2)]);
                    end
                  for (forvar330 = (1'h0); (forvar330 < (2'h2)); forvar330 = (forvar330 + (1'h1)))
                    begin
                      reg331 <= reg226[(3'h4):(2'h3)];
                      reg332 <= reg47;
                      reg333 <= reg349[(1'h0):(1'h0)];
                      reg334 <= (~^reg214);
                    end
                  for (forvar335 = (1'h0); (forvar335 < (1'h1)); forvar335 = (forvar335 + (1'h1)))
                    begin
                      reg336 <= reg344;
                      reg337 <= $signed(($signed((^reg318)) & (reg338[(3'h6):(2'h2)] * {reg318})));
                    end
                end
              for (forvar338 = (1'h0); (forvar338 < (1'h1)); forvar338 = (forvar338 + (1'h1)))
                begin
                  for (forvar339 = (1'h0); (forvar339 < (2'h3)); forvar339 = (forvar339 + (1'h1)))
                    begin
                      reg340 <= reg374[(4'ha):(3'h4)];
                      reg341 <= (^~reg296[(1'h0):(1'h0)]);
                    end
                  reg342 <= (wire173 ?
                      reg33[(3'h5):(1'h1)] : reg201[(4'ha):(2'h2)]);
                end
            end
          reg343 <= $unsigned((+$unsigned((~reg294))));
          reg344 <= (~^$unsigned($signed($signed(reg148))));
          reg345 <= ((8'hb5) << ((~(-reg199)) ?
              {{reg385}} : ($unsigned(forvar345) ?
                  ((8'hb7) - (8'hb7)) : reg243)));
        end
      if (reg349)
        begin
          if ((~|reg226[(4'hb):(3'h5)]))
            begin
              for (forvar391 = (1'h0); (forvar391 < (2'h2)); forvar391 = (forvar391 + (1'h1)))
                begin
                  reg392 <= $unsigned((reg226 ?
                      $unsigned((~&reg334)) : reg23[(3'h5):(3'h4)]));
                end
            end
          else
            begin
              if ($signed(($unsigned(reg47) ?
                  $unsigned(((8'hb9) ? reg246 : reg82)) : reg35)))
                begin
                  reg391 <= reg201;
                  if ((&(~^((~&reg259) ? reg88 : (reg262 ? reg34 : reg81)))))
                    begin
                      reg392 <= $unsigned((8'h9d));
                      reg393 <= (|reg223);
                      reg394 <= (^~$unsigned(($unsigned(reg258) ?
                          $unsigned(reg302) : {reg255})));
                    end
                  else
                    begin
                      reg392 <= (reg185[(2'h2):(1'h1)] ?
                          {$signed((reg220 <= reg24))} : reg221);
                    end
                  for (forvar395 = (1'h0); (forvar395 < (1'h0)); forvar395 = (forvar395 + (1'h1)))
                    begin
                      reg396 <= $unsigned($unsigned((~&((8'ha6) ?
                          reg301 : forvar372))));
                      reg397 <= reg354[(2'h3):(2'h2)];
                      reg398 <= $unsigned((~&$unsigned(reg279)));
                      reg399 <= (((~reg253) <= ($unsigned((8'ha2)) >= (reg49 ?
                          reg331 : (8'ha6)))) ~^ $unsigned(reg314[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar391 = (1'h0); (forvar391 < (1'h1)); forvar391 = (forvar391 + (1'h1)))
                    begin
                      reg392 <= $signed((($unsigned((8'hac)) + (^~reg252)) ?
                          ((reg43 ?
                              reg136 : (8'ha9)) >>> (reg206 << (8'hab))) : reg92[(1'h0):(1'h0)]));
                      reg393 <= reg145;
                      reg394 <= reg253[(4'h9):(3'h7)];
                    end
                  for (forvar395 = (1'h0); (forvar395 < (2'h2)); forvar395 = (forvar395 + (1'h1)))
                    begin
                      reg396 <= ((-{$unsigned(reg108)}) < (8'h9c));
                      reg397 <= $unsigned(reg391);
                      reg398 <= (~|$signed($signed((reg55 ? reg28 : reg242))));
                    end
                end
            end
          for (forvar400 = (1'h0); (forvar400 < (2'h3)); forvar400 = (forvar400 + (1'h1)))
            begin
              if (((reg320[(1'h1):(1'h0)] > (8'ha0)) ^ (((reg148 - (8'hb1)) ?
                  $unsigned(reg317) : (reg292 >>> reg297)) == $signed((forvar332 > reg296)))))
                begin
                  for (forvar401 = (1'h0); (forvar401 < (2'h3)); forvar401 = (forvar401 + (1'h1)))
                    begin
                      reg402 <= $unsigned(($unsigned($signed(forvar319)) || $unsigned({reg122})));
                    end
                  if (($unsigned((|(reg55 + reg180))) ?
                      reg212 : $unsigned($unsigned((reg256 ? reg99 : reg388)))))
                    begin
                      reg403 <= (8'ha8);
                      reg404 <= ((!(!(reg93 ?
                          reg136 : reg326))) >> (reg203[(1'h0):(1'h0)] && ((+reg17) != (reg116 <= reg352))));
                      reg405 <= (-reg117[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg403 <= reg24[(1'h1):(1'h0)];
                    end
                  for (forvar406 = (1'h0); (forvar406 < (2'h3)); forvar406 = (forvar406 + (1'h1)))
                    begin
                      reg407 <= (^reg226);
                    end
                  reg408 <= (($unsigned(forvar335[(4'hd):(1'h1)]) ?
                      $unsigned(reg57) : (reg34 ?
                          (~|reg40) : reg109)) || $unsigned({(reg92 > (8'hb9))}));
                end
              else
                begin
                  reg401 <= $unsigned($signed(((forvar332 ?
                      reg377 : reg129) - ((8'hb0) == reg35))));
                  for (forvar402 = (1'h0); (forvar402 < (1'h0)); forvar402 = (forvar402 + (1'h1)))
                    begin
                      reg403 <= ($unsigned($unsigned($signed(reg292))) ?
                          (reg370 ?
                              ($unsigned(wire12) ?
                                  reg197 : ((8'hac) ?
                                      reg234 : (8'ha6))) : ((reg32 >= reg394) ?
                                  {reg313} : ((8'ha1) ?
                                      forvar349 : reg401))) : $signed((|reg85[(4'ha):(1'h0)])));
                      reg404 <= ($signed(reg327) ~^ $signed($signed((reg393 + reg189))));
                      reg405 <= reg305;
                      reg406 <= $unsigned(reg383[(4'hd):(4'ha)]);
                    end
                  reg407 <= $unsigned(reg327);
                end
              for (forvar409 = (1'h0); (forvar409 < (2'h3)); forvar409 = (forvar409 + (1'h1)))
                begin
                  reg410 <= (reg258[(1'h1):(1'h0)] ?
                      (~{$signed(reg100)}) : $unsigned((8'hb2)));
                  if ($unsigned((|(~reg25[(2'h2):(2'h2)]))))
                    begin
                      reg411 <= ({reg364} ?
                          (reg69 != reg208) : {(~&reg340[(2'h2):(1'h1)])});
                    end
                  else
                    begin
                      reg411 <= ({(reg279[(4'h8):(1'h0)] ?
                                  reg77[(4'h9):(2'h3)] : $signed(reg217))} ?
                          $unsigned(reg239) : $signed(({reg99} >> $unsigned((8'ha7)))));
                      reg412 <= $unsigned((8'ha4));
                    end
                  if (reg19)
                    begin
                      reg413 <= (({((8'haa) ? reg210 : reg240)} ?
                              reg240[(2'h2):(2'h2)] : $unsigned($unsigned(reg147))) ?
                          reg137 : $unsigned($unsigned($signed(reg300))));
                      reg414 <= $signed($signed(((-reg304) >>> (forvar409 ?
                          reg192 : reg313))));
                    end
                  else
                    begin
                      reg413 <= (forvar304 * reg283[(1'h0):(1'h0)]);
                      reg414 <= (forvar318 ?
                          (($signed((8'ha2)) >> $unsigned(reg413)) ?
                              reg213[(1'h1):(1'h1)] : (^reg302[(2'h2):(1'h1)])) : (reg95[(1'h1):(1'h0)] ?
                              reg118[(4'hb):(3'h5)] : {reg312}));
                      reg415 <= ($signed({reg338}) & {reg142});
                      reg416 <= $signed(forvar391);
                    end
                end
            end
          if (reg182)
            begin
              for (forvar417 = (1'h0); (forvar417 < (2'h2)); forvar417 = (forvar417 + (1'h1)))
                begin
                  reg418 <= reg403;
                end
            end
          else
            begin
              reg417 <= ((($unsigned(reg214) ?
                      ((8'h9e) ?
                          (8'hba) : reg129) : (reg370 && reg337)) - reg317) ?
                  (((^reg34) ?
                      $unsigned(reg222) : $signed(reg21)) * reg235) : $unsigned($unsigned((+reg85))));
              if ($signed($unsigned(reg111[(2'h2):(1'h0)])))
                begin
                  for (forvar418 = (1'h0); (forvar418 < (1'h1)); forvar418 = (forvar418 + (1'h1)))
                    begin
                      reg419 <= reg358;
                      reg420 <= $unsigned(($unsigned((forvar332 ?
                          forvar409 : reg150)) || $signed($signed(reg259))));
                    end
                  reg421 <= ((-(^(^~reg97))) & reg396);
                end
              else
                begin
                  reg418 <= (reg370[(4'he):(3'h6)] ?
                      (~^forvar335) : {((reg134 ? reg394 : reg197) ?
                              (reg248 ? forvar321 : reg49) : $signed(reg35))});
                end
            end
          if ({reg254})
            begin
              if (reg238[(2'h3):(1'h1)])
                begin
                  if ({reg72})
                    begin
                      reg422 <= $unsigned(wire155[(3'h4):(3'h4)]);
                      reg423 <= $unsigned((&reg382[(3'h7):(3'h7)]));
                    end
                  else
                    begin
                      reg422 <= reg336;
                      reg423 <= $signed((&{(forvar372 < reg290)}));
                    end
                  reg424 <= $unsigned((((-reg77) ?
                          $unsigned(forvar418) : reg33[(2'h2):(2'h2)]) ?
                      reg136 : wire173[(4'hc):(2'h2)]));
                  if ($signed(reg362))
                    begin
                      reg425 <= {($unsigned({reg388}) ?
                              $signed(reg46[(3'h4):(3'h4)]) : (forvar349 ?
                                  reg398 : $unsigned(reg21)))};
                      reg426 <= {(((reg93 >= (8'ha6)) ?
                              (+reg330) : $unsigned(reg389)) ^~ reg64[(3'h4):(2'h2)])};
                      reg427 <= $unsigned(reg93);
                    end
                  else
                    begin
                      reg425 <= (~|(((reg84 ? reg422 : (8'haf)) ?
                          forvar305 : $signed((8'ha6))) && $unsigned((^reg280))));
                    end
                  reg428 <= {$unsigned($signed(reg263))};
                end
              else
                begin
                  for (forvar422 = (1'h0); (forvar422 < (1'h1)); forvar422 = (forvar422 + (1'h1)))
                    begin
                      reg423 <= forvar313[(1'h0):(1'h0)];
                      reg424 <= {$unsigned($unsigned(reg108[(3'h7):(3'h5)]))};
                    end
                  if ($unsigned($signed($unsigned((reg23 ? reg86 : reg280)))))
                    begin
                      reg425 <= ($unsigned((~((8'hb8) & (8'ha6)))) - $signed((~^(reg56 ?
                          (8'hab) : (8'hb2)))));
                      reg426 <= forvar324[(1'h1):(1'h0)];
                      reg427 <= $unsigned(($unsigned((reg212 | forvar325)) ?
                          $unsigned($unsigned(reg245)) : ((reg108 ^~ reg55) || $signed(reg129))));
                    end
                  else
                    begin
                      reg425 <= $unsigned(reg135[(4'h8):(1'h1)]);
                      reg426 <= $signed({$unsigned({(8'ha0)})});
                      reg427 <= reg335[(3'h5):(3'h5)];
                    end
                  for (forvar428 = (1'h0); (forvar428 < (1'h1)); forvar428 = (forvar428 + (1'h1)))
                    begin
                      reg429 <= $unsigned((reg311[(1'h0):(1'h0)] ?
                          $signed(forvar418) : reg261));
                    end
                end
              reg430 <= $unsigned(((~&(reg193 ? reg29 : reg145)) ?
                  $unsigned((reg27 <<< wire11)) : (8'ha5)));
            end
          else
            begin
              for (forvar422 = (1'h0); (forvar422 < (1'h1)); forvar422 = (forvar422 + (1'h1)))
                begin
                  reg423 <= (-reg264);
                end
              if ((-({(reg277 != reg250)} != (reg304[(3'h4):(3'h4)] ?
                  (forvar324 <= reg390) : (reg20 >= reg403)))))
                begin
                  for (forvar424 = (1'h0); (forvar424 < (1'h0)); forvar424 = (forvar424 + (1'h1)))
                    begin
                      reg425 <= {$signed({(reg359 ? (8'ha5) : reg47)})};
                      reg426 <= $unsigned(reg88);
                      reg427 <= (~|($signed($unsigned(reg93)) ^~ reg389));
                      reg428 <= forvar304[(3'h7):(2'h3)];
                    end
                  reg429 <= (~^(($signed((8'hb3)) ?
                      (~^reg21) : $unsigned(reg378)) > ((reg16 ?
                      (8'ha2) : forvar387) ^ (8'h9d))));
                end
              else
                begin
                  for (forvar424 = (1'h0); (forvar424 < (1'h0)); forvar424 = (forvar424 + (1'h1)))
                    begin
                      reg425 <= reg376[(4'h8):(3'h5)];
                      reg426 <= $unsigned($unsigned(reg271[(2'h2):(1'h0)]));
                      reg427 <= (8'ha1);
                    end
                  if (forvar309)
                    begin
                      reg428 <= reg332[(3'h6):(1'h0)];
                      reg429 <= (8'hb0);
                    end
                  else
                    begin
                      reg428 <= (~|($unsigned($signed(reg374)) ?
                          ({forvar311} | reg293) : $signed(((8'hb1) ?
                              reg63 : reg252))));
                      reg429 <= {{((reg343 ^ reg69) <<< reg133)}};
                      reg430 <= {$signed(((|(8'hb0)) & forvar342))};
                      reg431 <= reg358[(3'h6):(2'h3)];
                    end
                end
            end
        end
      else
        begin
          reg391 <= (~|(^{{reg49}}));
          reg392 <= ($signed($signed((~|reg63))) == forvar409);
          if ($signed(reg43))
            begin
              for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
                begin
                  if (reg329[(1'h1):(1'h0)])
                    begin
                      reg394 <= $signed(reg330[(3'h5):(2'h3)]);
                      reg395 <= $unsigned(reg253[(3'h5):(1'h1)]);
                      reg396 <= (((reg94[(3'h7):(3'h4)] ^ (^reg143)) ?
                              wire8 : (reg134[(2'h3):(2'h2)] - reg272[(2'h2):(2'h2)])) ?
                          $unsigned((|reg136[(1'h1):(1'h0)])) : reg423[(4'h8):(2'h3)]);
                    end
                  else
                    begin
                      reg394 <= {$signed((^(reg377 ? reg42 : reg276)))};
                      reg395 <= $signed(reg91);
                    end
                  for (forvar397 = (1'h0); (forvar397 < (1'h0)); forvar397 = (forvar397 + (1'h1)))
                    begin
                      reg398 <= ((~|$signed((reg75 >>> reg369))) ~^ $signed(((8'h9f) ?
                          reg22[(3'h4):(2'h3)] : reg144)));
                    end
                  reg399 <= (reg280 ? reg30[(4'h9):(3'h5)] : (|reg110));
                end
            end
          else
            begin
              if ($unsigned($unsigned((^~reg198))))
                begin
                  if (reg272)
                    begin
                      reg393 <= reg394[(3'h5):(2'h2)];
                      reg394 <= {(reg344 <= $signed((forvar349 ?
                              reg81 : reg397)))};
                      reg395 <= reg187[(2'h3):(1'h1)];
                      reg396 <= $unsigned(reg140[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg393 <= (|reg408);
                      reg394 <= reg72;
                      reg395 <= reg25;
                    end
                end
              else
                begin
                  reg393 <= reg97[(3'h4):(1'h0)];
                  for (forvar394 = (1'h0); (forvar394 < (2'h3)); forvar394 = (forvar394 + (1'h1)))
                    begin
                      reg395 <= $unsigned(reg242);
                      reg396 <= (^(-forvar387));
                    end
                  if ((+($signed({reg365}) | (~(forvar335 ?
                      wire173 : reg414)))))
                    begin
                      reg397 <= reg99[(1'h1):(1'h0)];
                      reg398 <= ((($unsigned(reg244) ?
                                  $unsigned(reg210) : reg133[(2'h3):(1'h1)]) ?
                              ($signed(reg252) ?
                                  (forvar335 == reg208) : {reg414}) : ((reg16 >= reg414) & (8'ha9))) ?
                          $unsigned((reg390[(1'h1):(1'h1)] ?
                              (8'ha9) : $signed(reg216))) : $signed(forvar332));
                      reg399 <= reg238;
                      reg400 <= {reg100};
                    end
                  else
                    begin
                      reg397 <= (~&$unsigned(((^~reg365) == $unsigned(forvar391))));
                      reg398 <= (+$unsigned(reg86[(1'h1):(1'h1)]));
                      reg399 <= (^(+((reg108 ? reg382 : reg249) ?
                          $unsigned(forvar394) : reg365)));
                    end
                end
              for (forvar401 = (1'h0); (forvar401 < (1'h1)); forvar401 = (forvar401 + (1'h1)))
                begin
                  for (forvar402 = (1'h0); (forvar402 < (1'h1)); forvar402 = (forvar402 + (1'h1)))
                    begin
                      reg403 <= reg262;
                      reg404 <= (!wire156);
                      reg405 <= $unsigned($signed(reg15[(3'h4):(3'h4)]));
                      reg406 <= (($signed($unsigned(reg307)) ?
                              $unsigned(reg149) : (reg314[(1'h0):(1'h0)] & (forvar332 * (8'hac)))) ?
                          reg400 : reg259);
                    end
                  for (forvar407 = (1'h0); (forvar407 < (1'h0)); forvar407 = (forvar407 + (1'h1)))
                    begin
                      reg408 <= reg389;
                      reg409 <= (reg109[(2'h3):(1'h1)] || reg101[(3'h4):(2'h3)]);
                    end
                  for (forvar410 = (1'h0); (forvar410 < (1'h1)); forvar410 = (forvar410 + (1'h1)))
                    begin
                      reg411 <= (|$unsigned(reg362));
                      reg412 <= $unsigned(({(~^reg360)} ?
                          {(~^forvar332)} : reg264[(4'hc):(4'hc)]));
                    end
                end
              for (forvar413 = (1'h0); (forvar413 < (1'h0)); forvar413 = (forvar413 + (1'h1)))
                begin
                  reg414 <= (&(8'hae));
                  for (forvar415 = (1'h0); (forvar415 < (1'h1)); forvar415 = (forvar415 + (1'h1)))
                    begin
                      reg416 <= (+reg294);
                    end
                end
              reg417 <= (&(forvar368 ?
                  {$signed(reg33)} : ($unsigned(reg315) ?
                      $signed(reg313) : (&reg338))));
            end
        end
      for (forvar432 = (1'h0); (forvar432 < (1'h1)); forvar432 = (forvar432 + (1'h1)))
        begin
          for (forvar433 = (1'h0); (forvar433 < (2'h3)); forvar433 = (forvar433 + (1'h1)))
            begin
              for (forvar434 = (1'h0); (forvar434 < (1'h1)); forvar434 = (forvar434 + (1'h1)))
                begin
                  for (forvar435 = (1'h0); (forvar435 < (1'h0)); forvar435 = (forvar435 + (1'h1)))
                    begin
                      reg436 <= $signed($unsigned({$unsigned(reg100)}));
                      reg437 <= (|$unsigned($signed(reg337[(3'h6):(3'h6)])));
                      reg438 <= (reg391[(3'h4):(3'h4)] ?
                          $signed({((8'ha9) >>> reg113)}) : reg419);
                      reg439 <= reg308[(3'h7):(3'h6)];
                    end
                  reg440 <= (reg279[(1'h1):(1'h0)] ?
                      $unsigned({(~|reg80)}) : reg71);
                end
              for (forvar441 = (1'h0); (forvar441 < (2'h2)); forvar441 = (forvar441 + (1'h1)))
                begin
                  reg442 <= (^~$signed(reg223));
                  for (forvar443 = (1'h0); (forvar443 < (1'h0)); forvar443 = (forvar443 + (1'h1)))
                    begin
                      reg444 <= ((~&forvar342) << reg252);
                    end
                  reg445 <= ($signed(reg345[(4'h8):(2'h2)]) ?
                      $unsigned((reg261[(2'h3):(2'h3)] ?
                          ((8'hac) ?
                              reg33 : reg270) : wire7)) : ($signed((~|reg49)) >= forvar342));
                end
              reg446 <= {$signed($unsigned(reg390))};
            end
        end
    end
  assign wire447 = $unsigned($unsigned(({reg421} ?
                       reg354 : (reg355 == reg149))));
  always
    @(posedge clk) begin
      for (forvar448 = (1'h0); (forvar448 < (2'h3)); forvar448 = (forvar448 + (1'h1)))
        begin
          if ({reg38[(3'h7):(3'h7)]})
            begin
              if (reg374)
                begin
                  for (forvar449 = (1'h0); (forvar449 < (1'h1)); forvar449 = (forvar449 + (1'h1)))
                    begin
                      reg450 <= ((^~{reg122[(1'h0):(1'h0)]}) ?
                          reg232 : reg217[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  if ((8'hb4))
                    begin
                      reg449 <= reg290;
                      reg450 <= reg322[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg449 <= (~|{$unsigned(reg145[(2'h2):(2'h2)])});
                    end
                  reg451 <= wire174[(1'h1):(1'h0)];
                end
              if ($unsigned($unsigned((reg311 | ((8'hb0) ? reg137 : reg334)))))
                begin
                  reg452 <= reg374;
                  if (reg358)
                    begin
                      reg453 <= $signed(($signed((-(8'ha9))) > ({(8'h9d)} ?
                          (reg182 ? reg183 : reg371) : reg260)));
                      reg454 <= (!$signed($signed((^reg223))));
                    end
                  else
                    begin
                      reg453 <= {(reg136[(2'h2):(1'h0)] | reg111)};
                      reg454 <= $signed($signed($unsigned($unsigned(reg416))));
                    end
                end
              else
                begin
                  for (forvar452 = (1'h0); (forvar452 < (2'h2)); forvar452 = (forvar452 + (1'h1)))
                    begin
                      reg453 <= ($signed(reg276[(2'h2):(1'h1)]) ?
                          ((((8'hb1) <<< reg261) != (reg388 ? reg40 : reg201)) ?
                              ($unsigned(reg431) ?
                                  {reg210} : $signed((8'hb7))) : {reg337[(3'h6):(3'h4)]}) : reg50);
                      reg454 <= reg329[(3'h4):(2'h2)];
                    end
                  if ($signed(((&reg323) ~^ (reg261 ?
                      ((8'hb0) ? reg56 : reg226) : (~^reg350)))))
                    begin
                      reg455 <= (reg408[(4'hd):(2'h3)] ?
                          $unsigned(reg154[(1'h0):(1'h0)]) : ((~|reg122) ?
                              (^$signed((8'ha6))) : {wire447[(3'h5):(2'h2)]}));
                      reg456 <= reg240[(2'h3):(1'h1)];
                      reg457 <= $signed((+(reg352[(3'h4):(2'h3)] << (!wire9))));
                      reg458 <= $unsigned($unsigned($signed(reg403[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg455 <= wire174;
                      reg456 <= $signed($unsigned(reg424[(1'h0):(1'h0)]));
                    end
                  if (reg20)
                    begin
                      reg459 <= ($unsigned(reg403) ?
                          (~|((reg43 ? reg438 : reg246) ?
                              (|reg427) : reg224[(1'h0):(1'h0)])) : reg94);
                    end
                  else
                    begin
                      reg459 <= $signed(reg424[(1'h1):(1'h1)]);
                      reg460 <= reg361;
                    end
                  reg461 <= $signed((((wire9 ? reg180 : (8'h9e)) & ((8'h9d) ?
                          reg137 : reg239)) ?
                      (((8'haa) ? reg221 : reg323) ^ {reg239}) : (!(reg249 ?
                          reg409 : reg21))));
                end
              if ($signed((reg258[(2'h3):(2'h3)] ?
                  reg256 : $unsigned($signed(reg256)))))
                begin
                  if (reg73[(2'h2):(1'h0)])
                    begin
                      reg462 <= $unsigned($unsigned(((reg319 >> reg34) && $unsigned(reg329))));
                      reg463 <= $unsigned($unsigned(($unsigned(reg354) ?
                          $unsigned(wire8) : $signed(reg228))));
                      reg464 <= $signed((^~$signed($unsigned(reg300))));
                      reg465 <= reg99[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg462 <= $unsigned(reg24[(2'h2):(1'h0)]);
                      reg463 <= $unsigned($unsigned((+(^reg368))));
                      reg464 <= $unsigned($unsigned(reg399[(1'h0):(1'h0)]));
                      reg465 <= (($unsigned(reg333) || reg312[(3'h5):(1'h1)]) ^ $signed($signed(reg376[(3'h5):(2'h3)])));
                    end
                end
              else
                begin
                  if ($signed((!(|$unsigned(reg365)))))
                    begin
                      reg462 <= ({$signed(reg428)} | {$signed(reg245[(2'h2):(2'h2)])});
                    end
                  else
                    begin
                      reg462 <= $signed(((~(!reg460)) <<< (reg331[(3'h5):(2'h3)] ~^ ((8'hb5) ?
                          reg74 : reg74))));
                    end
                  for (forvar463 = (1'h0); (forvar463 < (1'h0)); forvar463 = (forvar463 + (1'h1)))
                    begin
                      reg464 <= reg379;
                    end
                  if ($signed((((reg360 ? reg305 : reg241) ?
                      (+reg226) : reg238[(3'h5):(1'h0)]) ^~ $signed((~|(8'hba))))))
                    begin
                      reg465 <= reg197;
                      reg466 <= ((!((~reg221) <<< reg148[(3'h5):(1'h1)])) >> reg392);
                      reg467 <= ((!{((8'h9f) | (8'ha8))}) ?
                          ({reg64[(2'h3):(2'h3)]} <= reg271) : reg393);
                    end
                  else
                    begin
                      reg465 <= {reg264[(1'h1):(1'h0)]};
                      reg466 <= reg296[(3'h4):(1'h1)];
                      reg467 <= (&(reg191[(4'h8):(2'h2)] ?
                          $signed(reg259) : ((+reg80) ? reg328 : {reg412})));
                      reg468 <= (~^(((reg277 ? reg195 : reg227) ~^ (^~reg233)) ?
                          reg456 : (8'hb0)));
                    end
                end
              reg469 <= reg307;
            end
          else
            begin
              for (forvar449 = (1'h0); (forvar449 < (2'h2)); forvar449 = (forvar449 + (1'h1)))
                begin
                  reg450 <= {(&$unsigned((-(8'hae))))};
                  if ($unsigned(reg290[(2'h2):(2'h2)]))
                    begin
                      reg451 <= $signed($unsigned($signed((reg116 ?
                          reg410 : reg46))));
                      reg452 <= (~&reg403);
                      reg453 <= $unsigned((|($unsigned(reg337) * reg308)));
                    end
                  else
                    begin
                      reg451 <= $unsigned($unsigned($signed(reg110)));
                    end
                end
              reg454 <= $signed(forvar463);
            end
          if ($unsigned($signed($unsigned((reg273 ? reg389 : reg437)))))
            begin
              if (reg241)
                begin
                  for (forvar470 = (1'h0); (forvar470 < (1'h1)); forvar470 = (forvar470 + (1'h1)))
                    begin
                      reg471 <= $signed($unsigned((reg294[(1'h0):(1'h0)] ?
                          (!reg100) : (reg192 ? (8'hb5) : reg393))));
                    end
                end
              else
                begin
                  if ($signed((8'hae)))
                    begin
                      reg470 <= $unsigned($unsigned($signed((8'hb5))));
                      reg471 <= wire7[(1'h0):(1'h0)];
                      reg472 <= (|(|(+reg85[(3'h7):(3'h4)])));
                      reg473 <= (($signed((reg383 | (8'ha9))) ?
                          (reg54 ^~ (reg341 ?
                              reg56 : reg414)) : $signed(reg191)) - $unsigned((~|reg247[(4'hf):(2'h2)])));
                    end
                  else
                    begin
                      reg470 <= $unsigned((&$signed(reg209[(1'h0):(1'h0)])));
                    end
                end
            end
          else
            begin
              for (forvar470 = (1'h0); (forvar470 < (2'h3)); forvar470 = (forvar470 + (1'h1)))
                begin
                  if ({reg377})
                    begin
                      reg471 <= ((reg21 ^ reg91[(1'h1):(1'h0)]) >>> (($signed(reg284) | reg453[(4'h9):(4'h9)]) ?
                          (reg53[(2'h3):(2'h3)] ?
                              (reg88 | reg71) : reg416) : $signed(((8'hb5) >> reg298))));
                      reg472 <= (~^((8'ha9) <<< (~&(wire12 | reg417))));
                    end
                  else
                    begin
                      reg471 <= $signed(($unsigned({reg178}) == (reg20[(1'h0):(1'h0)] ?
                          (reg427 < (8'hba)) : reg370[(4'hd):(4'hd)])));
                      reg472 <= ((!{$unsigned(reg382)}) ?
                          ((reg469 == $signed(reg227)) ?
                              (reg80[(1'h1):(1'h0)] * $unsigned(reg36)) : reg82) : (($signed(reg254) ?
                              (reg208 ?
                                  reg105 : (8'ha2)) : (reg413 + reg331)) >> reg450));
                      reg473 <= ($unsigned({reg198[(3'h4):(2'h3)]}) < ($signed($signed(wire156)) ^~ ((reg426 || reg217) >>> $signed(reg116))));
                    end
                end
            end
        end
      for (forvar474 = (1'h0); (forvar474 < (2'h2)); forvar474 = (forvar474 + (1'h1)))
        begin
          for (forvar475 = (1'h0); (forvar475 < (2'h2)); forvar475 = (forvar475 + (1'h1)))
            begin
              if ((+reg371))
                begin
                  for (forvar476 = (1'h0); (forvar476 < (2'h3)); forvar476 = (forvar476 + (1'h1)))
                    begin
                      reg477 <= ((reg222 != $unsigned(reg197[(3'h7):(3'h5)])) ?
                          ({reg317} ?
                              {(8'hb9)} : {(forvar449 ?
                                      reg249 : reg279)}) : (({reg80} < reg338[(1'h1):(1'h1)]) < (reg223 == ((8'hab) == reg94))));
                      reg478 <= (((&(reg103 ? reg457 : reg19)) | reg358) ?
                          {((reg289 <= reg244) < (reg209 || reg52))} : {$unsigned($unsigned(reg134))});
                      reg479 <= reg75;
                    end
                end
              else
                begin
                  for (forvar476 = (1'h0); (forvar476 < (2'h2)); forvar476 = (forvar476 + (1'h1)))
                    begin
                      reg477 <= (~^reg122[(3'h4):(1'h1)]);
                    end
                  for (forvar478 = (1'h0); (forvar478 < (2'h2)); forvar478 = (forvar478 + (1'h1)))
                    begin
                      reg479 <= $unsigned(($signed(reg135) ?
                          $unsigned($signed(reg381)) : ($signed(reg218) * (~&reg208))));
                      reg480 <= (((8'hab) || {reg183[(2'h3):(2'h3)]}) * (reg299[(4'hd):(3'h6)] ?
                          ($signed((8'hb7)) && (reg234 <= reg439)) : ($unsigned(reg479) * (!reg37))));
                    end
                end
              if ((reg406[(1'h0):(1'h0)] ?
                  reg305 : $unsigned($unsigned((reg275 ? reg307 : reg236)))))
                begin
                  for (forvar481 = (1'h0); (forvar481 < (2'h2)); forvar481 = (forvar481 + (1'h1)))
                    begin
                      reg482 <= reg43[(4'hc):(3'h7)];
                    end
                  if ((8'h9e))
                    begin
                      reg483 <= reg37;
                      reg484 <= (^~(~^($unsigned(reg98) ?
                          (reg281 ? (8'hb7) : reg242) : (~reg305))));
                      reg485 <= reg467;
                      reg486 <= reg379;
                    end
                  else
                    begin
                      reg483 <= $unsigned((!((&reg188) ?
                          (-reg140) : $signed((8'ha9)))));
                    end
                  reg487 <= reg341;
                  if (($unsigned($signed(reg320)) && $unsigned((^(reg463 ^~ reg185)))))
                    begin
                      reg488 <= ($unsigned((8'hba)) ~^ (~|($signed(reg264) ?
                          (reg396 >> reg479) : $unsigned(reg412))));
                      reg489 <= (8'ha1);
                      reg490 <= {$signed($unsigned($signed(reg480)))};
                    end
                  else
                    begin
                      reg488 <= (($signed($unsigned(reg224)) ?
                              reg185 : $signed((reg488 ? (8'hb0) : reg260))) ?
                          {(~$unsigned(reg299))} : $unsigned(reg148));
                    end
                end
              else
                begin
                  reg481 <= reg449;
                end
              reg491 <= {{($signed(reg454) ?
                          {(8'h9c)} : reg206[(1'h0):(1'h0)])}};
            end
          if (({$unsigned((+reg201))} ?
              $signed($signed((^~reg491))) : (&reg36)))
            begin
              for (forvar492 = (1'h0); (forvar492 < (2'h2)); forvar492 = (forvar492 + (1'h1)))
                begin
                  reg493 <= {(!$signed($signed(reg260)))};
                end
            end
          else
            begin
              for (forvar492 = (1'h0); (forvar492 < (2'h3)); forvar492 = (forvar492 + (1'h1)))
                begin
                  for (forvar493 = (1'h0); (forvar493 < (1'h0)); forvar493 = (forvar493 + (1'h1)))
                    begin
                      reg494 <= (reg145[(1'h1):(1'h0)] ?
                          reg358 : $unsigned(((8'ha6) ?
                              $unsigned(reg100) : reg83[(1'h1):(1'h0)])));
                      reg495 <= $unsigned($signed(reg316));
                      reg496 <= reg275[(2'h2):(1'h1)];
                    end
                  if ($unsigned(($signed(reg134) ? reg74 : (^~{(8'had)}))))
                    begin
                      reg497 <= (!(~|reg446));
                    end
                  else
                    begin
                      reg497 <= (|$signed($signed((reg349 || reg105))));
                      reg498 <= wire13;
                    end
                end
              if (reg285)
                begin
                  if ({(reg362 ? {$signed(reg345)} : (&reg428[(3'h7):(3'h6)]))})
                    begin
                      reg499 <= $unsigned($unsigned($unsigned((~^reg410))));
                      reg500 <= {$signed($unsigned((+reg357)))};
                      reg501 <= ((reg28[(4'hd):(4'hd)] ^~ reg100) ^~ reg27);
                      reg502 <= $signed(reg23);
                    end
                  else
                    begin
                      reg499 <= reg415;
                      reg500 <= {reg297};
                    end
                  for (forvar503 = (1'h0); (forvar503 < (2'h3)); forvar503 = (forvar503 + (1'h1)))
                    begin
                      reg504 <= reg410[(2'h2):(1'h1)];
                    end
                  if ((reg199[(1'h0):(1'h0)] ?
                      (reg317[(4'h8):(3'h6)] ?
                          $signed($signed(reg25)) : reg221[(3'h6):(2'h3)]) : reg440))
                    begin
                      reg505 <= (-reg409);
                      reg506 <= {(|$unsigned(reg61[(2'h3):(2'h3)]))};
                    end
                  else
                    begin
                      reg505 <= reg232;
                      reg506 <= (($signed((~|reg222)) ?
                          reg364 : ((reg299 > (8'hb2)) >>> (reg44 - reg73))) + $unsigned((~{reg142})));
                      reg507 <= reg401[(2'h2):(2'h2)];
                      reg508 <= {reg216};
                    end
                end
              else
                begin
                  reg499 <= ($signed(forvar448[(2'h3):(2'h3)]) >>> ({$unsigned(reg100)} - ((reg426 > reg450) ?
                      reg70 : {reg338})));
                  for (forvar500 = (1'h0); (forvar500 < (1'h1)); forvar500 = (forvar500 + (1'h1)))
                    begin
                      reg501 <= reg390;
                      reg502 <= $signed((({reg305} - reg377[(1'h0):(1'h0)]) ?
                          reg465 : $unsigned({reg446})));
                      reg503 <= $signed((&reg449));
                      reg504 <= (8'ha4);
                    end
                  if (($unsigned($unsigned({(8'hba)})) ?
                      forvar500[(1'h0):(1'h0)] : {$unsigned($unsigned(reg281))}))
                    begin
                      reg505 <= (~|((~|(~reg421)) ?
                          reg327 : $signed((reg344 == reg427))));
                      reg506 <= reg32;
                    end
                  else
                    begin
                      reg505 <= $signed(reg285[(3'h4):(2'h2)]);
                    end
                end
              for (forvar509 = (1'h0); (forvar509 < (1'h1)); forvar509 = (forvar509 + (1'h1)))
                begin
                  if ((~|($unsigned($signed(reg223)) ?
                      (~|reg55) : {(~&reg312)})))
                    begin
                      reg510 <= $signed((8'hb2));
                      reg511 <= (+($signed($unsigned(reg30)) < $signed((reg151 * reg411))));
                    end
                  else
                    begin
                      reg510 <= (reg105 ?
                          {reg394} : ($signed((~&reg35)) <<< {(&reg23)}));
                      reg511 <= $unsigned({($signed(reg71) * $unsigned(reg500))});
                      reg512 <= (($unsigned(reg285) ?
                          $signed(reg507) : (8'hab)) == $unsigned($unsigned($unsigned(reg379))));
                    end
                  if ((~&reg326))
                    begin
                      reg513 <= $unsigned(({reg452[(2'h3):(1'h0)]} >= ($signed((8'ha2)) ?
                          (^~reg450) : {reg488})));
                      reg514 <= reg513;
                    end
                  else
                    begin
                      reg513 <= (reg256[(3'h4):(1'h1)] | $signed(reg430[(2'h3):(1'h1)]));
                    end
                  if ($signed(reg396))
                    begin
                      reg515 <= $unsigned(reg378[(2'h3):(1'h1)]);
                      reg516 <= (+$unsigned(reg341));
                      reg517 <= reg494;
                    end
                  else
                    begin
                      reg515 <= ($unsigned((^reg392)) <= $unsigned(({(8'hb0)} + reg438[(3'h4):(2'h3)])));
                    end
                  for (forvar518 = (1'h0); (forvar518 < (2'h3)); forvar518 = (forvar518 + (1'h1)))
                    begin
                      reg519 <= wire447;
                    end
                end
              reg520 <= $unsigned($unsigned((+(reg477 | reg355))));
            end
          if ($unsigned((($unsigned(reg241) <= reg412[(4'h9):(3'h4)]) >= $unsigned($signed(reg220)))))
            begin
              for (forvar521 = (1'h0); (forvar521 < (1'h1)); forvar521 = (forvar521 + (1'h1)))
                begin
                  for (forvar522 = (1'h0); (forvar522 < (1'h1)); forvar522 = (forvar522 + (1'h1)))
                    begin
                      reg523 <= reg120[(1'h0):(1'h0)];
                    end
                  if (reg104)
                    begin
                      reg524 <= $signed(reg272[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg524 <= {((reg490 ?
                              (~|reg361) : forvar492[(4'h9):(3'h5)]) | $signed((reg311 + reg259)))};
                      reg525 <= (!$unsigned($unsigned((reg512 < reg356))));
                      reg526 <= $signed($unsigned(reg496[(4'hb):(3'h5)]));
                      reg527 <= {reg123[(3'h5):(1'h0)]};
                    end
                  for (forvar528 = (1'h0); (forvar528 < (1'h1)); forvar528 = (forvar528 + (1'h1)))
                    begin
                      reg529 <= wire9;
                      reg530 <= (~|(reg216[(1'h0):(1'h0)] ? reg63 : reg417));
                    end
                  reg531 <= reg316[(3'h5):(3'h5)];
                end
              for (forvar532 = (1'h0); (forvar532 < (1'h1)); forvar532 = (forvar532 + (1'h1)))
                begin
                  if ($unsigned(reg424))
                    begin
                      reg533 <= (reg346[(2'h3):(1'h0)] < (reg365 ?
                          $unsigned((reg125 >>> reg29)) : reg135));
                      reg534 <= reg33;
                      reg535 <= ((-(8'ha5)) >>> (~|$signed(((8'hb5) ?
                          (8'hb6) : (8'hb4)))));
                    end
                  else
                    begin
                      reg533 <= $signed(reg481);
                      reg534 <= $signed((&$unsigned((8'h9c))));
                    end
                  for (forvar536 = (1'h0); (forvar536 < (2'h2)); forvar536 = (forvar536 + (1'h1)))
                    begin
                      reg537 <= $signed((reg506 || $signed(reg242)));
                    end
                end
              reg538 <= $signed(reg70);
            end
          else
            begin
              for (forvar521 = (1'h0); (forvar521 < (2'h3)); forvar521 = (forvar521 + (1'h1)))
                begin
                  for (forvar522 = (1'h0); (forvar522 < (1'h0)); forvar522 = (forvar522 + (1'h1)))
                    begin
                      reg523 <= reg134;
                      reg524 <= reg305[(4'h9):(2'h2)];
                      reg525 <= (^$signed(((reg377 < (8'hab)) && (8'h9d))));
                    end
                  for (forvar526 = (1'h0); (forvar526 < (2'h2)); forvar526 = (forvar526 + (1'h1)))
                    begin
                      reg527 <= ($signed(reg373[(1'h1):(1'h1)]) <= {{(reg261 >> reg538)}});
                      reg528 <= $unsigned(reg523[(3'h4):(3'h4)]);
                      reg529 <= (8'hb5);
                      reg530 <= $signed(reg324[(2'h3):(1'h0)]);
                    end
                end
              reg531 <= reg494[(1'h0):(1'h0)];
            end
          reg539 <= reg386;
        end
      for (forvar540 = (1'h0); (forvar540 < (2'h2)); forvar540 = (forvar540 + (1'h1)))
        begin
          for (forvar541 = (1'h0); (forvar541 < (2'h2)); forvar541 = (forvar541 + (1'h1)))
            begin
              reg542 <= reg333;
              for (forvar543 = (1'h0); (forvar543 < (1'h0)); forvar543 = (forvar543 + (1'h1)))
                begin
                  if (reg135[(3'h5):(2'h3)])
                    begin
                      reg544 <= (reg400[(4'h9):(3'h5)] ?
                          $unsigned(($signed(reg234) < reg130[(1'h0):(1'h0)])) : (^~(8'hb8)));
                      reg545 <= {reg188[(1'h0):(1'h0)]};
                      reg546 <= $signed(reg139[(1'h0):(1'h0)]);
                      reg547 <= reg338[(4'he):(3'h5)];
                    end
                  else
                    begin
                      reg544 <= $signed((((+reg117) ?
                          {reg95} : $unsigned(reg241)) << reg285[(3'h6):(1'h1)]));
                      reg545 <= (($unsigned({reg21}) != $signed(reg415[(3'h7):(2'h2)])) * {((8'ha1) != (~|(8'ha2)))});
                    end
                  for (forvar548 = (1'h0); (forvar548 < (1'h0)); forvar548 = (forvar548 + (1'h1)))
                    begin
                      reg549 <= reg338;
                      reg550 <= (&reg146);
                      reg551 <= ((~&(^$signed(reg138))) ?
                          {{(reg367 ?
                                      reg418 : (8'hb2))}} : ($signed($signed(reg549)) ?
                              reg360[(4'ha):(4'ha)] : $unsigned(reg338[(3'h6):(1'h0)])));
                      reg552 <= reg489[(4'ha):(1'h0)];
                    end
                  for (forvar553 = (1'h0); (forvar553 < (2'h3)); forvar553 = (forvar553 + (1'h1)))
                    begin
                      reg554 <= (forvar522[(4'ha):(3'h4)] ?
                          (($signed(reg446) ?
                              {(8'ha1)} : (forvar521 ?
                                  reg125 : reg18)) < forvar463) : reg187);
                    end
                end
              for (forvar555 = (1'h0); (forvar555 < (1'h0)); forvar555 = (forvar555 + (1'h1)))
                begin
                  if (($unsigned((~^$unsigned((8'h9c)))) ?
                      ($unsigned(reg192[(1'h1):(1'h0)]) ?
                          $signed($signed(reg308)) : $signed((~^reg469))) : ((8'hb3) <= ({reg368} * reg182[(3'h6):(3'h6)]))))
                    begin
                      reg556 <= (~&reg391[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg556 <= {reg370};
                      reg557 <= reg349[(1'h1):(1'h1)];
                      reg558 <= reg472[(4'h9):(4'h8)];
                    end
                  if ((8'ha5))
                    begin
                      reg559 <= $signed(($signed((forvar481 * (8'haf))) ~^ forvar492));
                    end
                  else
                    begin
                      reg559 <= {(^~$signed((~reg421)))};
                    end
                  if ($signed(reg108[(3'h7):(3'h5)]))
                    begin
                      reg560 <= $signed($signed($signed((reg23 < reg279))));
                      reg561 <= $unsigned((reg206 << $signed((reg545 ?
                          reg508 : reg272))));
                      reg562 <= ($signed(reg498) > $signed($signed($unsigned(reg100))));
                    end
                  else
                    begin
                      reg560 <= $signed(($signed($unsigned(reg355)) & $signed(reg38[(1'h0):(1'h0)])));
                      reg561 <= $signed((-(!(reg231 ? (8'hb8) : reg227))));
                      reg562 <= (reg220 ?
                          ((8'ha8) != (reg467 ?
                              reg377[(4'h9):(3'h7)] : $unsigned(reg98))) : $unsigned((+$signed(reg472))));
                      reg563 <= (reg393 ?
                          $signed(($signed(reg189) ?
                              (wire155 <= reg562) : (+reg412))) : reg377[(4'h8):(3'h4)]);
                    end
                  if ((reg452[(1'h0):(1'h0)] >> $signed({$unsigned(reg328)})))
                    begin
                      reg564 <= ($signed(((8'hb4) ?
                              (-reg182) : $unsigned(reg417))) ?
                          $signed((reg52 ?
                              $unsigned(reg469) : (8'haf))) : {reg212});
                      reg565 <= $unsigned(({(|reg22)} > (8'hb2)));
                    end
                  else
                    begin
                      reg564 <= {(reg36 ?
                              forvar553[(3'h7):(3'h5)] : $unsigned({reg150}))};
                    end
                end
              for (forvar566 = (1'h0); (forvar566 < (1'h1)); forvar566 = (forvar566 + (1'h1)))
                begin
                  if (($signed((8'haa)) ?
                      $signed(($signed(reg56) > {reg271})) : $unsigned($signed((^reg322)))))
                    begin
                      reg567 <= reg61[(3'h7):(1'h0)];
                      reg568 <= $unsigned($unsigned((-$unsigned((8'ha3)))));
                      reg569 <= ($signed($signed((reg320 ? reg17 : reg264))) ?
                          ({reg206[(4'hc):(1'h0)]} ?
                              (&$signed(reg418)) : {{forvar503}}) : ((~|reg517) ?
                              reg306 : reg351));
                      reg570 <= forvar553[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg567 <= ($unsigned(reg326) | ($signed((reg296 ?
                          reg277 : reg325)) || reg27));
                    end
                end
            end
          for (forvar571 = (1'h0); (forvar571 < (2'h3)); forvar571 = (forvar571 + (1'h1)))
            begin
              if (reg72[(4'ha):(3'h6)])
                begin
                  if ((~^reg245))
                    begin
                      reg572 <= (reg189 ^ (~&({reg283} ?
                          reg242[(4'he):(1'h1)] : (reg113 ^~ (8'haa)))));
                      reg573 <= ($signed((reg567 ?
                              reg299[(4'hb):(3'h5)] : {reg386})) ?
                          (~^((reg525 ?
                              reg193 : reg524) && $signed(reg64))) : forvar553);
                      reg574 <= {$unsigned($unsigned($signed(forvar474)))};
                      reg575 <= reg426;
                    end
                  else
                    begin
                      reg572 <= (~|(!reg234));
                      reg573 <= reg84[(4'hb):(1'h0)];
                      reg574 <= $signed(({(reg397 ? reg336 : reg275)} ?
                          reg527 : $signed($unsigned(reg352))));
                      reg575 <= ($unsigned(($signed(reg489) ?
                          (reg99 ^ reg519) : (reg557 ?
                              reg143 : reg417))) + (|$unsigned(reg71[(2'h3):(1'h1)])));
                    end
                  reg576 <= reg123[(1'h1):(1'h0)];
                  for (forvar577 = (1'h0); (forvar577 < (2'h2)); forvar577 = (forvar577 + (1'h1)))
                    begin
                      reg578 <= (~|$unsigned(((8'hb3) < $unsigned(reg15))));
                      reg579 <= reg322[(3'h5):(2'h3)];
                    end
                end
              else
                begin
                  reg572 <= (-$unsigned(reg426[(3'h7):(3'h7)]));
                  if (({$signed((reg272 ?
                          forvar452 : reg252))} + $unsigned($unsigned((reg393 ?
                      reg123 : reg531)))))
                    begin
                      reg573 <= reg256;
                      reg574 <= ((+reg116) >= $unsigned((|((8'hb2) ?
                          (8'ha5) : (8'hb0)))));
                    end
                  else
                    begin
                      reg573 <= $signed((^($signed(reg47) - (reg429 ?
                          reg487 : reg245))));
                      reg574 <= $signed(((&((8'hb3) ?
                          reg345 : reg189)) == ({(8'haf)} <= $signed(reg308))));
                      reg575 <= $unsigned($unsigned((+{reg471})));
                      reg576 <= reg564[(3'h4):(1'h0)];
                    end
                  if ($signed(reg228[(2'h3):(2'h2)]))
                    begin
                      reg577 <= ($signed($signed((8'ha6))) << (8'had));
                      reg578 <= $signed(reg523[(4'h8):(3'h7)]);
                    end
                  else
                    begin
                      reg577 <= (|(((reg337 > reg333) < ((8'ha8) ?
                          reg477 : reg32)) + $signed((reg560 == reg391))));
                      reg578 <= reg314;
                    end
                  for (forvar579 = (1'h0); (forvar579 < (1'h0)); forvar579 = (forvar579 + (1'h1)))
                    begin
                      reg580 <= (reg261 <<< reg254[(1'h0):(1'h0)]);
                      reg581 <= (($signed(reg531[(3'h4):(1'h1)]) ?
                              $signed((reg104 << (8'hb9))) : reg528) ?
                          (^forvar481[(4'hd):(3'h6)]) : {($unsigned(reg276) >= {reg40})});
                      reg582 <= ((-reg508[(2'h3):(1'h1)]) ?
                          ($unsigned(reg106[(3'h4):(2'h3)]) ?
                              ((reg342 ?
                                  reg112 : (8'h9e)) ~^ $signed(reg232)) : reg144[(3'h5):(2'h2)]) : $signed((^(reg258 ?
                              reg393 : reg354))));
                    end
                end
            end
          reg583 <= ((($signed(reg468) ? $unsigned(reg460) : $unsigned(reg35)) ?
                  (reg358[(2'h3):(2'h2)] >> (~^reg185)) : reg489[(1'h1):(1'h0)]) ?
              $signed(reg87) : ($unsigned(reg246[(2'h3):(1'h0)]) ?
                  {reg212[(1'h1):(1'h1)]} : (~^reg327)));
        end
      for (forvar584 = (1'h0); (forvar584 < (2'h2)); forvar584 = (forvar584 + (1'h1)))
        begin
          for (forvar585 = (1'h0); (forvar585 < (2'h2)); forvar585 = (forvar585 + (1'h1)))
            begin
              if ((&$unsigned(((reg84 & reg368) ?
                  $unsigned(reg444) : $unsigned(forvar528)))))
                begin
                  for (forvar586 = (1'h0); (forvar586 < (1'h1)); forvar586 = (forvar586 + (1'h1)))
                    begin
                      reg587 <= $signed((reg401 ?
                          {((8'ha3) + reg111)} : ($unsigned(reg507) && $signed(reg284))));
                      reg588 <= ($unsigned((reg302 ?
                              reg499 : ((8'hac) >= forvar541))) ?
                          (8'hb2) : reg199);
                      reg589 <= (reg588[(2'h3):(1'h0)] ?
                          (-(&$unsigned(reg486))) : ((-reg203) + ((reg45 ?
                                  reg65 : reg399) ?
                              reg424[(3'h4):(2'h3)] : reg336)));
                    end
                  if (reg344)
                    begin
                      reg590 <= {(&(+(reg130 ? reg399 : reg247)))};
                    end
                  else
                    begin
                      reg590 <= $signed({{(reg556 ? reg263 : reg92)}});
                      reg591 <= reg567[(2'h3):(2'h2)];
                      reg592 <= reg288;
                    end
                  reg593 <= $unsigned(reg529[(3'h5):(3'h4)]);
                  if ($unsigned({(~((8'hb8) ? (8'hb2) : reg313))}))
                    begin
                      reg594 <= {$signed($unsigned(reg400[(3'h6):(3'h6)]))};
                      reg595 <= (($unsigned((reg398 ^~ (8'hb2))) ~^ ($unsigned((8'h9c)) ?
                          reg125 : $signed(reg197))) >>> reg108[(3'h7):(3'h4)]);
                      reg596 <= (reg224[(4'h9):(1'h1)] ?
                          (reg91 > $unsigned((reg594 ^~ reg246))) : $unsigned((^reg593[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg594 <= (({(+(8'ha5))} - reg16) ?
                          (-$unsigned((^(8'ha3)))) : ({$signed(reg53)} ?
                              (~$signed(reg52)) : (-{reg531})));
                      reg595 <= reg61[(4'h9):(4'h8)];
                    end
                end
              else
                begin
                  if ($unsigned($unsigned(reg87[(1'h1):(1'h0)])))
                    begin
                      reg586 <= (8'ha5);
                      reg587 <= {(($signed(reg236) - ((8'hb2) ?
                              reg80 : reg241)) ~^ $signed({forvar478}))};
                      reg588 <= $signed((^$signed(reg527)));
                      reg589 <= {reg30};
                    end
                  else
                    begin
                      reg586 <= ($signed(($unsigned((8'ha6)) ^ (reg563 - reg209))) ?
                          {({reg413} ?
                                  (~|reg339) : $unsigned((8'ha5)))} : (((~reg345) << (reg406 ^~ reg440)) ?
                              (|$signed(reg71)) : (reg97 <<< (reg535 ^~ reg16))));
                      reg587 <= reg451;
                    end
                  for (forvar590 = (1'h0); (forvar590 < (1'h1)); forvar590 = (forvar590 + (1'h1)))
                    begin
                      reg591 <= $unsigned(reg65);
                      reg592 <= $unsigned(((^(reg95 > reg104)) ^~ ((~&reg260) ^~ (reg109 ?
                          reg419 : wire7))));
                    end
                end
              for (forvar597 = (1'h0); (forvar597 < (1'h1)); forvar597 = (forvar597 + (1'h1)))
                begin
                  if (($unsigned(reg323) || reg336[(2'h2):(1'h0)]))
                    begin
                      reg598 <= $signed((reg342 ?
                          $signed(reg299) : (reg340 ?
                              (reg358 | wire155) : $unsigned((8'hb9)))));
                    end
                  else
                    begin
                      reg598 <= (reg485[(1'h0):(1'h0)] ?
                          $signed((&$unsigned(reg374))) : reg439);
                      reg599 <= $unsigned(wire7[(2'h2):(1'h0)]);
                      reg600 <= $unsigned(($signed($unsigned((8'hb6))) ?
                          $unsigned($unsigned(reg499)) : {reg369[(3'h6):(3'h6)]}));
                    end
                  for (forvar601 = (1'h0); (forvar601 < (2'h2)); forvar601 = (forvar601 + (1'h1)))
                    begin
                      reg602 <= $signed((!((reg43 == reg42) ^~ (~&(8'h9e)))));
                      reg603 <= (reg249[(3'h4):(2'h3)] ^~ (^~(&reg139[(3'h7):(2'h3)])));
                      reg604 <= ($unsigned(((reg582 > forvar528) && (reg101 ?
                              reg259 : reg595))) ?
                          {(&(reg569 ?
                                  forvar541 : forvar522))} : $signed((reg477[(3'h6):(3'h6)] > {reg214})));
                      reg605 <= $signed((~(~(reg42 == reg102))));
                    end
                end
              reg606 <= (reg72[(3'h4):(2'h3)] ? reg410 : reg30[(4'h8):(1'h1)]);
              for (forvar607 = (1'h0); (forvar607 < (2'h3)); forvar607 = (forvar607 + (1'h1)))
                begin
                  reg608 <= (&(~^$signed($signed(reg278))));
                end
            end
        end
    end
  assign wire609 = {reg354};
  assign wire610 = $signed(((|{reg48}) || reg261[(1'h0):(1'h0)]));
  module611 #() modinst830 (wire829, clk, reg600, wire8, reg91, reg490, reg379);
  assign wire831 = ((((reg370 + reg472) >> (+reg272)) ?
                       reg444 : (&(wire155 <= reg111))) < $signed((reg326 != $signed(reg36))));
  assign wire832 = (reg482 ? reg425[(1'h1):(1'h1)] : $signed(reg456));
  assign wire833 = $signed($unsigned($signed(reg22)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module611
#(parameter param828 = ((({(8'ha6)} ? (8'hb5) : (!(8'hba))) ? ((&(8'hb4)) ? ((8'hb2) > (8'ha3)) : (~|(8'hb3))) : (-(-(8'hba)))) ~^ ({((8'had) || (8'ha7))} && ((+(8'hb3)) ~^ ((8'hb5) * (8'ha2))))))
(y, clk, wire616, wire615, wire614, wire613, wire612);
  output wire [(32'h870):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire616;
  input wire [(2'h2):(1'h0)] wire615;
  input wire signed [(3'h4):(1'h0)] wire614;
  input wire signed [(3'h5):(1'h0)] wire613;
  input wire [(4'h8):(1'h0)] wire612;
  wire [(4'hc):(1'h0)] wire827;
  wire [(3'h5):(1'h0)] wire826;
  wire [(3'h7):(1'h0)] wire825;
  wire signed [(3'h6):(1'h0)] wire824;
  wire [(3'h7):(1'h0)] wire823;
  wire signed [(4'ha):(1'h0)] wire822;
  wire signed [(3'h7):(1'h0)] wire821;
  wire signed [(2'h3):(1'h0)] wire820;
  wire signed [(4'hf):(1'h0)] wire781;
  wire [(4'hc):(1'h0)] wire780;
  wire [(3'h7):(1'h0)] wire779;
  wire signed [(4'h8):(1'h0)] wire778;
  wire signed [(4'hf):(1'h0)] wire617;
  reg signed [(3'h4):(1'h0)] reg788 = (1'h0);
  reg [(4'hd):(1'h0)] reg819 = (1'h0);
  reg [(2'h2):(1'h0)] reg818 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg817 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg814 = (1'h0);
  reg [(2'h3):(1'h0)] reg813 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg811 = (1'h0);
  reg signed [(4'he):(1'h0)] reg810 = (1'h0);
  reg [(3'h4):(1'h0)] reg809 = (1'h0);
  reg [(4'ha):(1'h0)] reg806 = (1'h0);
  reg [(4'he):(1'h0)] reg804 = (1'h0);
  reg [(2'h2):(1'h0)] reg799 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg807 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg805 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg803 = (1'h0);
  reg [(3'h7):(1'h0)] reg802 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg801 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg800 = (1'h0);
  reg [(3'h4):(1'h0)] reg798 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg797 = (1'h0);
  reg [(4'hd):(1'h0)] reg795 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg794 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg793 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg792 = (1'h0);
  reg [(4'he):(1'h0)] reg789 = (1'h0);
  reg [(4'hd):(1'h0)] reg787 = (1'h0);
  reg [(4'h9):(1'h0)] reg786 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg784 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg783 = (1'h0);
  reg [(2'h3):(1'h0)] reg777 = (1'h0);
  reg [(4'hf):(1'h0)] reg716 = (1'h0);
  reg [(3'h5):(1'h0)] reg709 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg754 = (1'h0);
  reg [(4'h9):(1'h0)] reg775 = (1'h0);
  reg [(3'h5):(1'h0)] reg774 = (1'h0);
  reg [(4'hb):(1'h0)] reg773 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg771 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg770 = (1'h0);
  reg [(3'h6):(1'h0)] reg769 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg768 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg767 = (1'h0);
  reg [(4'hc):(1'h0)] reg766 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg765 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg762 = (1'h0);
  reg [(4'h8):(1'h0)] reg761 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg760 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg759 = (1'h0);
  reg [(4'h8):(1'h0)] reg758 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg757 = (1'h0);
  reg [(4'h9):(1'h0)] reg756 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg755 = (1'h0);
  reg [(4'ha):(1'h0)] reg753 = (1'h0);
  reg [(3'h6):(1'h0)] reg752 = (1'h0);
  reg [(5'h10):(1'h0)] reg751 = (1'h0);
  reg [(4'hd):(1'h0)] reg748 = (1'h0);
  reg [(4'hd):(1'h0)] reg747 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg746 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg745 = (1'h0);
  reg [(2'h2):(1'h0)] reg744 = (1'h0);
  reg [(4'h9):(1'h0)] reg743 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg741 = (1'h0);
  reg [(4'ha):(1'h0)] reg740 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg737 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg734 = (1'h0);
  reg [(5'h10):(1'h0)] reg733 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg732 = (1'h0);
  reg [(3'h5):(1'h0)] reg731 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg730 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg729 = (1'h0);
  reg [(4'hd):(1'h0)] reg728 = (1'h0);
  reg [(3'h6):(1'h0)] reg727 = (1'h0);
  reg [(4'hf):(1'h0)] reg726 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg725 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg724 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg722 = (1'h0);
  reg [(5'h10):(1'h0)] reg721 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg720 = (1'h0);
  reg [(4'hb):(1'h0)] reg719 = (1'h0);
  reg [(4'hb):(1'h0)] reg718 = (1'h0);
  reg [(4'hf):(1'h0)] reg717 = (1'h0);
  reg [(3'h5):(1'h0)] reg715 = (1'h0);
  reg [(3'h6):(1'h0)] reg714 = (1'h0);
  reg [(3'h4):(1'h0)] reg710 = (1'h0);
  reg [(4'hb):(1'h0)] reg707 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg713 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg712 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg711 = (1'h0);
  reg [(4'hf):(1'h0)] reg708 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg706 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg705 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg704 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg703 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg702 = (1'h0);
  reg [(3'h7):(1'h0)] reg701 = (1'h0);
  reg [(4'hf):(1'h0)] reg700 = (1'h0);
  reg [(4'ha):(1'h0)] reg699 = (1'h0);
  reg [(4'hc):(1'h0)] reg696 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg694 = (1'h0);
  reg [(4'h9):(1'h0)] reg693 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg692 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg691 = (1'h0);
  reg [(4'hf):(1'h0)] reg690 = (1'h0);
  reg signed [(4'he):(1'h0)] reg688 = (1'h0);
  reg [(3'h5):(1'h0)] reg687 = (1'h0);
  reg signed [(4'he):(1'h0)] reg686 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg685 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg682 = (1'h0);
  reg [(2'h2):(1'h0)] reg675 = (1'h0);
  reg [(2'h3):(1'h0)] reg673 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg666 = (1'h0);
  reg [(3'h4):(1'h0)] reg663 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg684 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg683 = (1'h0);
  reg [(4'hb):(1'h0)] reg681 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg680 = (1'h0);
  reg [(2'h2):(1'h0)] reg679 = (1'h0);
  reg [(4'h8):(1'h0)] reg678 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg676 = (1'h0);
  reg signed [(4'he):(1'h0)] reg674 = (1'h0);
  reg [(2'h3):(1'h0)] reg672 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg671 = (1'h0);
  reg [(3'h5):(1'h0)] reg670 = (1'h0);
  reg [(3'h5):(1'h0)] reg668 = (1'h0);
  reg [(4'h9):(1'h0)] reg667 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg665 = (1'h0);
  reg [(4'h9):(1'h0)] reg664 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg661 = (1'h0);
  reg [(4'hf):(1'h0)] reg660 = (1'h0);
  reg [(3'h7):(1'h0)] reg659 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg658 = (1'h0);
  reg [(4'hf):(1'h0)] reg657 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg656 = (1'h0);
  reg [(3'h6):(1'h0)] reg655 = (1'h0);
  reg [(3'h6):(1'h0)] reg654 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg652 = (1'h0);
  reg [(4'he):(1'h0)] reg651 = (1'h0);
  reg [(3'h7):(1'h0)] reg650 = (1'h0);
  reg [(5'h10):(1'h0)] reg642 = (1'h0);
  reg [(3'h4):(1'h0)] reg647 = (1'h0);
  reg [(4'h8):(1'h0)] reg646 = (1'h0);
  reg [(3'h6):(1'h0)] reg645 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg644 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg643 = (1'h0);
  reg [(3'h4):(1'h0)] reg641 = (1'h0);
  reg [(2'h2):(1'h0)] reg640 = (1'h0);
  reg signed [(4'he):(1'h0)] reg639 = (1'h0);
  reg signed [(4'he):(1'h0)] reg638 = (1'h0);
  reg [(4'h9):(1'h0)] reg637 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg636 = (1'h0);
  reg [(4'hf):(1'h0)] reg635 = (1'h0);
  reg [(2'h2):(1'h0)] reg634 = (1'h0);
  reg [(4'he):(1'h0)] reg633 = (1'h0);
  reg [(4'h9):(1'h0)] reg632 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg631 = (1'h0);
  reg [(3'h6):(1'h0)] reg630 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg628 = (1'h0);
  reg [(3'h6):(1'h0)] reg627 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg621 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg626 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg625 = (1'h0);
  reg [(3'h4):(1'h0)] reg624 = (1'h0);
  reg [(4'hb):(1'h0)] reg623 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg622 = (1'h0);
  reg [(4'h8):(1'h0)] reg619 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar816 = (1'h0);
  reg [(4'hc):(1'h0)] forvar815 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar812 = (1'h0);
  reg [(4'h8):(1'h0)] forvar808 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar806 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar804 = (1'h0);
  reg [(4'hb):(1'h0)] forvar799 = (1'h0);
  reg [(2'h2):(1'h0)] forvar796 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar791 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar790 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar788 = (1'h0);
  reg [(3'h4):(1'h0)] forvar785 = (1'h0);
  reg [(4'hc):(1'h0)] forvar782 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar776 = (1'h0);
  reg [(4'ha):(1'h0)] forvar724 = (1'h0);
  reg [(2'h2):(1'h0)] forvar722 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar718 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar714 = (1'h0);
  reg [(4'hd):(1'h0)] forvar772 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar764 = (1'h0);
  reg [(3'h4):(1'h0)] forvar763 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar754 = (1'h0);
  reg [(3'h7):(1'h0)] forvar750 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar749 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar742 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar739 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar738 = (1'h0);
  reg [(5'h10):(1'h0)] forvar736 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar735 = (1'h0);
  reg [(2'h3):(1'h0)] forvar732 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar723 = (1'h0);
  reg [(4'ha):(1'h0)] forvar716 = (1'h0);
  reg [(4'h8):(1'h0)] forvar712 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar708 = (1'h0);
  reg [(4'hd):(1'h0)] forvar710 = (1'h0);
  reg [(3'h7):(1'h0)] forvar709 = (1'h0);
  reg [(3'h4):(1'h0)] forvar707 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar698 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar697 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar695 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar690 = (1'h0);
  reg [(2'h2):(1'h0)] forvar689 = (1'h0);
  reg [(4'hb):(1'h0)] forvar681 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar674 = (1'h0);
  reg [(4'hd):(1'h0)] forvar664 = (1'h0);
  reg [(3'h5):(1'h0)] forvar682 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar677 = (1'h0);
  reg [(4'h9):(1'h0)] forvar675 = (1'h0);
  reg [(5'h10):(1'h0)] forvar673 = (1'h0);
  reg [(2'h3):(1'h0)] forvar669 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar666 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar663 = (1'h0);
  reg [(4'he):(1'h0)] forvar662 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar625 = (1'h0);
  reg [(3'h7):(1'h0)] forvar622 = (1'h0);
  reg [(4'he):(1'h0)] forvar653 = (1'h0);
  reg [(4'h8):(1'h0)] forvar649 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar648 = (1'h0);
  reg [(3'h6):(1'h0)] forvar641 = (1'h0);
  reg [(5'h10):(1'h0)] forvar638 = (1'h0);
  reg [(3'h5):(1'h0)] forvar642 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar629 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar621 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar620 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar618 = (1'h0);
  assign y = {wire827,
                 wire826,
                 wire825,
                 wire824,
                 wire823,
                 wire822,
                 wire821,
                 wire820,
                 wire781,
                 wire780,
                 wire779,
                 wire778,
                 wire617,
                 reg788,
                 reg819,
                 reg818,
                 reg817,
                 reg814,
                 reg813,
                 reg811,
                 reg810,
                 reg809,
                 reg806,
                 reg804,
                 reg799,
                 reg807,
                 reg805,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 reg798,
                 reg797,
                 reg795,
                 reg794,
                 reg793,
                 reg792,
                 reg789,
                 reg787,
                 reg786,
                 reg784,
                 reg783,
                 reg777,
                 reg716,
                 reg709,
                 reg754,
                 reg775,
                 reg774,
                 reg773,
                 reg771,
                 reg770,
                 reg769,
                 reg768,
                 reg767,
                 reg766,
                 reg765,
                 reg762,
                 reg761,
                 reg760,
                 reg759,
                 reg758,
                 reg757,
                 reg756,
                 reg755,
                 reg753,
                 reg752,
                 reg751,
                 reg748,
                 reg747,
                 reg746,
                 reg745,
                 reg744,
                 reg743,
                 reg741,
                 reg740,
                 reg737,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 reg730,
                 reg729,
                 reg728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 reg722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg715,
                 reg714,
                 reg710,
                 reg707,
                 reg713,
                 reg712,
                 reg711,
                 reg708,
                 reg706,
                 reg705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 reg699,
                 reg696,
                 reg694,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg688,
                 reg687,
                 reg686,
                 reg685,
                 reg682,
                 reg675,
                 reg673,
                 reg666,
                 reg663,
                 reg684,
                 reg683,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 reg676,
                 reg674,
                 reg672,
                 reg671,
                 reg670,
                 reg668,
                 reg667,
                 reg665,
                 reg664,
                 reg661,
                 reg660,
                 reg659,
                 reg658,
                 reg657,
                 reg656,
                 reg655,
                 reg654,
                 reg652,
                 reg651,
                 reg650,
                 reg642,
                 reg647,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 reg641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 reg628,
                 reg627,
                 reg621,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 reg619,
                 forvar816,
                 forvar815,
                 forvar812,
                 forvar808,
                 forvar806,
                 forvar804,
                 forvar799,
                 forvar796,
                 forvar791,
                 forvar790,
                 forvar788,
                 forvar785,
                 forvar782,
                 forvar776,
                 forvar724,
                 forvar722,
                 forvar718,
                 forvar714,
                 forvar772,
                 forvar764,
                 forvar763,
                 forvar754,
                 forvar750,
                 forvar749,
                 forvar742,
                 forvar739,
                 forvar738,
                 forvar736,
                 forvar735,
                 forvar732,
                 forvar723,
                 forvar716,
                 forvar712,
                 forvar708,
                 forvar710,
                 forvar709,
                 forvar707,
                 forvar698,
                 forvar697,
                 forvar695,
                 forvar690,
                 forvar689,
                 forvar681,
                 forvar674,
                 forvar664,
                 forvar682,
                 forvar677,
                 forvar675,
                 forvar673,
                 forvar669,
                 forvar666,
                 forvar663,
                 forvar662,
                 forvar625,
                 forvar622,
                 forvar653,
                 forvar649,
                 forvar648,
                 forvar641,
                 forvar638,
                 forvar642,
                 forvar629,
                 forvar621,
                 forvar620,
                 forvar618,
                 (1'h0)};
  assign wire617 = (+(+(~&$unsigned(wire616))));
  always
    @(posedge clk) begin
      for (forvar618 = (1'h0); (forvar618 < (1'h1)); forvar618 = (forvar618 + (1'h1)))
        begin
          reg619 <= ((-wire612[(3'h5):(3'h5)]) ?
              wire617 : {(wire616[(3'h4):(2'h3)] ?
                      wire614 : (wire617 * (8'hab)))});
        end
      for (forvar620 = (1'h0); (forvar620 < (1'h0)); forvar620 = (forvar620 + (1'h1)))
        begin
          if ($unsigned(($unsigned($signed(wire614)) ?
              {(forvar618 == wire613)} : ((&wire616) ?
                  (wire615 > (8'ha7)) : wire614[(1'h1):(1'h0)]))))
            begin
              if ((({(wire613 != wire616)} ?
                      (8'ha8) : $unsigned((wire615 ^~ wire615))) ?
                  {($signed(wire615) ?
                          (^forvar618) : {forvar618})} : {((8'haa) != $unsigned(wire614))}))
                begin
                  for (forvar621 = (1'h0); (forvar621 < (2'h3)); forvar621 = (forvar621 + (1'h1)))
                    begin
                      reg622 <= $signed(wire617);
                      reg623 <= wire613;
                    end
                  if ({$signed((^{reg622}))})
                    begin
                      reg624 <= (~&(^((^~forvar618) ?
                          (forvar621 ?
                              reg622 : forvar621) : $unsigned(wire614))));
                      reg625 <= reg622;
                    end
                  else
                    begin
                      reg624 <= wire612[(2'h2):(1'h0)];
                      reg625 <= $unsigned($signed((^(reg622 ?
                          (8'ha5) : reg624))));
                      reg626 <= ((|$unsigned(((8'h9d) ? reg624 : wire616))) ?
                          ((~(wire613 ? (8'hb4) : forvar618)) ?
                              (wire615[(1'h0):(1'h0)] ?
                                  (~|reg625) : forvar620) : ({forvar620} ?
                                  (wire617 ?
                                      (8'h9c) : wire614) : ((8'ha0) * reg623))) : $signed({$signed(reg622)}));
                    end
                end
              else
                begin
                  reg621 <= $signed((~|((~&wire617) ? wire615 : (~&(8'hb5)))));
                  if (reg621)
                    begin
                      reg622 <= (reg622 ?
                          (~|$unsigned($unsigned(reg625))) : {reg621[(4'h8):(3'h6)]});
                      reg623 <= {wire615};
                      reg624 <= $unsigned($unsigned($unsigned((reg625 <<< forvar621))));
                    end
                  else
                    begin
                      reg622 <= $signed(((wire612 ?
                          wire612[(3'h6):(3'h4)] : (-reg625)) || $unsigned(wire612[(3'h5):(3'h5)])));
                      reg623 <= (((reg624 ?
                                  (wire616 >> reg624) : (wire612 & reg619)) ?
                              ((8'ha2) * (reg626 & reg621)) : $unsigned($unsigned(forvar618))) ?
                          ((^~(forvar618 == (8'hab))) - {$unsigned((8'hab))}) : forvar618);
                      reg624 <= (forvar621[(4'hd):(3'h4)] ?
                          (-forvar620[(3'h4):(3'h4)]) : $signed($signed(wire617[(4'h8):(4'h8)])));
                      reg625 <= $signed((~((wire614 ? reg626 : reg619) ?
                          wire612 : $signed(reg624))));
                    end
                  if ($unsigned({{wire617}}))
                    begin
                      reg626 <= (({$unsigned((8'had))} < reg625[(2'h2):(2'h2)]) != (|$signed(reg624[(2'h3):(1'h0)])));
                      reg627 <= (!$signed(reg621));
                      reg628 <= $unsigned(($signed($unsigned((8'hb8))) ?
                          $signed((reg624 ? reg619 : reg623)) : (~{reg626})));
                    end
                  else
                    begin
                      reg626 <= (^~((((8'hab) ?
                              reg626 : wire612) <<< (forvar618 ?
                              reg622 : wire613)) ?
                          $unsigned((reg627 ?
                              forvar618 : wire615)) : {forvar618[(3'h6):(2'h2)]}));
                      reg627 <= ({$signed(wire617)} <<< $signed(wire617));
                    end
                end
              for (forvar629 = (1'h0); (forvar629 < (2'h2)); forvar629 = (forvar629 + (1'h1)))
                begin
                  if (((((wire617 ~^ wire613) ?
                          wire615[(1'h1):(1'h0)] : reg625) - ({reg622} - (reg622 ^~ forvar618))) ?
                      (~$unsigned((-(8'had)))) : reg619))
                    begin
                      reg630 <= (^~(reg619[(1'h1):(1'h0)] * {$signed(wire617)}));
                      reg631 <= $unsigned({$unsigned($unsigned((8'hb9)))});
                      reg632 <= {reg619[(4'h8):(2'h2)]};
                      reg633 <= (^~forvar629);
                    end
                  else
                    begin
                      reg630 <= {forvar621[(3'h6):(3'h4)]};
                      reg631 <= (8'ha8);
                    end
                  if (forvar629[(2'h3):(1'h0)])
                    begin
                      reg634 <= ((^((forvar618 ? wire612 : forvar621) ?
                          (reg633 ?
                              (8'hb2) : (8'ha8)) : $signed(wire616))) + (((8'ha4) ?
                              (forvar618 ^ reg628) : reg633[(4'hd):(4'h8)]) ?
                          (forvar629[(1'h0):(1'h0)] == ((8'hb9) ?
                              wire617 : reg621)) : {(reg627 >= reg626)}));
                    end
                  else
                    begin
                      reg634 <= $signed(reg624);
                    end
                  if (($signed(reg622[(3'h4):(1'h0)]) >>> $unsigned($unsigned($unsigned(wire613)))))
                    begin
                      reg635 <= (8'hb0);
                      reg636 <= ($signed(forvar621[(3'h6):(3'h5)]) > ((!{reg624}) + $unsigned((wire616 != reg627))));
                      reg637 <= ((~|{reg635[(4'hb):(4'hb)]}) ?
                          ($unsigned((reg622 ?
                              forvar621 : reg619)) << forvar618[(4'h8):(3'h4)]) : $unsigned((~&(reg630 && reg636))));
                    end
                  else
                    begin
                      reg635 <= $signed(($unsigned(reg637[(3'h5):(1'h1)]) > $signed($unsigned(reg625))));
                      reg636 <= forvar618[(2'h3):(1'h0)];
                    end
                end
              if ((reg621[(4'ha):(3'h6)] >> {(^forvar629)}))
                begin
                  if ((~^$signed((reg619 >>> (wire615 ? (8'haf) : reg632)))))
                    begin
                      reg638 <= (~&$signed($signed(wire617)));
                      reg639 <= wire617[(4'h9):(4'h8)];
                      reg640 <= ({(^(forvar618 ? reg631 : forvar620))} ?
                          (^$signed(forvar620[(3'h4):(1'h0)])) : reg619[(3'h6):(2'h3)]);
                      reg641 <= $signed((reg632[(2'h3):(2'h3)] ?
                          {(reg639 ?
                                  reg626 : reg632)} : ({reg624} != $signed(reg638))));
                    end
                  else
                    begin
                      reg638 <= {(~^reg622)};
                      reg639 <= (+((~^forvar629[(2'h2):(2'h2)]) > $unsigned((&wire615))));
                      reg640 <= (~&reg622);
                      reg641 <= wire614;
                    end
                  for (forvar642 = (1'h0); (forvar642 < (1'h0)); forvar642 = (forvar642 + (1'h1)))
                    begin
                      reg643 <= reg634;
                      reg644 <= (forvar629[(1'h1):(1'h1)] ?
                          $signed(((reg631 + reg638) ?
                              reg637 : (|forvar629))) : ($unsigned((~|reg638)) ?
                              (8'ha5) : ((-(8'hb0)) ?
                                  (wire615 ~^ reg637) : (wire615 * (8'hb8)))));
                    end
                  if ($signed({(wire614 >> (wire614 & reg626))}))
                    begin
                      reg645 <= ((($signed(reg641) <= (8'hac)) ?
                          (|(reg634 ? reg622 : reg627)) : $signed((reg635 ?
                              wire615 : reg641))) * (wire614 ?
                          ((!reg626) ?
                              $signed((8'ha3)) : reg636) : {(&reg633)}));
                    end
                  else
                    begin
                      reg645 <= ($unsigned(reg627) ?
                          $signed({$unsigned(reg619)}) : reg644);
                      reg646 <= forvar618;
                      reg647 <= reg639;
                    end
                end
              else
                begin
                  for (forvar638 = (1'h0); (forvar638 < (2'h2)); forvar638 = (forvar638 + (1'h1)))
                    begin
                      reg639 <= $unsigned($unsigned((wire614 ^~ $unsigned(forvar642))));
                    end
                  reg640 <= ((|(&((8'had) ?
                      reg631 : reg630))) <<< wire613[(3'h5):(1'h1)]);
                  for (forvar641 = (1'h0); (forvar641 < (1'h0)); forvar641 = (forvar641 + (1'h1)))
                    begin
                      reg642 <= reg621;
                      reg643 <= ($unsigned(reg625[(3'h4):(1'h1)]) ?
                          (8'ha7) : $signed(reg625));
                      reg644 <= wire616[(4'ha):(3'h4)];
                    end
                  if (wire616)
                    begin
                      reg645 <= (reg634 * $unsigned(reg638));
                      reg646 <= reg623[(4'ha):(3'h5)];
                      reg647 <= $unsigned({({(8'ha2)} && (+reg632))});
                    end
                  else
                    begin
                      reg645 <= ((forvar641 - ($unsigned(reg619) > reg627)) >> {((^~reg635) >> reg639)});
                      reg646 <= (^{$unsigned((wire615 ? reg642 : reg646))});
                    end
                end
              for (forvar648 = (1'h0); (forvar648 < (2'h2)); forvar648 = (forvar648 + (1'h1)))
                begin
                  for (forvar649 = (1'h0); (forvar649 < (1'h1)); forvar649 = (forvar649 + (1'h1)))
                    begin
                      reg650 <= (($signed($unsigned(forvar638)) ?
                              {wire612[(3'h5):(1'h0)]} : ((reg639 * reg640) + (+forvar621))) ?
                          reg623[(2'h3):(2'h2)] : $unsigned((&(reg619 <= reg624))));
                      reg651 <= wire615[(1'h0):(1'h0)];
                      reg652 <= $signed((reg651 >> $signed(reg633)));
                    end
                  for (forvar653 = (1'h0); (forvar653 < (2'h2)); forvar653 = (forvar653 + (1'h1)))
                    begin
                      reg654 <= $unsigned($unsigned((8'h9d)));
                    end
                  if (($unsigned($unsigned($unsigned(forvar621))) < $unsigned(reg641[(2'h2):(2'h2)])))
                    begin
                      reg655 <= reg639[(4'h9):(3'h5)];
                      reg656 <= (&$unsigned(((&reg641) || reg636)));
                      reg657 <= ($signed(((reg641 ?
                          reg646 : (8'hba)) & reg642)) - ((!(wire614 ?
                          reg641 : wire616)) && (-reg639[(4'hd):(4'ha)])));
                    end
                  else
                    begin
                      reg655 <= wire613[(2'h3):(2'h3)];
                    end
                  if ($unsigned((forvar629 ?
                      {$signed((8'hb6))} : ((reg634 << reg642) ?
                          (|(8'ha8)) : (reg655 ? forvar620 : reg642)))))
                    begin
                      reg658 <= wire612[(2'h3):(2'h2)];
                      reg659 <= $unsigned($unsigned(((~wire617) < $signed(reg630))));
                    end
                  else
                    begin
                      reg658 <= reg650[(2'h3):(2'h3)];
                      reg659 <= ({($unsigned(wire615) && wire616)} <= reg631[(3'h7):(1'h0)]);
                      reg660 <= (-reg621[(4'hb):(4'h9)]);
                      reg661 <= {reg631[(3'h7):(3'h7)]};
                    end
                end
            end
          else
            begin
              for (forvar621 = (1'h0); (forvar621 < (1'h0)); forvar621 = (forvar621 + (1'h1)))
                begin
                  for (forvar622 = (1'h0); (forvar622 < (2'h2)); forvar622 = (forvar622 + (1'h1)))
                    begin
                      reg623 <= $signed(reg650[(3'h7):(1'h1)]);
                    end
                end
              if ((($signed($unsigned(forvar629)) ?
                  reg652[(1'h0):(1'h0)] : (!(~forvar649))) >>> (|$signed(forvar642))))
                begin
                  if (wire612[(1'h0):(1'h0)])
                    begin
                      reg624 <= $signed((&$signed({reg626})));
                      reg625 <= reg655[(2'h3):(1'h0)];
                      reg626 <= $signed(reg622[(3'h4):(2'h3)]);
                      reg627 <= $unsigned(forvar638);
                    end
                  else
                    begin
                      reg624 <= {(reg656 ?
                              ($signed((8'ha9)) ?
                                  reg631[(4'hb):(3'h7)] : wire612) : (reg632[(4'h9):(4'h9)] ?
                                  reg630[(1'h1):(1'h1)] : $unsigned(reg650)))};
                      reg625 <= (^~$signed(((8'ha9) ?
                          $unsigned(reg658) : reg634)));
                      reg626 <= (~^$signed($signed((reg647 < reg632))));
                    end
                end
              else
                begin
                  reg624 <= (^reg640);
                  for (forvar625 = (1'h0); (forvar625 < (1'h0)); forvar625 = (forvar625 + (1'h1)))
                    begin
                      reg626 <= forvar621;
                      reg627 <= reg632;
                      reg628 <= ($unsigned($signed(reg661)) ?
                          $unsigned($unsigned(reg619)) : reg657[(1'h1):(1'h1)]);
                    end
                end
            end
          if ($signed((($signed(reg646) ? $signed(reg633) : (~&forvar648)) ?
              reg651 : forvar622[(3'h4):(2'h3)])))
            begin
              for (forvar662 = (1'h0); (forvar662 < (1'h0)); forvar662 = (forvar662 + (1'h1)))
                begin
                  for (forvar663 = (1'h0); (forvar663 < (2'h3)); forvar663 = (forvar663 + (1'h1)))
                    begin
                      reg664 <= $signed(((~^(&wire613)) * ($unsigned(reg654) ?
                          (reg641 ? reg645 : wire614) : wire614)));
                      reg665 <= reg630[(2'h3):(1'h1)];
                    end
                  for (forvar666 = (1'h0); (forvar666 < (1'h1)); forvar666 = (forvar666 + (1'h1)))
                    begin
                      reg667 <= (wire616 ?
                          (^~$signed({reg657})) : ($unsigned($signed(wire612)) ?
                              ($unsigned(wire612) + reg656) : ((reg621 >>> (8'ha7)) - $signed(reg634))));
                      reg668 <= forvar642;
                    end
                  for (forvar669 = (1'h0); (forvar669 < (2'h3)); forvar669 = (forvar669 + (1'h1)))
                    begin
                      reg670 <= reg667;
                      reg671 <= $unsigned(reg639);
                    end
                  reg672 <= (8'hb3);
                end
              for (forvar673 = (1'h0); (forvar673 < (1'h1)); forvar673 = (forvar673 + (1'h1)))
                begin
                  reg674 <= {$unsigned($unsigned({forvar625}))};
                  for (forvar675 = (1'h0); (forvar675 < (1'h0)); forvar675 = (forvar675 + (1'h1)))
                    begin
                      reg676 <= ($signed((forvar648 + $signed((8'hb5)))) < (8'ha9));
                    end
                end
              for (forvar677 = (1'h0); (forvar677 < (2'h2)); forvar677 = (forvar677 + (1'h1)))
                begin
                  if ({reg655})
                    begin
                      reg678 <= reg619[(3'h5):(1'h0)];
                      reg679 <= ($unsigned((+(reg639 ~^ reg643))) ~^ $signed((reg630 == reg665[(4'h8):(3'h7)])));
                      reg680 <= $signed({({forvar662} ?
                              (~&reg645) : {reg639})});
                    end
                  else
                    begin
                      reg678 <= reg619[(1'h0):(1'h0)];
                    end
                  reg681 <= reg651;
                  for (forvar682 = (1'h0); (forvar682 < (1'h0)); forvar682 = (forvar682 + (1'h1)))
                    begin
                      reg683 <= reg627[(2'h2):(1'h0)];
                      reg684 <= {($unsigned((forvar622 ?
                              reg625 : reg651)) <<< reg658[(2'h3):(1'h1)])};
                    end
                end
            end
          else
            begin
              for (forvar662 = (1'h0); (forvar662 < (1'h0)); forvar662 = (forvar662 + (1'h1)))
                begin
                  reg663 <= ((forvar648[(4'h8):(2'h3)] ?
                          $unsigned(reg645) : ((&(8'hb6)) ?
                              reg641[(1'h0):(1'h0)] : $signed(reg679))) ?
                      reg639[(3'h4):(2'h3)] : (~|wire617[(3'h5):(1'h0)]));
                end
              for (forvar664 = (1'h0); (forvar664 < (1'h1)); forvar664 = (forvar664 + (1'h1)))
                begin
                  if ({wire617})
                    begin
                      reg665 <= $signed((reg658[(3'h4):(3'h4)] && wire616[(3'h7):(3'h5)]));
                      reg666 <= (wire617 ?
                          ((~&(wire614 ? reg625 : forvar622)) ?
                              $signed(((8'hb8) * reg658)) : $unsigned((forvar642 << forvar663))) : reg631[(3'h7):(3'h5)]);
                      reg667 <= $signed($unsigned(((forvar629 ^~ reg634) ?
                          (forvar673 ? reg628 : forvar664) : $signed(reg666))));
                      reg668 <= {($unsigned(((8'h9c) <= reg621)) ?
                              ($signed(forvar666) * (wire614 ^ reg646)) : reg664[(3'h5):(1'h0)])};
                    end
                  else
                    begin
                      reg665 <= ((~$unsigned((reg621 < reg642))) <= (~^(~^$unsigned(reg650))));
                      reg666 <= (~&reg658);
                      reg667 <= forvar673[(3'h4):(2'h2)];
                      reg668 <= ((((|reg642) ~^ $signed(reg632)) <<< reg679[(2'h2):(2'h2)]) >>> $unsigned(reg652[(4'ha):(3'h6)]));
                    end
                  for (forvar669 = (1'h0); (forvar669 < (2'h2)); forvar669 = (forvar669 + (1'h1)))
                    begin
                      reg670 <= (((forvar663[(2'h3):(2'h2)] << (~reg643)) ?
                          ((!(8'ha3)) ?
                              $unsigned(reg659) : reg634) : ((&reg624) ?
                              (~&reg655) : (8'h9d))) & reg672[(1'h1):(1'h1)]);
                      reg671 <= (~|({forvar673[(1'h1):(1'h1)]} || (reg684 ~^ $signed(reg622))));
                      reg672 <= reg619;
                      reg673 <= (reg641 ?
                          reg660 : $signed(($unsigned(reg659) && (reg644 | forvar666))));
                    end
                  for (forvar674 = (1'h0); (forvar674 < (2'h2)); forvar674 = (forvar674 + (1'h1)))
                    begin
                      reg675 <= {(~forvar622[(1'h0):(1'h0)])};
                      reg676 <= (8'had);
                    end
                end
              for (forvar677 = (1'h0); (forvar677 < (1'h0)); forvar677 = (forvar677 + (1'h1)))
                begin
                  if ((^reg639))
                    begin
                      reg678 <= reg661[(1'h1):(1'h0)];
                      reg679 <= $unsigned(reg679[(1'h0):(1'h0)]);
                      reg680 <= ((|(reg644 ?
                          forvar662[(4'ha):(3'h4)] : (forvar666 ?
                              (8'ha2) : forvar664))) | $signed(reg621[(4'hd):(3'h6)]));
                    end
                  else
                    begin
                      reg678 <= forvar642;
                      reg679 <= reg639[(4'hd):(4'h8)];
                    end
                  for (forvar681 = (1'h0); (forvar681 < (1'h1)); forvar681 = (forvar681 + (1'h1)))
                    begin
                      reg682 <= {wire615[(2'h2):(2'h2)]};
                      reg683 <= (^reg640);
                    end
                  if (wire616[(3'h5):(1'h1)])
                    begin
                      reg684 <= forvar648;
                    end
                  else
                    begin
                      reg684 <= ((((forvar664 * reg651) <<< $signed(reg656)) ?
                              reg641 : $signed((reg642 || reg668))) ?
                          ($signed(forvar625) ?
                              reg668 : (~|{(8'ha2)})) : $unsigned($unsigned((8'ha5))));
                      reg685 <= (forvar625[(1'h1):(1'h1)] ?
                          (^(8'hb3)) : $signed((|$unsigned(reg658))));
                      reg686 <= (+$signed(reg640[(1'h1):(1'h0)]));
                    end
                  if ((^forvar648))
                    begin
                      reg687 <= reg656;
                    end
                  else
                    begin
                      reg687 <= ({$unsigned((reg636 ? (8'haf) : reg636))} ?
                          reg619[(2'h3):(2'h3)] : forvar653[(4'hb):(2'h3)]);
                    end
                end
              reg688 <= reg660;
            end
          for (forvar689 = (1'h0); (forvar689 < (2'h2)); forvar689 = (forvar689 + (1'h1)))
            begin
              if ($signed(reg642[(4'hf):(1'h1)]))
                begin
                  if ($unsigned(reg645))
                    begin
                      reg690 <= forvar682;
                      reg691 <= (~^forvar682);
                      reg692 <= (reg635[(3'h6):(2'h2)] > (((+(8'h9f)) ?
                              ((8'hb2) ? reg686 : reg682) : $signed(wire616)) ?
                          $unsigned((forvar642 ?
                              forvar662 : reg684)) : ((reg645 ?
                                  wire617 : forvar621) ?
                              (wire612 ? reg631 : reg672) : ((8'h9e) ?
                                  reg685 : reg635))));
                      reg693 <= $unsigned($signed(reg672[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg690 <= (8'ha8);
                      reg691 <= reg660;
                    end
                end
              else
                begin
                  for (forvar690 = (1'h0); (forvar690 < (1'h0)); forvar690 = (forvar690 + (1'h1)))
                    begin
                      reg691 <= ($signed($unsigned(forvar622)) ?
                          $signed((((8'hb4) ^~ wire613) ?
                              $unsigned(forvar620) : (^~reg627))) : {{reg685[(2'h2):(1'h1)]}});
                      reg692 <= (({{wire614}} >> ((reg655 - (8'haf)) && {reg665})) ?
                          reg668[(1'h0):(1'h0)] : (reg658[(3'h6):(3'h4)] ?
                              (reg623[(2'h2):(2'h2)] ?
                                  reg643[(2'h2):(1'h1)] : {reg657}) : $unsigned($unsigned((8'hab)))));
                      reg693 <= reg684;
                    end
                  reg694 <= reg686[(4'h8):(1'h1)];
                  for (forvar695 = (1'h0); (forvar695 < (2'h3)); forvar695 = (forvar695 + (1'h1)))
                    begin
                      reg696 <= (reg672[(1'h1):(1'h1)] ?
                          (reg623 ?
                              $unsigned((reg656 >> (8'hac))) : reg665[(3'h6):(1'h0)]) : $signed(((^reg665) < reg628[(1'h0):(1'h0)])));
                    end
                end
              for (forvar697 = (1'h0); (forvar697 < (2'h3)); forvar697 = (forvar697 + (1'h1)))
                begin
                  for (forvar698 = (1'h0); (forvar698 < (1'h0)); forvar698 = (forvar698 + (1'h1)))
                    begin
                      reg699 <= {$signed($unsigned((wire617 != forvar677)))};
                      reg700 <= (reg654 >= reg663);
                      reg701 <= (~^(^~$signed($unsigned(reg623))));
                    end
                  if ({wire617[(4'h9):(3'h7)]})
                    begin
                      reg702 <= ((~^$signed(reg667[(1'h1):(1'h1)])) || $signed($unsigned({reg676})));
                    end
                  else
                    begin
                      reg702 <= (+((((8'haf) ?
                          forvar621 : reg674) | $unsigned(reg666)) - $signed((~^reg701))));
                      reg703 <= (-(8'ha7));
                      reg704 <= reg692;
                    end
                  reg705 <= forvar620;
                  reg706 <= (~reg694);
                end
            end
        end
      if (({$signed($signed(reg682))} || (8'hb5)))
        begin
          if (reg703)
            begin
              for (forvar707 = (1'h0); (forvar707 < (1'h0)); forvar707 = (forvar707 + (1'h1)))
                begin
                  reg708 <= (reg674[(2'h3):(2'h3)] <= $unsigned({$signed(forvar648)}));
                end
              for (forvar709 = (1'h0); (forvar709 < (2'h2)); forvar709 = (forvar709 + (1'h1)))
                begin
                  for (forvar710 = (1'h0); (forvar710 < (2'h3)); forvar710 = (forvar710 + (1'h1)))
                    begin
                      reg711 <= $unsigned($signed($signed((forvar621 ?
                          reg641 : reg679))));
                      reg712 <= $signed(((~&(wire617 ?
                          (8'ha2) : reg641)) != (~$signed((8'ha9)))));
                      reg713 <= $signed(reg703);
                    end
                end
            end
          else
            begin
              reg707 <= (reg642 || ($unsigned(reg639) ?
                  ((!reg622) ?
                      $signed(reg634) : reg667) : (((8'hb6) && reg630) | forvar664[(1'h1):(1'h0)])));
              for (forvar708 = (1'h0); (forvar708 < (1'h1)); forvar708 = (forvar708 + (1'h1)))
                begin
                  for (forvar709 = (1'h0); (forvar709 < (2'h2)); forvar709 = (forvar709 + (1'h1)))
                    begin
                      reg710 <= $unsigned(reg621);
                      reg711 <= $unsigned(((reg661 >>> reg656[(2'h2):(1'h0)]) && {(8'hac)}));
                    end
                  for (forvar712 = (1'h0); (forvar712 < (1'h1)); forvar712 = (forvar712 + (1'h1)))
                    begin
                      reg713 <= reg655[(2'h3):(2'h2)];
                      reg714 <= reg622[(2'h3):(1'h0)];
                      reg715 <= ((reg661 >>> $unsigned($signed((8'hba)))) ^~ reg632[(2'h3):(2'h3)]);
                    end
                  for (forvar716 = (1'h0); (forvar716 < (2'h2)); forvar716 = (forvar716 + (1'h1)))
                    begin
                      reg717 <= wire616;
                      reg718 <= $unsigned($unsigned((&$signed(reg714))));
                    end
                end
              if ((8'ha5))
                begin
                  if ($signed($unsigned({reg623})))
                    begin
                      reg719 <= reg654;
                      reg720 <= reg719[(3'h5):(1'h0)];
                      reg721 <= ((~((forvar653 <= reg642) >>> (reg644 ?
                          forvar641 : reg666))) - ($signed($unsigned(reg637)) ?
                          (((8'haf) ?
                              reg665 : (8'haa)) ~^ $signed((8'hba))) : $unsigned(reg644[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg719 <= (~^reg682);
                      reg720 <= (~&$signed($signed((reg679 | reg626))));
                      reg721 <= reg692[(4'hb):(4'ha)];
                      reg722 <= ($signed({(~|reg644)}) <= (|({reg636} >= reg644[(1'h0):(1'h0)])));
                    end
                  for (forvar723 = (1'h0); (forvar723 < (2'h3)); forvar723 = (forvar723 + (1'h1)))
                    begin
                      reg724 <= $signed($unsigned(reg640));
                      reg725 <= (^(($signed(wire612) == (forvar712 ?
                              forvar723 : reg672)) ?
                          forvar712[(1'h1):(1'h0)] : $signed((reg713 >= wire612))));
                      reg726 <= (((!$unsigned(reg693)) ?
                          $signed(reg635) : {$unsigned(reg713)}) >> ($signed((|(8'hab))) ?
                          $signed((|reg696)) : reg619[(2'h2):(1'h1)]));
                      reg727 <= forvar642[(3'h4):(3'h4)];
                    end
                  if ((8'ha6))
                    begin
                      reg728 <= ($signed((^(~&reg659))) > ($unsigned($signed(reg706)) ?
                          $signed((reg684 ?
                              (8'hac) : reg692)) : ((reg681 && reg725) ?
                              reg636[(3'h7):(1'h0)] : forvar620)));
                      reg729 <= ((forvar708[(1'h1):(1'h1)] ?
                          ($signed(reg694) ?
                              reg630 : (8'h9f)) : (~|$unsigned((8'ha6)))) + (^((~&reg711) ?
                          $unsigned(reg726) : $unsigned(reg708))));
                    end
                  else
                    begin
                      reg728 <= ($signed(reg678[(3'h4):(3'h4)]) <<< reg707[(4'h9):(2'h2)]);
                      reg729 <= ((~$signed(reg646)) == ((|{forvar629}) ~^ forvar621));
                      reg730 <= reg708;
                      reg731 <= wire613[(3'h4):(3'h4)];
                    end
                end
              else
                begin
                  if (reg628[(1'h0):(1'h0)])
                    begin
                      reg719 <= $unsigned(($unsigned((reg687 ?
                          reg730 : reg654)) | (reg667 ^~ $unsigned(reg647))));
                    end
                  else
                    begin
                      reg719 <= (reg685 ?
                          $signed((reg700[(4'hd):(2'h3)] ~^ (8'ha0))) : (((8'hb6) ~^ (reg659 <= (8'ha6))) ?
                              $signed(reg715[(2'h2):(1'h1)]) : (~^$unsigned(reg619))));
                      reg720 <= ($signed(((-reg681) * (^(8'ha9)))) ?
                          (-$signed(forvar620[(1'h1):(1'h0)])) : (reg660 ?
                              (8'hb0) : $unsigned({reg708})));
                      reg721 <= forvar681[(4'h9):(1'h1)];
                    end
                end
            end
          if ($unsigned((-(8'ha9))))
            begin
              reg732 <= (~&$unsigned($signed($unsigned(reg710))));
            end
          else
            begin
              for (forvar732 = (1'h0); (forvar732 < (1'h0)); forvar732 = (forvar732 + (1'h1)))
                begin
                  if ((((8'had) <<< $unsigned((-wire616))) || ($unsigned($unsigned(reg720)) ?
                      (~|(reg650 - reg624)) : $signed(forvar681[(2'h3):(1'h1)]))))
                    begin
                      reg733 <= ((~^reg651[(4'h9):(1'h0)]) ?
                          (((~(8'h9f)) ? $unsigned(reg700) : (8'h9c)) ?
                              reg658[(3'h6):(3'h6)] : reg708[(1'h0):(1'h0)]) : (reg731 ?
                              $unsigned((~^reg720)) : {(8'h9e)}));
                      reg734 <= reg729;
                    end
                  else
                    begin
                      reg733 <= reg636;
                    end
                end
              for (forvar735 = (1'h0); (forvar735 < (1'h1)); forvar735 = (forvar735 + (1'h1)))
                begin
                  for (forvar736 = (1'h0); (forvar736 < (1'h0)); forvar736 = (forvar736 + (1'h1)))
                    begin
                      reg737 <= ({reg651[(4'h8):(4'h8)]} ?
                          reg686[(4'hc):(3'h6)] : (!forvar716));
                    end
                end
              for (forvar738 = (1'h0); (forvar738 < (2'h2)); forvar738 = (forvar738 + (1'h1)))
                begin
                  for (forvar739 = (1'h0); (forvar739 < (1'h0)); forvar739 = (forvar739 + (1'h1)))
                    begin
                      reg740 <= $unsigned($signed((|$signed(reg687))));
                      reg741 <= forvar716;
                    end
                  for (forvar742 = (1'h0); (forvar742 < (1'h1)); forvar742 = (forvar742 + (1'h1)))
                    begin
                      reg743 <= $unsigned((wire613[(3'h5):(1'h0)] ?
                          ((-forvar618) ?
                              (^~forvar689) : (8'ha3)) : {reg721[(3'h7):(2'h3)]}));
                      reg744 <= (reg687[(3'h5):(2'h3)] ?
                          $signed($unsigned((~^reg658))) : ((reg630 ?
                              (~&reg676) : ((8'h9e) & reg733)) <= wire613));
                      reg745 <= $unsigned(forvar677[(3'h4):(1'h0)]);
                    end
                  if ($unsigned(forvar618[(3'h7):(3'h5)]))
                    begin
                      reg746 <= {$signed(reg650[(2'h3):(1'h1)])};
                      reg747 <= $signed({reg630});
                      reg748 <= (reg708 && ((((8'haa) * reg702) > forvar710) != {reg732[(1'h0):(1'h0)]}));
                    end
                  else
                    begin
                      reg746 <= $unsigned((reg676 | (&(reg722 * reg628))));
                      reg747 <= ((~({forvar742} ?
                          {forvar649} : ((8'hb2) ?
                              reg643 : wire614))) >>> ((reg733 ?
                          ((8'h9f) && reg706) : reg658[(3'h4):(1'h1)]) + {$signed((8'ha4))}));
                      reg748 <= ((~|($unsigned(wire617) < $signed(reg732))) ?
                          ($signed($unsigned(reg658)) * ($signed(reg682) ?
                              $signed(reg693) : (forvar723 || reg628))) : {(~reg701)});
                    end
                end
            end
          if (($unsigned((~reg684[(4'hb):(1'h0)])) - {reg717[(4'hd):(4'hb)]}))
            begin
              for (forvar749 = (1'h0); (forvar749 < (1'h1)); forvar749 = (forvar749 + (1'h1)))
                begin
                  for (forvar750 = (1'h0); (forvar750 < (2'h2)); forvar750 = (forvar750 + (1'h1)))
                    begin
                      reg751 <= {reg673};
                      reg752 <= (($signed($signed(reg751)) ?
                              (-{reg713}) : ($unsigned(reg672) <<< (|reg703))) ?
                          ((((8'ha9) ? reg663 : forvar736) ?
                              $signed(reg712) : reg685[(4'h9):(3'h7)]) ~^ $unsigned($signed((8'haa)))) : $unsigned($signed((~forvar620))));
                    end
                  reg753 <= forvar695[(4'h8):(1'h0)];
                  for (forvar754 = (1'h0); (forvar754 < (1'h1)); forvar754 = (forvar754 + (1'h1)))
                    begin
                      reg755 <= ((reg701 ?
                          $unsigned((8'h9d)) : reg672) * reg663[(1'h1):(1'h0)]);
                      reg756 <= (+(8'hb9));
                      reg757 <= (8'h9f);
                    end
                  if ((&($signed((reg659 ?
                      reg630 : reg743)) << reg757[(1'h0):(1'h0)])))
                    begin
                      reg758 <= $signed($signed((8'hb1)));
                      reg759 <= reg651[(4'hd):(4'h9)];
                      reg760 <= $signed(((^~(reg672 ? reg694 : (8'ha1))) ?
                          reg757 : reg641));
                      reg761 <= $signed($unsigned(((reg746 ?
                          reg643 : forvar750) == {reg686})));
                    end
                  else
                    begin
                      reg758 <= ($unsigned(forvar662[(1'h1):(1'h0)]) > (($unsigned(reg667) ?
                          forvar690 : ((8'hb6) && reg727)) << ((reg636 ?
                          reg725 : reg621) || {reg635})));
                      reg759 <= (+((~reg619) | reg680));
                      reg760 <= reg703;
                    end
                end
              reg762 <= {reg651};
              for (forvar763 = (1'h0); (forvar763 < (2'h2)); forvar763 = (forvar763 + (1'h1)))
                begin
                  for (forvar764 = (1'h0); (forvar764 < (1'h1)); forvar764 = (forvar764 + (1'h1)))
                    begin
                      reg765 <= $signed(forvar629);
                      reg766 <= (reg733[(2'h2):(1'h1)] == (({reg712} == (forvar663 ?
                              forvar625 : reg668)) ?
                          reg744[(2'h2):(1'h0)] : $unsigned((reg696 ?
                              (8'haf) : forvar653))));
                      reg767 <= (+(~|((reg668 >= forvar682) ?
                          (forvar709 ?
                              reg690 : (8'hb7)) : $unsigned(forvar710))));
                    end
                end
              if (reg647)
                begin
                  reg768 <= $signed((~&$signed((8'hb7))));
                end
              else
                begin
                  if (($signed({$signed(reg760)}) ?
                      {$signed({forvar712})} : $signed(($signed(reg744) ?
                          forvar675[(3'h5):(1'h1)] : (^~(8'ha7))))))
                    begin
                      reg768 <= (~&$unsigned({forvar649[(1'h1):(1'h0)]}));
                      reg769 <= reg753;
                    end
                  else
                    begin
                      reg768 <= $signed(((8'ha6) ^~ $signed(reg706)));
                      reg769 <= $unsigned(($unsigned($unsigned(forvar620)) + reg672[(2'h2):(2'h2)]));
                      reg770 <= ($signed($signed($unsigned(reg727))) | (($signed(reg745) ?
                          (|reg719) : (~(8'hb9))) && (forvar674 ^~ reg727[(2'h3):(2'h2)])));
                      reg771 <= reg740;
                    end
                  for (forvar772 = (1'h0); (forvar772 < (2'h3)); forvar772 = (forvar772 + (1'h1)))
                    begin
                      reg773 <= ((~&(~|forvar666[(3'h6):(2'h3)])) ?
                          reg757 : {$unsigned(reg751[(2'h3):(2'h2)])});
                      reg774 <= ((-$unsigned(forvar749[(2'h3):(2'h2)])) ?
                          $signed((8'ha8)) : reg664[(4'h9):(1'h0)]);
                      reg775 <= $signed(reg715);
                    end
                end
            end
          else
            begin
              for (forvar749 = (1'h0); (forvar749 < (1'h0)); forvar749 = (forvar749 + (1'h1)))
                begin
                  for (forvar750 = (1'h0); (forvar750 < (1'h1)); forvar750 = (forvar750 + (1'h1)))
                    begin
                      reg751 <= $signed(($unsigned(forvar673[(4'hb):(3'h5)]) * (reg681 ?
                          {(8'ha2)} : {(8'ha0)})));
                      reg752 <= $unsigned($signed(reg651));
                      reg753 <= $signed($signed(reg759));
                      reg754 <= $signed(reg675);
                    end
                end
            end
        end
      else
        begin
          for (forvar707 = (1'h0); (forvar707 < (1'h1)); forvar707 = (forvar707 + (1'h1)))
            begin
              if (($unsigned((^reg705[(3'h6):(2'h3)])) ?
                  {(~|((8'ha0) ?
                          reg720 : reg637))} : ({reg639[(4'h8):(3'h6)]} - (~&$signed(forvar677)))))
                begin
                  if (reg706)
                    begin
                      reg708 <= $unsigned({((8'hae) >>> forvar749[(4'ha):(3'h7)])});
                      reg709 <= (({forvar735} ?
                              ((reg708 ? reg717 : reg761) ?
                                  reg650[(3'h6):(1'h1)] : {forvar690}) : (^reg741)) ?
                          $unsigned(reg681[(3'h4):(3'h4)]) : ((~^(reg631 && reg627)) ?
                              (8'hb5) : ((+(8'h9f)) ?
                                  $signed(forvar669) : $unsigned(reg710))));
                      reg710 <= reg684[(4'hd):(4'h9)];
                      reg711 <= $signed(reg640);
                    end
                  else
                    begin
                      reg708 <= $unsigned({reg771});
                      reg709 <= $unsigned((~^((~forvar674) == $unsigned(forvar772))));
                      reg710 <= {reg668[(2'h3):(2'h3)]};
                    end
                  reg712 <= {($signed((forvar749 || reg732)) ?
                          $unsigned(forvar772[(3'h4):(2'h2)]) : (((8'ha3) ?
                                  reg719 : forvar735) ?
                              {reg624} : (^reg621)))};
                  if (($signed($unsigned(reg644)) && (reg771[(3'h4):(2'h2)] ?
                      (~{(8'hb0)}) : {(reg720 ~^ reg709)})))
                    begin
                      reg713 <= ($unsigned(((!reg770) * reg630)) * $signed({(reg724 ?
                              reg706 : reg638)}));
                      reg714 <= $signed($signed(forvar750));
                      reg715 <= $unsigned($unsigned((forvar677 ?
                          $unsigned(reg746) : $signed(reg743))));
                      reg716 <= ($unsigned($signed((8'hab))) >= (reg744[(1'h0):(1'h0)] <<< (reg634[(2'h2):(1'h0)] != (forvar669 ?
                          reg693 : (8'ha9)))));
                    end
                  else
                    begin
                      reg713 <= forvar675;
                      reg714 <= $unsigned(reg715);
                      reg715 <= forvar750[(3'h6):(3'h6)];
                    end
                end
              else
                begin
                  if ($unsigned($unsigned((|$unsigned(reg678)))))
                    begin
                      reg708 <= $signed((~$signed(reg632[(1'h0):(1'h0)])));
                      reg709 <= {(((^reg714) + {reg643}) ?
                              ((reg703 || reg758) >> reg655[(3'h5):(1'h0)]) : $signed((reg683 & forvar707)))};
                    end
                  else
                    begin
                      reg708 <= $signed((($signed(reg741) ?
                          forvar749[(3'h7):(2'h3)] : {forvar736}) * $signed(reg758[(1'h1):(1'h1)])));
                      reg709 <= reg645;
                    end
                  if ((~|$unsigned($unsigned(reg657))))
                    begin
                      reg710 <= (-(~&reg762));
                      reg711 <= {{((+forvar664) ~^ $signed(reg625))}};
                      reg712 <= reg733[(1'h1):(1'h1)];
                      reg713 <= reg711;
                    end
                  else
                    begin
                      reg710 <= (forvar754[(4'hc):(4'hb)] <= reg659[(3'h5):(3'h5)]);
                      reg711 <= ($unsigned(reg654[(2'h2):(2'h2)]) ?
                          ($signed((forvar754 ?
                              forvar723 : reg753)) & (reg700[(2'h2):(1'h1)] ~^ $unsigned(reg707))) : reg674);
                      reg712 <= reg682;
                      reg713 <= (((~|(8'hb2)) != reg711) ?
                          (reg625[(2'h2):(2'h2)] ?
                              ({reg687} ?
                                  reg746[(1'h1):(1'h0)] : $signed(reg756)) : (!wire614[(2'h2):(1'h0)])) : forvar642[(1'h1):(1'h1)]);
                    end
                  for (forvar714 = (1'h0); (forvar714 < (1'h1)); forvar714 = (forvar714 + (1'h1)))
                    begin
                      reg715 <= reg701;
                      reg716 <= (~(+reg700[(2'h2):(1'h0)]));
                      reg717 <= $unsigned(reg692);
                    end
                  for (forvar718 = (1'h0); (forvar718 < (2'h2)); forvar718 = (forvar718 + (1'h1)))
                    begin
                      reg719 <= $signed($signed(forvar750[(3'h5):(3'h4)]));
                      reg720 <= reg639;
                      reg721 <= $signed($unsigned((~^{forvar709})));
                    end
                end
            end
          for (forvar722 = (1'h0); (forvar722 < (2'h3)); forvar722 = (forvar722 + (1'h1)))
            begin
              for (forvar723 = (1'h0); (forvar723 < (1'h1)); forvar723 = (forvar723 + (1'h1)))
                begin
                  for (forvar724 = (1'h0); (forvar724 < (1'h0)); forvar724 = (forvar724 + (1'h1)))
                    begin
                      reg725 <= $signed($signed($signed((reg626 ^~ wire616))));
                      reg726 <= (!((+((8'hb6) || reg628)) >> {reg663[(3'h4):(1'h1)]}));
                      reg727 <= (~|(~|(forvar642 ? $signed((8'ha6)) : reg643)));
                      reg728 <= forvar708[(4'ha):(3'h7)];
                    end
                end
            end
        end
      for (forvar776 = (1'h0); (forvar776 < (1'h1)); forvar776 = (forvar776 + (1'h1)))
        begin
          reg777 <= forvar642;
        end
    end
  assign wire778 = {reg681};
  assign wire779 = $unsigned(reg666);
  assign wire780 = reg642;
  assign wire781 = reg679;
  always
    @(posedge clk) begin
      for (forvar782 = (1'h0); (forvar782 < (1'h1)); forvar782 = (forvar782 + (1'h1)))
        begin
          reg783 <= (reg645[(3'h4):(3'h4)] ?
              {((reg741 ?
                      reg674 : wire615) << $signed(reg707))} : ($unsigned((reg619 ?
                  reg635 : wire780)) == wire613));
          reg784 <= $unsigned(reg718[(3'h6):(3'h6)]);
          for (forvar785 = (1'h0); (forvar785 < (1'h1)); forvar785 = (forvar785 + (1'h1)))
            begin
              reg786 <= $unsigned($signed(reg753[(4'h8):(4'h8)]));
            end
        end
      reg787 <= (({(reg633 ? reg773 : reg747)} ? reg672 : {(reg729 + reg773)}) ?
          (reg652[(3'h5):(1'h0)] | reg680) : ($signed($signed(reg672)) | (((8'h9e) - reg725) && (reg674 ?
              reg771 : reg696))));
      if ({$signed($unsigned(reg666))})
        begin
          for (forvar788 = (1'h0); (forvar788 < (2'h3)); forvar788 = (forvar788 + (1'h1)))
            begin
              reg789 <= $unsigned({$unsigned((reg684 ? (8'ha0) : reg755))});
            end
          for (forvar790 = (1'h0); (forvar790 < (2'h2)); forvar790 = (forvar790 + (1'h1)))
            begin
              if (reg661)
                begin
                  for (forvar791 = (1'h0); (forvar791 < (2'h2)); forvar791 = (forvar791 + (1'h1)))
                    begin
                      reg792 <= (reg719 < $unsigned(wire780[(1'h0):(1'h0)]));
                      reg793 <= (-reg701[(3'h6):(1'h1)]);
                    end
                  if (reg622[(3'h4):(2'h3)])
                    begin
                      reg794 <= ((~^(^{reg757})) != (-($signed(reg657) ?
                          reg719[(4'h8):(1'h0)] : (~|reg773))));
                      reg795 <= ((~^$signed((reg667 >= (8'ha4)))) ?
                          reg707[(2'h3):(1'h1)] : reg756[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg794 <= {forvar791};
                    end
                  for (forvar796 = (1'h0); (forvar796 < (2'h2)); forvar796 = (forvar796 + (1'h1)))
                    begin
                      reg797 <= (-$unsigned((~$unsigned(wire612))));
                      reg798 <= reg769[(2'h2):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar791 = (1'h0); (forvar791 < (2'h2)); forvar791 = (forvar791 + (1'h1)))
                    begin
                      reg792 <= ($signed($signed($unsigned(reg789))) ?
                          $unsigned((~^{reg692})) : ((^(reg711 ?
                                  reg663 : reg729)) ?
                              (-$unsigned((8'hb4))) : $unsigned((|reg625))));
                      reg793 <= $signed(($unsigned(reg671[(4'hd):(2'h3)]) >> ({(8'ha9)} ~^ (~^reg702))));
                      reg794 <= (~reg760[(4'he):(2'h3)]);
                      reg795 <= (^$unsigned(($signed(wire617) > reg640[(1'h0):(1'h0)])));
                    end
                end
              if ($signed((8'ha6)))
                begin
                  for (forvar799 = (1'h0); (forvar799 < (1'h1)); forvar799 = (forvar799 + (1'h1)))
                    begin
                      reg800 <= {((~|(^reg632)) ?
                              (8'hb2) : $signed((&(8'h9c))))};
                      reg801 <= {(((wire780 ^~ forvar788) ?
                                  forvar785 : (wire612 >= reg646)) ?
                              reg767[(2'h2):(2'h2)] : (~(~|(8'ha8))))};
                      reg802 <= (reg740 ?
                          $signed($unsigned((forvar791 ?
                              reg623 : reg793))) : reg718[(1'h0):(1'h0)]);
                    end
                  reg803 <= $signed({$signed((reg733 ~^ reg626))});
                  for (forvar804 = (1'h0); (forvar804 < (1'h1)); forvar804 = (forvar804 + (1'h1)))
                    begin
                      reg805 <= ((reg794 - {$signed(reg752)}) != reg692[(1'h1):(1'h1)]);
                    end
                  for (forvar806 = (1'h0); (forvar806 < (1'h0)); forvar806 = (forvar806 + (1'h1)))
                    begin
                      reg807 <= (~|reg712);
                    end
                end
              else
                begin
                  if (reg730)
                    begin
                      reg799 <= reg663[(1'h1):(1'h1)];
                      reg800 <= (^((reg758[(3'h6):(3'h4)] ?
                          reg694 : $unsigned((8'had))) * ($signed(reg655) ?
                          reg755[(3'h6):(3'h4)] : (reg655 ?
                              (8'h9c) : reg740))));
                      reg801 <= (-reg761[(2'h2):(1'h1)]);
                      reg802 <= ((((forvar799 ? (8'hb2) : reg722) ?
                          (~&reg673) : (reg766 || (8'hb4))) == reg762[(4'h9):(3'h4)]) & $unsigned($unsigned((reg664 >= reg799))));
                    end
                  else
                    begin
                      reg799 <= (|$signed(wire779));
                    end
                  reg803 <= $unsigned((~^(|(reg795 - reg798))));
                  if ((($unsigned(reg702) > reg774[(2'h2):(1'h0)]) == (8'hae)))
                    begin
                      reg804 <= ((($unsigned(reg730) == $unsigned(wire778)) | reg798) << (reg752 << ((reg711 ~^ reg650) >>> {reg727})));
                      reg805 <= $unsigned($signed(reg667));
                    end
                  else
                    begin
                      reg804 <= reg802[(2'h3):(2'h2)];
                      reg805 <= reg800[(2'h3):(1'h1)];
                      reg806 <= wire615;
                      reg807 <= (+reg804[(4'h9):(3'h4)]);
                    end
                end
              for (forvar808 = (1'h0); (forvar808 < (1'h1)); forvar808 = (forvar808 + (1'h1)))
                begin
                  if ((reg792 ?
                      {$signed(reg671[(3'h6):(3'h4)])} : $unsigned((|$unsigned((8'hb1))))))
                    begin
                      reg809 <= $signed({({reg733} | (forvar790 || reg758))});
                      reg810 <= (+$signed(((^~reg658) ? (8'hb9) : {reg679})));
                      reg811 <= $signed($unsigned($signed(reg666)));
                    end
                  else
                    begin
                      reg809 <= $signed(reg766);
                      reg810 <= (|forvar790);
                    end
                  for (forvar812 = (1'h0); (forvar812 < (1'h1)); forvar812 = (forvar812 + (1'h1)))
                    begin
                      reg813 <= (8'hb9);
                      reg814 <= ($unsigned(reg703[(2'h2):(1'h0)]) ?
                          $signed(reg711) : $signed(reg767[(1'h0):(1'h0)]));
                    end
                end
              for (forvar815 = (1'h0); (forvar815 < (2'h2)); forvar815 = (forvar815 + (1'h1)))
                begin
                  for (forvar816 = (1'h0); (forvar816 < (2'h3)); forvar816 = (forvar816 + (1'h1)))
                    begin
                      reg817 <= $unsigned($signed($signed(reg783)));
                      reg818 <= (^reg775[(3'h6):(2'h2)]);
                      reg819 <= $unsigned($signed(reg753[(3'h4):(1'h0)]));
                    end
                end
            end
        end
      else
        begin
          reg788 <= reg708[(4'ha):(4'h8)];
        end
    end
  assign wire820 = reg718;
  assign wire821 = $unsigned(($unsigned($signed(reg641)) ^ ((reg678 <<< reg755) + ((8'ha6) + reg641))));
  assign wire822 = reg733;
  assign wire823 = (($unsigned(reg751[(5'h10):(4'hc)]) ?
                           reg717 : (^(^~reg800))) ?
                       ((!((8'hb7) < reg690)) | wire820[(2'h3):(1'h1)]) : (~&(-(reg621 ?
                           (8'hb2) : reg809))));
  assign wire824 = {{reg729}};
  assign wire825 = ({((reg728 >> reg642) ? {wire780} : $signed((8'haa)))} ?
                       reg682 : {reg664[(1'h0):(1'h0)]});
  assign wire826 = wire778;
  assign wire827 = $signed(($unsigned(reg753[(4'h8):(2'h2)]) << (-$unsigned(reg814))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module157  (y, clk, wire161, wire160, wire159, wire158);
  output wire [(32'h60):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire161;
  input wire signed [(4'h9):(1'h0)] wire160;
  input wire signed [(4'h9):(1'h0)] wire159;
  input wire signed [(2'h3):(1'h0)] wire158;
  wire [(4'hc):(1'h0)] wire170;
  wire [(3'h4):(1'h0)] wire169;
  wire signed [(4'hc):(1'h0)] wire168;
  wire signed [(3'h5):(1'h0)] wire167;
  wire signed [(3'h7):(1'h0)] wire166;
  wire [(4'hc):(1'h0)] wire165;
  wire [(4'hd):(1'h0)] wire164;
  wire [(4'he):(1'h0)] wire163;
  wire [(5'h10):(1'h0)] wire162;
  assign y = {wire170,
                 wire169,
                 wire168,
                 wire167,
                 wire166,
                 wire165,
                 wire164,
                 wire163,
                 wire162,
                 (1'h0)};
  assign wire162 = $signed({((wire161 ^ (8'ha5)) >> (8'hb9))});
  assign wire163 = (~$unsigned((8'ha3)));
  assign wire164 = $unsigned($unsigned(($signed(wire163) >> wire160)));
  assign wire165 = wire162[(2'h2):(1'h0)];
  assign wire166 = $signed((wire164[(3'h6):(1'h0)] && $unsigned($unsigned(wire165))));
  assign wire167 = (^({(wire164 <<< (8'hb1))} ?
                       ((!wire165) > (~&wire165)) : ($unsigned(wire160) ?
                           $unsigned(wire158) : $signed((8'ha2)))));
  assign wire168 = (~^wire160[(1'h1):(1'h0)]);
  assign wire169 = (((^(8'hb6)) && wire168[(2'h3):(1'h1)]) || wire160);
  assign wire170 = {{(-(wire168 ^~ wire166))}};
endmodule