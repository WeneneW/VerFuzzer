(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param4726 = ((((|(8'ha7)) ^ (&(8'hab))) ? (~^((8'hb7) == (8'hb1))) : (^~((8'hb4) ? (8'ha2) : (8'hb1)))) ~^ {(((8'hb8) ? (8'ha2) : (8'ha5)) << ((8'hb4) ? (8'ha3) : (8'h9f)))}))
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h26):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire0;
  input wire [(5'h10):(1'h0)] wire1;
  input wire [(4'he):(1'h0)] wire2;
  input wire [(4'hf):(1'h0)] wire3;
  wire signed [(3'h5):(1'h0)] wire4725;
  wire [(3'h4):(1'h0)] wire4724;
  wire [(4'hd):(1'h0)] wire4;
  wire signed [(2'h3):(1'h0)] wire3405;
  wire signed [(4'hc):(1'h0)] wire4722;
  assign y = {wire4725, wire4724, wire4, wire3405, wire4722, (1'h0)};
  assign wire4 = ((+wire2[(4'h8):(3'h5)]) ? $signed(wire3) : {wire3});
  module5 #() modinst3406 (.wire6(wire2), .wire8(wire0), .wire7(wire1), .clk(clk), .y(wire3405), .wire9(wire3));
  module3407 #() modinst4723 (.wire3408(wire2), .wire3409(wire3), .wire3410(wire1), .wire3411(wire4), .y(wire4722), .clk(clk), .wire3412(wire0));
  assign wire4724 = $signed($signed((8'hac)));
  assign wire4725 = ((~^$signed({wire0})) ?
                        ((|(wire4724 ? wire4722 : wire2)) + wire4722) : wire1);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3407
#(parameter param4721 = (~(^~(|((8'h9f) ^~ (8'hab))))))
(y, clk, wire3412, wire3411, wire3410, wire3409, wire3408);
  output wire [(32'h2a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire3412;
  input wire signed [(3'h4):(1'h0)] wire3411;
  input wire signed [(5'h10):(1'h0)] wire3410;
  input wire signed [(4'hf):(1'h0)] wire3409;
  input wire signed [(4'hc):(1'h0)] wire3408;
  wire signed [(4'hf):(1'h0)] wire3898;
  wire signed [(4'hf):(1'h0)] wire3413;
  wire signed [(3'h6):(1'h0)] wire3900;
  wire signed [(3'h5):(1'h0)] wire4719;
  assign y = {wire3898, wire3413, wire3900, wire4719, (1'h0)};
  assign wire3413 = ((wire3408 ?
                        wire3411[(1'h0):(1'h0)] : wire3408) ~^ $signed(wire3412));
  module3414 #() modinst3899 (.wire3416(wire3410), .clk(clk), .y(wire3898), .wire3417(wire3408), .wire3419(wire3409), .wire3418(wire3412), .wire3415(wire3413));
  assign wire3900 = wire3412;
  module3901 #() modinst4720 (wire4719, clk, wire3900, wire3409, wire3411, wire3898, wire3408);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module5
#(parameter param3404 = ({(((8'ha3) ? (8'hb6) : (8'hb8)) | (!(8'ha3)))} ? ((((8'ha4) && (8'h9d)) <<< ((8'had) ? (8'hb4) : (8'ha7))) ? ({(8'hb2)} ^ ((8'ha0) ? (8'ha3) : (8'ha1))) : (((8'hb5) ^~ (8'hb6)) ? ((8'hb8) ^~ (8'h9f)) : ((8'h9f) ? (8'h9d) : (8'ha4)))) : (~&(8'ha2))))
(y, clk, wire9, wire8, wire7, wire6);
  output wire [(32'h265d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire9;
  input wire [(3'h4):(1'h0)] wire8;
  input wire [(4'hc):(1'h0)] wire7;
  input wire [(4'he):(1'h0)] wire6;
  wire signed [(2'h2):(1'h0)] wire3402;
  wire [(4'h8):(1'h0)] wire1179;
  wire signed [(5'h10):(1'h0)] wire1040;
  wire [(3'h5):(1'h0)] wire964;
  wire [(3'h7):(1'h0)] wire708;
  wire signed [(4'h9):(1'h0)] wire707;
  wire [(4'hf):(1'h0)] wire492;
  reg signed [(4'ha):(1'h0)] reg1176 = (1'h0);
  reg [(4'h8):(1'h0)] reg1167 = (1'h0);
  reg [(4'h9):(1'h0)] reg1178 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1177 = (1'h0);
  reg [(4'hb):(1'h0)] reg1175 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1174 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1173 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1172 = (1'h0);
  reg [(3'h5):(1'h0)] reg1170 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1169 = (1'h0);
  reg [(3'h6):(1'h0)] reg1168 = (1'h0);
  reg [(3'h5):(1'h0)] reg1145 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1165 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1164 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1163 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1161 = (1'h0);
  reg [(2'h3):(1'h0)] reg1160 = (1'h0);
  reg [(3'h7):(1'h0)] reg1159 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1158 = (1'h0);
  reg [(4'h8):(1'h0)] reg1157 = (1'h0);
  reg [(4'hc):(1'h0)] reg1156 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1155 = (1'h0);
  reg [(4'ha):(1'h0)] reg1154 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1153 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1152 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1151 = (1'h0);
  reg [(2'h2):(1'h0)] reg1150 = (1'h0);
  reg [(4'h9):(1'h0)] reg1149 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1148 = (1'h0);
  reg [(4'hc):(1'h0)] reg1147 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1146 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1133 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1143 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1142 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1141 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1140 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1138 = (1'h0);
  reg [(4'h8):(1'h0)] reg1137 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1136 = (1'h0);
  reg [(4'hd):(1'h0)] reg1135 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1134 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1132 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1125 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1131 = (1'h0);
  reg [(4'hf):(1'h0)] reg1130 = (1'h0);
  reg [(4'hd):(1'h0)] reg1129 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1128 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1127 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1126 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1124 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1123 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1122 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1120 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1119 = (1'h0);
  reg [(3'h7):(1'h0)] reg1118 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1116 = (1'h0);
  reg [(4'h8):(1'h0)] reg1113 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1115 = (1'h0);
  reg [(5'h10):(1'h0)] reg1114 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1112 = (1'h0);
  reg [(3'h7):(1'h0)] reg1111 = (1'h0);
  reg [(4'hd):(1'h0)] reg1110 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1109 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1108 = (1'h0);
  reg [(3'h6):(1'h0)] reg1107 = (1'h0);
  reg [(4'hb):(1'h0)] reg1106 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1105 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1104 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1103 = (1'h0);
  reg [(3'h4):(1'h0)] reg1102 = (1'h0);
  reg [(4'ha):(1'h0)] reg1101 = (1'h0);
  reg [(4'h9):(1'h0)] reg1090 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1099 = (1'h0);
  reg [(3'h5):(1'h0)] reg1097 = (1'h0);
  reg [(4'he):(1'h0)] reg1096 = (1'h0);
  reg [(4'hd):(1'h0)] reg1095 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1094 = (1'h0);
  reg [(4'hd):(1'h0)] reg1093 = (1'h0);
  reg [(4'hf):(1'h0)] reg1092 = (1'h0);
  reg [(5'h10):(1'h0)] reg1091 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1089 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1088 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1087 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1086 = (1'h0);
  reg [(5'h10):(1'h0)] reg1085 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1084 = (1'h0);
  reg [(4'h8):(1'h0)] reg1082 = (1'h0);
  reg [(3'h5):(1'h0)] reg1081 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1080 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1079 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1076 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1075 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1073 = (1'h0);
  reg [(4'hf):(1'h0)] reg1072 = (1'h0);
  reg [(5'h10):(1'h0)] reg1071 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1070 = (1'h0);
  reg [(3'h6):(1'h0)] reg1069 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1065 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1064 = (1'h0);
  reg [(3'h4):(1'h0)] reg1045 = (1'h0);
  reg [(3'h4):(1'h0)] reg1042 = (1'h0);
  reg [(4'ha):(1'h0)] reg1062 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1061 = (1'h0);
  reg [(5'h10):(1'h0)] reg1060 = (1'h0);
  reg [(3'h6):(1'h0)] reg1059 = (1'h0);
  reg [(4'hc):(1'h0)] reg1058 = (1'h0);
  reg [(4'hb):(1'h0)] reg1057 = (1'h0);
  reg [(3'h5):(1'h0)] reg1056 = (1'h0);
  reg [(2'h3):(1'h0)] reg1055 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1053 = (1'h0);
  reg [(2'h3):(1'h0)] reg1052 = (1'h0);
  reg [(2'h3):(1'h0)] reg1051 = (1'h0);
  reg [(4'h8):(1'h0)] reg1046 = (1'h0);
  reg [(2'h3):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1049 = (1'h0);
  reg [(2'h3):(1'h0)] reg1048 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1047 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1044 = (1'h0);
  reg [(4'hb):(1'h0)] reg1043 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1041 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1039 = (1'h0);
  reg [(3'h6):(1'h0)] reg1037 = (1'h0);
  reg [(3'h4):(1'h0)] reg1036 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1035 = (1'h0);
  reg [(4'hb):(1'h0)] reg1034 = (1'h0);
  reg [(3'h7):(1'h0)] reg1031 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1030 = (1'h0);
  reg [(4'hd):(1'h0)] reg1029 = (1'h0);
  reg [(3'h6):(1'h0)] reg1027 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1026 = (1'h0);
  reg [(5'h10):(1'h0)] reg1025 = (1'h0);
  reg [(2'h2):(1'h0)] reg1024 = (1'h0);
  reg [(4'h9):(1'h0)] reg1023 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1022 = (1'h0);
  reg [(4'h9):(1'h0)] reg1021 = (1'h0);
  reg [(4'h8):(1'h0)] reg1020 = (1'h0);
  reg [(3'h4):(1'h0)] reg1019 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1018 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1017 = (1'h0);
  reg [(3'h4):(1'h0)] reg1011 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1016 = (1'h0);
  reg [(3'h6):(1'h0)] reg1015 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1013 = (1'h0);
  reg [(4'ha):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1010 = (1'h0);
  reg [(4'hd):(1'h0)] reg1009 = (1'h0);
  reg [(4'h9):(1'h0)] reg1008 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1007 = (1'h0);
  reg [(4'h8):(1'h0)] reg993 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1004 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1003 = (1'h0);
  reg [(4'h9):(1'h0)] reg1002 = (1'h0);
  reg [(4'hb):(1'h0)] reg1001 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1000 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg999 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg998 = (1'h0);
  reg [(2'h2):(1'h0)] reg997 = (1'h0);
  reg [(5'h10):(1'h0)] reg995 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg994 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg992 = (1'h0);
  reg [(4'hc):(1'h0)] reg991 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg979 = (1'h0);
  reg [(2'h3):(1'h0)] reg986 = (1'h0);
  reg [(4'h8):(1'h0)] reg981 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg974 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg990 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg989 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg988 = (1'h0);
  reg [(4'h9):(1'h0)] reg987 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg985 = (1'h0);
  reg [(3'h6):(1'h0)] reg984 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg983 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg982 = (1'h0);
  reg [(3'h7):(1'h0)] reg980 = (1'h0);
  reg signed [(4'he):(1'h0)] reg969 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg978 = (1'h0);
  reg [(3'h7):(1'h0)] reg977 = (1'h0);
  reg [(4'hc):(1'h0)] reg976 = (1'h0);
  reg [(4'ha):(1'h0)] reg975 = (1'h0);
  reg [(2'h2):(1'h0)] reg973 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg972 = (1'h0);
  reg [(4'ha):(1'h0)] reg971 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg970 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg968 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg967 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg966 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg965 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg963 = (1'h0);
  reg [(4'hd):(1'h0)] reg962 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg961 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg960 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg959 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg958 = (1'h0);
  reg [(4'hf):(1'h0)] reg956 = (1'h0);
  reg [(4'ha):(1'h0)] reg953 = (1'h0);
  reg [(2'h3):(1'h0)] reg952 = (1'h0);
  reg [(4'ha):(1'h0)] reg949 = (1'h0);
  reg [(3'h6):(1'h0)] reg947 = (1'h0);
  reg [(2'h3):(1'h0)] reg946 = (1'h0);
  reg [(4'ha):(1'h0)] reg945 = (1'h0);
  reg [(2'h3):(1'h0)] reg943 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg942 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg932 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg930 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg940 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg939 = (1'h0);
  reg [(4'h8):(1'h0)] reg938 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg937 = (1'h0);
  reg [(4'hb):(1'h0)] reg935 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg934 = (1'h0);
  reg [(3'h6):(1'h0)] reg933 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg931 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg929 = (1'h0);
  reg [(4'hc):(1'h0)] reg928 = (1'h0);
  reg signed [(4'he):(1'h0)] reg927 = (1'h0);
  reg [(3'h6):(1'h0)] reg926 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg925 = (1'h0);
  reg [(3'h6):(1'h0)] reg924 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg923 = (1'h0);
  reg [(4'hc):(1'h0)] reg922 = (1'h0);
  reg [(4'hc):(1'h0)] reg921 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg920 = (1'h0);
  reg signed [(4'he):(1'h0)] reg919 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg918 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg917 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg916 = (1'h0);
  reg [(4'ha):(1'h0)] reg915 = (1'h0);
  reg [(3'h7):(1'h0)] reg913 = (1'h0);
  reg [(2'h3):(1'h0)] reg912 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg908 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg907 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg906 = (1'h0);
  reg [(3'h4):(1'h0)] reg905 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg903 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg902 = (1'h0);
  reg [(3'h6):(1'h0)] reg901 = (1'h0);
  reg [(4'hf):(1'h0)] reg898 = (1'h0);
  reg [(4'hf):(1'h0)] reg897 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg896 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg895 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg893 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg892 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg890 = (1'h0);
  reg [(4'hf):(1'h0)] reg891 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg889 = (1'h0);
  reg [(4'h9):(1'h0)] reg888 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg887 = (1'h0);
  reg [(4'hb):(1'h0)] reg883 = (1'h0);
  reg [(4'ha):(1'h0)] reg882 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg881 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg880 = (1'h0);
  reg [(2'h3):(1'h0)] reg879 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg877 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg875 = (1'h0);
  reg [(4'hf):(1'h0)] reg874 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg873 = (1'h0);
  reg [(4'h8):(1'h0)] reg872 = (1'h0);
  reg [(5'h10):(1'h0)] reg871 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg868 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg867 = (1'h0);
  reg [(2'h3):(1'h0)] reg866 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg865 = (1'h0);
  reg [(4'he):(1'h0)] reg864 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg862 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg861 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg860 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg859 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg858 = (1'h0);
  reg [(5'h10):(1'h0)] reg857 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg856 = (1'h0);
  reg signed [(4'he):(1'h0)] reg855 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg854 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg853 = (1'h0);
  reg [(4'ha):(1'h0)] reg852 = (1'h0);
  reg [(4'h9):(1'h0)] reg850 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg849 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg847 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg846 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg845 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg843 = (1'h0);
  reg signed [(4'he):(1'h0)] reg842 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg841 = (1'h0);
  reg [(3'h6):(1'h0)] reg840 = (1'h0);
  reg [(4'hc):(1'h0)] reg839 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg838 = (1'h0);
  reg [(4'hc):(1'h0)] reg837 = (1'h0);
  reg [(5'h10):(1'h0)] reg836 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg835 = (1'h0);
  reg [(3'h5):(1'h0)] reg834 = (1'h0);
  reg [(4'ha):(1'h0)] reg833 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg832 = (1'h0);
  reg [(4'ha):(1'h0)] reg831 = (1'h0);
  reg [(2'h2):(1'h0)] reg830 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg829 = (1'h0);
  reg [(3'h6):(1'h0)] reg828 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg783 = (1'h0);
  reg [(4'he):(1'h0)] reg824 = (1'h0);
  reg [(4'hc):(1'h0)] reg823 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg822 = (1'h0);
  reg [(4'he):(1'h0)] reg821 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg820 = (1'h0);
  reg [(5'h10):(1'h0)] reg819 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg818 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg817 = (1'h0);
  reg [(4'hb):(1'h0)] reg816 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg815 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg814 = (1'h0);
  reg [(4'he):(1'h0)] reg813 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg793 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg798 = (1'h0);
  reg [(4'he):(1'h0)] reg796 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg811 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg808 = (1'h0);
  reg [(4'h9):(1'h0)] reg807 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg806 = (1'h0);
  reg [(4'ha):(1'h0)] reg805 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg804 = (1'h0);
  reg signed [(4'he):(1'h0)] reg803 = (1'h0);
  reg [(2'h3):(1'h0)] reg802 = (1'h0);
  reg [(4'h9):(1'h0)] reg801 = (1'h0);
  reg [(3'h6):(1'h0)] reg800 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg799 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg797 = (1'h0);
  reg [(2'h3):(1'h0)] reg795 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg794 = (1'h0);
  reg [(4'h8):(1'h0)] reg792 = (1'h0);
  reg [(4'hc):(1'h0)] reg791 = (1'h0);
  reg [(5'h10):(1'h0)] reg790 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg789 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg788 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg785 = (1'h0);
  reg [(4'h8):(1'h0)] reg787 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg786 = (1'h0);
  reg [(4'h8):(1'h0)] reg784 = (1'h0);
  reg [(5'h10):(1'h0)] reg782 = (1'h0);
  reg [(2'h3):(1'h0)] reg781 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg780 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg779 = (1'h0);
  reg [(4'hb):(1'h0)] reg775 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg774 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg773 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg772 = (1'h0);
  reg [(3'h7):(1'h0)] reg768 = (1'h0);
  reg [(4'h9):(1'h0)] reg771 = (1'h0);
  reg [(2'h3):(1'h0)] reg770 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg769 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg762 = (1'h0);
  reg [(2'h3):(1'h0)] reg756 = (1'h0);
  reg [(4'h9):(1'h0)] reg767 = (1'h0);
  reg [(3'h5):(1'h0)] reg766 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg765 = (1'h0);
  reg [(5'h10):(1'h0)] reg764 = (1'h0);
  reg [(4'hf):(1'h0)] reg763 = (1'h0);
  reg [(3'h5):(1'h0)] reg761 = (1'h0);
  reg [(4'ha):(1'h0)] reg760 = (1'h0);
  reg [(2'h2):(1'h0)] reg759 = (1'h0);
  reg [(4'hb):(1'h0)] reg758 = (1'h0);
  reg [(4'h9):(1'h0)] reg757 = (1'h0);
  reg [(4'h8):(1'h0)] reg753 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg748 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg746 = (1'h0);
  reg [(3'h6):(1'h0)] reg745 = (1'h0);
  reg [(3'h7):(1'h0)] reg737 = (1'h0);
  reg [(4'hc):(1'h0)] reg732 = (1'h0);
  reg [(4'h8):(1'h0)] reg714 = (1'h0);
  reg [(4'he):(1'h0)] reg755 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg754 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg752 = (1'h0);
  reg signed [(4'he):(1'h0)] reg751 = (1'h0);
  reg [(4'he):(1'h0)] reg750 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg749 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg747 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg744 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg743 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg742 = (1'h0);
  reg [(3'h7):(1'h0)] reg741 = (1'h0);
  reg [(4'hf):(1'h0)] reg740 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg739 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg738 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg735 = (1'h0);
  reg [(3'h7):(1'h0)] reg734 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg733 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg731 = (1'h0);
  reg signed [(4'he):(1'h0)] reg730 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg729 = (1'h0);
  reg [(4'hb):(1'h0)] reg728 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg727 = (1'h0);
  reg [(3'h6):(1'h0)] reg720 = (1'h0);
  reg [(4'hf):(1'h0)] reg722 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg726 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg725 = (1'h0);
  reg [(4'he):(1'h0)] reg724 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg723 = (1'h0);
  reg [(4'hf):(1'h0)] reg721 = (1'h0);
  reg [(4'hc):(1'h0)] reg719 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg718 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg717 = (1'h0);
  reg [(4'he):(1'h0)] reg716 = (1'h0);
  reg [(3'h6):(1'h0)] reg715 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg713 = (1'h0);
  reg [(4'hb):(1'h0)] reg712 = (1'h0);
  reg [(4'hb):(1'h0)] reg711 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg710 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg709 = (1'h0);
  reg [(2'h3):(1'h0)] reg706 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg705 = (1'h0);
  reg [(4'hd):(1'h0)] reg704 = (1'h0);
  reg [(4'hf):(1'h0)] reg701 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg698 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg697 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg685 = (1'h0);
  reg signed [(4'he):(1'h0)] reg702 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg700 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg699 = (1'h0);
  reg [(4'h8):(1'h0)] reg696 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg695 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg694 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg693 = (1'h0);
  reg [(2'h3):(1'h0)] reg692 = (1'h0);
  reg [(3'h5):(1'h0)] reg691 = (1'h0);
  reg [(3'h5):(1'h0)] reg690 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg689 = (1'h0);
  reg [(3'h5):(1'h0)] reg688 = (1'h0);
  reg [(4'hf):(1'h0)] reg687 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg686 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg684 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg683 = (1'h0);
  reg [(2'h2):(1'h0)] reg682 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg681 = (1'h0);
  reg [(4'hb):(1'h0)] reg680 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg679 = (1'h0);
  reg [(3'h4):(1'h0)] reg678 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg677 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg675 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg674 = (1'h0);
  reg signed [(4'he):(1'h0)] reg673 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg668 = (1'h0);
  reg signed [(4'he):(1'h0)] reg672 = (1'h0);
  reg signed [(4'he):(1'h0)] reg671 = (1'h0);
  reg [(4'he):(1'h0)] reg670 = (1'h0);
  reg [(2'h3):(1'h0)] reg669 = (1'h0);
  reg [(3'h5):(1'h0)] reg667 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg666 = (1'h0);
  reg [(2'h2):(1'h0)] reg665 = (1'h0);
  reg [(4'hf):(1'h0)] reg660 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg655 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg664 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg663 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg662 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg661 = (1'h0);
  reg [(4'ha):(1'h0)] reg659 = (1'h0);
  reg [(3'h4):(1'h0)] reg658 = (1'h0);
  reg [(4'hd):(1'h0)] reg657 = (1'h0);
  reg [(4'he):(1'h0)] reg656 = (1'h0);
  reg [(4'he):(1'h0)] reg651 = (1'h0);
  reg [(3'h5):(1'h0)] reg636 = (1'h0);
  reg [(2'h2):(1'h0)] reg654 = (1'h0);
  reg [(3'h6):(1'h0)] reg653 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg652 = (1'h0);
  reg signed [(4'he):(1'h0)] reg650 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg649 = (1'h0);
  reg [(4'hb):(1'h0)] reg648 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg647 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg646 = (1'h0);
  reg [(4'ha):(1'h0)] reg645 = (1'h0);
  reg [(2'h2):(1'h0)] reg644 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg643 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg642 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg641 = (1'h0);
  reg [(2'h3):(1'h0)] reg639 = (1'h0);
  reg [(4'hc):(1'h0)] reg638 = (1'h0);
  reg [(4'hc):(1'h0)] reg637 = (1'h0);
  reg [(3'h5):(1'h0)] reg635 = (1'h0);
  reg [(4'hc):(1'h0)] reg614 = (1'h0);
  reg [(3'h4):(1'h0)] reg634 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg633 = (1'h0);
  reg [(4'h8):(1'h0)] reg631 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg630 = (1'h0);
  reg signed [(4'he):(1'h0)] reg629 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg628 = (1'h0);
  reg [(2'h2):(1'h0)] reg627 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg626 = (1'h0);
  reg [(2'h2):(1'h0)] reg624 = (1'h0);
  reg [(4'hf):(1'h0)] reg623 = (1'h0);
  reg [(2'h3):(1'h0)] reg622 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg621 = (1'h0);
  reg [(2'h3):(1'h0)] reg618 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg617 = (1'h0);
  reg [(4'he):(1'h0)] reg616 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg615 = (1'h0);
  reg [(4'hb):(1'h0)] reg587 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg598 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg613 = (1'h0);
  reg [(2'h2):(1'h0)] reg612 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg610 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg609 = (1'h0);
  reg [(4'hb):(1'h0)] reg608 = (1'h0);
  reg [(3'h7):(1'h0)] reg606 = (1'h0);
  reg [(4'hd):(1'h0)] reg599 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg586 = (1'h0);
  reg signed [(4'he):(1'h0)] reg605 = (1'h0);
  reg [(4'ha):(1'h0)] reg604 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg603 = (1'h0);
  reg [(4'hc):(1'h0)] reg602 = (1'h0);
  reg [(4'h9):(1'h0)] reg601 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg600 = (1'h0);
  reg [(4'ha):(1'h0)] reg597 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg596 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg595 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg594 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg593 = (1'h0);
  reg [(3'h5):(1'h0)] reg592 = (1'h0);
  reg [(2'h2):(1'h0)] reg591 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg590 = (1'h0);
  reg signed [(4'he):(1'h0)] reg589 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg588 = (1'h0);
  reg [(2'h2):(1'h0)] reg585 = (1'h0);
  reg [(3'h7):(1'h0)] reg584 = (1'h0);
  reg [(4'hb):(1'h0)] reg583 = (1'h0);
  reg signed [(4'he):(1'h0)] reg578 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg573 = (1'h0);
  reg signed [(4'he):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg581 = (1'h0);
  reg [(4'hb):(1'h0)] reg580 = (1'h0);
  reg [(3'h5):(1'h0)] reg579 = (1'h0);
  reg [(2'h2):(1'h0)] reg577 = (1'h0);
  reg [(4'ha):(1'h0)] reg576 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg575 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg574 = (1'h0);
  reg [(4'hc):(1'h0)] reg571 = (1'h0);
  reg [(3'h6):(1'h0)] reg525 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg516 = (1'h0);
  reg [(2'h3):(1'h0)] reg514 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg526 = (1'h0);
  reg [(3'h4):(1'h0)] reg517 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg509 = (1'h0);
  reg [(4'ha):(1'h0)] reg501 = (1'h0);
  reg [(4'hd):(1'h0)] reg500 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg545 = (1'h0);
  reg [(3'h4):(1'h0)] reg542 = (1'h0);
  reg [(5'h10):(1'h0)] reg541 = (1'h0);
  reg [(4'he):(1'h0)] reg570 = (1'h0);
  reg [(4'he):(1'h0)] reg569 = (1'h0);
  reg [(2'h3):(1'h0)] reg568 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg567 = (1'h0);
  reg [(3'h7):(1'h0)] reg566 = (1'h0);
  reg [(4'h9):(1'h0)] reg565 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg564 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg563 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg562 = (1'h0);
  reg [(5'h10):(1'h0)] reg561 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg560 = (1'h0);
  reg [(2'h3):(1'h0)] reg559 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg558 = (1'h0);
  reg [(2'h2):(1'h0)] reg557 = (1'h0);
  reg [(3'h6):(1'h0)] reg556 = (1'h0);
  reg [(3'h4):(1'h0)] reg555 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg554 = (1'h0);
  reg [(3'h4):(1'h0)] reg553 = (1'h0);
  reg [(2'h2):(1'h0)] reg552 = (1'h0);
  reg [(2'h2):(1'h0)] reg551 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg548 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg547 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg546 = (1'h0);
  reg signed [(4'he):(1'h0)] reg544 = (1'h0);
  reg [(4'hf):(1'h0)] reg543 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg540 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg539 = (1'h0);
  reg [(5'h10):(1'h0)] reg538 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg537 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg536 = (1'h0);
  reg [(3'h6):(1'h0)] reg535 = (1'h0);
  reg [(3'h6):(1'h0)] reg534 = (1'h0);
  reg [(4'h9):(1'h0)] reg533 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg531 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg530 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg529 = (1'h0);
  reg [(4'ha):(1'h0)] reg528 = (1'h0);
  reg [(3'h7):(1'h0)] reg527 = (1'h0);
  reg [(3'h7):(1'h0)] reg524 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg523 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg522 = (1'h0);
  reg [(4'hc):(1'h0)] reg521 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg520 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg519 = (1'h0);
  reg signed [(4'he):(1'h0)] reg518 = (1'h0);
  reg [(4'hb):(1'h0)] reg505 = (1'h0);
  reg [(3'h7):(1'h0)] reg515 = (1'h0);
  reg [(4'he):(1'h0)] reg513 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg512 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg511 = (1'h0);
  reg signed [(4'he):(1'h0)] reg510 = (1'h0);
  reg [(4'hf):(1'h0)] reg508 = (1'h0);
  reg [(4'hb):(1'h0)] reg507 = (1'h0);
  reg [(3'h6):(1'h0)] reg506 = (1'h0);
  reg [(4'hb):(1'h0)] reg504 = (1'h0);
  reg [(5'h10):(1'h0)] reg503 = (1'h0);
  reg [(3'h5):(1'h0)] reg502 = (1'h0);
  reg [(3'h6):(1'h0)] reg499 = (1'h0);
  reg [(4'ha):(1'h0)] reg498 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg497 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg496 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg495 = (1'h0);
  reg [(2'h3):(1'h0)] reg494 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg10 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg13 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg14 = (1'h0);
  reg [(4'ha):(1'h0)] reg16 = (1'h0);
  reg [(4'hf):(1'h0)] reg17 = (1'h0);
  reg signed [(4'he):(1'h0)] reg18 = (1'h0);
  reg [(3'h5):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg21 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg22 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg26 = (1'h0);
  reg [(2'h3):(1'h0)] reg27 = (1'h0);
  reg [(2'h2):(1'h0)] reg30 = (1'h0);
  reg [(4'h8):(1'h0)] reg32 = (1'h0);
  reg [(3'h6):(1'h0)] reg33 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg34 = (1'h0);
  reg [(3'h7):(1'h0)] reg36 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg37 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg38 = (1'h0);
  reg [(3'h5):(1'h0)] reg39 = (1'h0);
  reg [(4'h9):(1'h0)] reg40 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg42 = (1'h0);
  reg [(4'ha):(1'h0)] reg43 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg45 = (1'h0);
  reg [(4'hb):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg47 = (1'h0);
  reg [(4'hb):(1'h0)] reg48 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg50 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg51 = (1'h0);
  reg [(3'h5):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg54 = (1'h0);
  reg [(3'h5):(1'h0)] reg55 = (1'h0);
  reg [(4'hd):(1'h0)] reg56 = (1'h0);
  reg [(4'hd):(1'h0)] reg57 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg59 = (1'h0);
  reg [(4'h9):(1'h0)] reg60 = (1'h0);
  reg [(4'hc):(1'h0)] reg64 = (1'h0);
  reg [(4'h9):(1'h0)] reg65 = (1'h0);
  reg [(4'hc):(1'h0)] reg66 = (1'h0);
  reg [(3'h4):(1'h0)] reg68 = (1'h0);
  reg [(3'h7):(1'h0)] reg69 = (1'h0);
  reg [(2'h3):(1'h0)] reg70 = (1'h0);
  reg [(3'h6):(1'h0)] reg73 = (1'h0);
  reg [(3'h5):(1'h0)] reg75 = (1'h0);
  reg [(3'h5):(1'h0)] reg76 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg79 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg80 = (1'h0);
  reg [(4'he):(1'h0)] reg81 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg83 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg77 = (1'h0);
  reg [(4'hb):(1'h0)] reg82 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg84 = (1'h0);
  reg [(3'h5):(1'h0)] reg85 = (1'h0);
  reg [(4'hf):(1'h0)] reg88 = (1'h0);
  reg [(4'ha):(1'h0)] reg89 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg90 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg92 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg95 = (1'h0);
  reg [(4'he):(1'h0)] reg96 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg97 = (1'h0);
  reg [(4'hb):(1'h0)] reg98 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg100 = (1'h0);
  reg [(4'ha):(1'h0)] reg102 = (1'h0);
  reg [(4'hf):(1'h0)] reg104 = (1'h0);
  reg [(2'h2):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg106 = (1'h0);
  reg [(2'h3):(1'h0)] reg108 = (1'h0);
  reg [(3'h6):(1'h0)] reg109 = (1'h0);
  reg [(4'h8):(1'h0)] reg110 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg111 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg114 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg115 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg107 = (1'h0);
  reg [(3'h7):(1'h0)] reg112 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg101 = (1'h0);
  reg [(4'he):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg118 = (1'h0);
  reg [(3'h4):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg121 = (1'h0);
  reg [(3'h4):(1'h0)] reg124 = (1'h0);
  reg [(4'h9):(1'h0)] reg125 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg127 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg128 = (1'h0);
  reg [(4'ha):(1'h0)] reg99 = (1'h0);
  reg [(5'h10):(1'h0)] reg117 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg122 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg123 = (1'h0);
  reg [(4'he):(1'h0)] reg129 = (1'h0);
  reg [(3'h6):(1'h0)] reg130 = (1'h0);
  reg [(4'h9):(1'h0)] reg131 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg132 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg133 = (1'h0);
  reg [(4'h8):(1'h0)] reg134 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg135 = (1'h0);
  reg [(3'h7):(1'h0)] reg116 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg139 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg140 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg141 = (1'h0);
  reg [(2'h3):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg143 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg144 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg146 = (1'h0);
  reg [(2'h3):(1'h0)] reg147 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg148 = (1'h0);
  reg [(4'h9):(1'h0)] reg149 = (1'h0);
  reg [(4'h9):(1'h0)] reg150 = (1'h0);
  reg [(4'h9):(1'h0)] reg151 = (1'h0);
  reg [(4'h9):(1'h0)] reg152 = (1'h0);
  reg [(4'ha):(1'h0)] reg154 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg155 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg156 = (1'h0);
  reg [(2'h2):(1'h0)] reg157 = (1'h0);
  reg [(2'h3):(1'h0)] reg145 = (1'h0);
  reg [(4'h9):(1'h0)] reg159 = (1'h0);
  reg [(5'h10):(1'h0)] reg160 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg161 = (1'h0);
  reg [(3'h4):(1'h0)] reg164 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg166 = (1'h0);
  reg [(4'hb):(1'h0)] reg168 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg169 = (1'h0);
  reg [(4'h8):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg171 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg173 = (1'h0);
  reg [(2'h3):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg175 = (1'h0);
  reg [(2'h3):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg178 = (1'h0);
  reg [(5'h10):(1'h0)] reg179 = (1'h0);
  reg [(4'hc):(1'h0)] reg180 = (1'h0);
  reg [(3'h4):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg183 = (1'h0);
  reg [(4'he):(1'h0)] reg184 = (1'h0);
  reg signed [(4'he):(1'h0)] reg186 = (1'h0);
  reg [(4'hc):(1'h0)] reg187 = (1'h0);
  reg [(3'h4):(1'h0)] reg188 = (1'h0);
  reg signed [(4'he):(1'h0)] reg190 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg191 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg162 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg163 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg167 = (1'h0);
  reg signed [(4'he):(1'h0)] reg172 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg176 = (1'h0);
  reg [(4'h8):(1'h0)] reg185 = (1'h0);
  reg [(3'h4):(1'h0)] reg189 = (1'h0);
  reg signed [(4'he):(1'h0)] reg192 = (1'h0);
  reg [(4'h9):(1'h0)] reg193 = (1'h0);
  reg [(2'h2):(1'h0)] reg195 = (1'h0);
  reg [(5'h10):(1'h0)] reg194 = (1'h0);
  reg [(2'h2):(1'h0)] reg196 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg198 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg199 = (1'h0);
  reg [(4'he):(1'h0)] reg200 = (1'h0);
  reg [(5'h10):(1'h0)] reg201 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg197 = (1'h0);
  reg [(4'hb):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg204 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg205 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg206 = (1'h0);
  reg [(4'hd):(1'h0)] reg208 = (1'h0);
  reg [(4'hc):(1'h0)] reg209 = (1'h0);
  reg signed [(4'he):(1'h0)] reg210 = (1'h0);
  reg [(5'h10):(1'h0)] reg211 = (1'h0);
  reg signed [(4'he):(1'h0)] reg212 = (1'h0);
  reg [(4'hb):(1'h0)] reg213 = (1'h0);
  reg [(4'he):(1'h0)] reg207 = (1'h0);
  reg [(2'h3):(1'h0)] reg214 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg216 = (1'h0);
  reg [(2'h3):(1'h0)] reg217 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg219 = (1'h0);
  reg [(3'h7):(1'h0)] reg215 = (1'h0);
  reg [(4'h8):(1'h0)] reg220 = (1'h0);
  reg [(2'h3):(1'h0)] reg221 = (1'h0);
  reg [(4'ha):(1'h0)] reg222 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg223 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg225 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1176 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1171 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1167 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1166 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1151 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1146 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1162 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1145 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1144 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1139 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1133 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1125 = (1'h0);
  reg [(4'he):(1'h0)] forvar1121 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1117 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1113 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1110 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1103 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1100 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1098 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1090 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1083 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1078 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1077 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1074 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1068 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1067 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1066 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1063 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1058 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1056 = (1'h0);
  reg [(4'he):(1'h0)] forvar1044 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1043 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1060 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1054 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1050 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1046 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1045 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1042 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1038 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1033 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1032 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1028 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1024 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1009 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1014 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1011 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1006 = (1'h0);
  reg [(4'he):(1'h0)] forvar1005 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar996 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar993 = (1'h0);
  reg [(4'hc):(1'h0)] forvar982 = (1'h0);
  reg [(3'h6):(1'h0)] forvar978 = (1'h0);
  reg [(4'hc):(1'h0)] forvar968 = (1'h0);
  reg [(4'hb):(1'h0)] forvar966 = (1'h0);
  reg [(2'h3):(1'h0)] forvar973 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar975 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar965 = (1'h0);
  reg [(4'he):(1'h0)] forvar986 = (1'h0);
  reg [(3'h6):(1'h0)] forvar981 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar979 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar974 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar969 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar957 = (1'h0);
  reg [(3'h5):(1'h0)] forvar955 = (1'h0);
  reg [(3'h7):(1'h0)] forvar954 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar951 = (1'h0);
  reg [(5'h10):(1'h0)] forvar950 = (1'h0);
  reg [(3'h4):(1'h0)] forvar948 = (1'h0);
  reg [(2'h3):(1'h0)] forvar944 = (1'h0);
  reg [(4'hc):(1'h0)] forvar941 = (1'h0);
  reg [(4'hd):(1'h0)] forvar936 = (1'h0);
  reg [(4'hb):(1'h0)] forvar932 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar930 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar914 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar911 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar910 = (1'h0);
  reg [(3'h6):(1'h0)] forvar909 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar904 = (1'h0);
  reg [(3'h6):(1'h0)] forvar900 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar899 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar894 = (1'h0);
  reg [(4'h8):(1'h0)] forvar890 = (1'h0);
  reg [(4'ha):(1'h0)] forvar886 = (1'h0);
  reg [(3'h4):(1'h0)] forvar885 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar884 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar878 = (1'h0);
  reg [(4'h9):(1'h0)] forvar876 = (1'h0);
  reg [(4'hd):(1'h0)] forvar870 = (1'h0);
  reg [(2'h3):(1'h0)] forvar869 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar863 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar851 = (1'h0);
  reg [(3'h6):(1'h0)] forvar848 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar844 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar827 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar826 = (1'h0);
  reg [(3'h5):(1'h0)] forvar825 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar792 = (1'h0);
  reg [(3'h5):(1'h0)] forvar786 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar784 = (1'h0);
  reg [(4'hc):(1'h0)] forvar819 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar818 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar812 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar797 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar810 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar809 = (1'h0);
  reg [(3'h5):(1'h0)] forvar803 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar798 = (1'h0);
  reg [(4'h9):(1'h0)] forvar796 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar793 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar787 = (1'h0);
  reg [(3'h7):(1'h0)] forvar785 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar783 = (1'h0);
  reg [(4'h8):(1'h0)] forvar778 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar777 = (1'h0);
  reg [(3'h6):(1'h0)] forvar776 = (1'h0);
  reg [(5'h10):(1'h0)] forvar769 = (1'h0);
  reg [(4'hd):(1'h0)] forvar768 = (1'h0);
  reg [(4'hd):(1'h0)] forvar763 = (1'h0);
  reg [(3'h7):(1'h0)] forvar760 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar762 = (1'h0);
  reg [(4'he):(1'h0)] forvar756 = (1'h0);
  reg [(4'ha):(1'h0)] forvar749 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar744 = (1'h0);
  reg [(4'hb):(1'h0)] forvar743 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar738 = (1'h0);
  reg [(4'ha):(1'h0)] forvar729 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar727 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar719 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar717 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar711 = (1'h0);
  reg [(3'h4):(1'h0)] forvar710 = (1'h0);
  reg [(2'h2):(1'h0)] forvar753 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar748 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar746 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar745 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar737 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar736 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar730 = (1'h0);
  reg [(4'hb):(1'h0)] forvar732 = (1'h0);
  reg [(4'he):(1'h0)] forvar724 = (1'h0);
  reg [(5'h10):(1'h0)] forvar722 = (1'h0);
  reg [(4'he):(1'h0)] forvar720 = (1'h0);
  reg [(4'h9):(1'h0)] forvar714 = (1'h0);
  reg [(3'h5):(1'h0)] forvar709 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar661 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar658 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar656 = (1'h0);
  reg [(4'hc):(1'h0)] forvar703 = (1'h0);
  reg [(4'h9):(1'h0)] forvar700 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar696 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar692 = (1'h0);
  reg [(3'h4):(1'h0)] forvar684 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar701 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar698 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar697 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar685 = (1'h0);
  reg [(2'h2):(1'h0)] forvar678 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar676 = (1'h0);
  reg [(4'hd):(1'h0)] forvar669 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar668 = (1'h0);
  reg [(4'hf):(1'h0)] forvar660 = (1'h0);
  reg [(4'h8):(1'h0)] forvar655 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar652 = (1'h0);
  reg [(4'hb):(1'h0)] forvar647 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar639 = (1'h0);
  reg [(4'h8):(1'h0)] forvar635 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar651 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar640 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar636 = (1'h0);
  reg [(2'h2):(1'h0)] forvar632 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar625 = (1'h0);
  reg [(3'h7):(1'h0)] forvar620 = (1'h0);
  reg [(4'he):(1'h0)] forvar619 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar614 = (1'h0);
  reg [(2'h2):(1'h0)] forvar591 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar611 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar607 = (1'h0);
  reg [(4'hf):(1'h0)] forvar604 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar601 = (1'h0);
  reg [(4'h8):(1'h0)] forvar597 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar590 = (1'h0);
  reg [(4'h9):(1'h0)] forvar571 = (1'h0);
  reg [(4'hf):(1'h0)] forvar599 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar598 = (1'h0);
  reg [(2'h2):(1'h0)] forvar587 = (1'h0);
  reg [(4'hb):(1'h0)] forvar586 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar582 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar578 = (1'h0);
  reg [(3'h7):(1'h0)] forvar573 = (1'h0);
  reg [(4'h9):(1'h0)] forvar572 = (1'h0);
  reg [(4'he):(1'h0)] forvar512 = (1'h0);
  reg [(4'hd):(1'h0)] forvar519 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar511 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar524 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar520 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar510 = (1'h0);
  reg [(4'hf):(1'h0)] forvar508 = (1'h0);
  reg [(3'h6):(1'h0)] forvar499 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar496 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar502 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar536 = (1'h0);
  reg [(4'he):(1'h0)] forvar531 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar530 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar550 = (1'h0);
  reg [(2'h3):(1'h0)] forvar549 = (1'h0);
  reg [(4'ha):(1'h0)] forvar545 = (1'h0);
  reg [(4'hf):(1'h0)] forvar542 = (1'h0);
  reg [(3'h4):(1'h0)] forvar541 = (1'h0);
  reg [(4'hf):(1'h0)] forvar526 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar525 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar495 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar517 = (1'h0);
  reg [(2'h2):(1'h0)] forvar516 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar514 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar509 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar505 = (1'h0);
  reg [(4'hd):(1'h0)] forvar501 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar500 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar497 = (1'h0);
  reg [(4'h8):(1'h0)] forvar494 = (1'h0);
  reg [(4'hd):(1'h0)] forvar209 = (1'h0);
  reg [(4'hf):(1'h0)] forvar224 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar219 = (1'h0);
  reg [(3'h4):(1'h0)] forvar214 = (1'h0);
  reg [(3'h6):(1'h0)] forvar215 = (1'h0);
  reg [(5'h10):(1'h0)] forvar205 = (1'h0);
  reg [(3'h6):(1'h0)] forvar207 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar202 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar195 = (1'h0);
  reg [(3'h4):(1'h0)] forvar192 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar197 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar193 = (1'h0);
  reg [(4'h8):(1'h0)] forvar191 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar187 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar194 = (1'h0);
  reg [(4'h9):(1'h0)] forvar186 = (1'h0);
  reg [(4'h8):(1'h0)] forvar166 = (1'h0);
  reg [(3'h5):(1'h0)] forvar174 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar169 = (1'h0);
  reg [(3'h6):(1'h0)] forvar164 = (1'h0);
  reg [(3'h5):(1'h0)] forvar189 = (1'h0);
  reg [(4'h9):(1'h0)] forvar185 = (1'h0);
  reg [(2'h3):(1'h0)] forvar181 = (1'h0);
  reg [(4'hc):(1'h0)] forvar176 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar172 = (1'h0);
  reg [(4'hb):(1'h0)] forvar167 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar163 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar162 = (1'h0);
  reg [(3'h6):(1'h0)] forvar158 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar153 = (1'h0);
  reg [(2'h2):(1'h0)] forvar145 = (1'h0);
  reg [(3'h7):(1'h0)] forvar138 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar137 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar136 = (1'h0);
  reg [(4'hf):(1'h0)] forvar125 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar121 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar114 = (1'h0);
  reg [(3'h6):(1'h0)] forvar131 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar127 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar115 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar108 = (1'h0);
  reg [(4'hf):(1'h0)] forvar109 = (1'h0);
  reg [(4'hc):(1'h0)] forvar123 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar122 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar117 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar116 = (1'h0);
  reg [(4'hf):(1'h0)] forvar104 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar105 = (1'h0);
  reg [(2'h2):(1'h0)] forvar112 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar107 = (1'h0);
  reg [(4'ha):(1'h0)] forvar103 = (1'h0);
  reg [(3'h6):(1'h0)] forvar101 = (1'h0);
  reg [(3'h5):(1'h0)] forvar99 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar94 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar91 = (1'h0);
  reg [(4'ha):(1'h0)] forvar87 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar86 = (1'h0);
  reg [(3'h6):(1'h0)] forvar78 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar82 = (1'h0);
  reg [(3'h5):(1'h0)] forvar77 = (1'h0);
  reg [(4'he):(1'h0)] forvar74 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar72 = (1'h0);
  reg [(4'he):(1'h0)] forvar71 = (1'h0);
  reg [(3'h7):(1'h0)] forvar67 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar63 = (1'h0);
  reg [(4'hd):(1'h0)] forvar62 = (1'h0);
  reg [(4'hd):(1'h0)] forvar61 = (1'h0);
  reg [(4'hc):(1'h0)] forvar58 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar53 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar49 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar46 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar40 = (1'h0);
  reg [(3'h7):(1'h0)] forvar41 = (1'h0);
  reg [(3'h4):(1'h0)] forvar35 = (1'h0);
  reg [(3'h6):(1'h0)] forvar31 = (1'h0);
  reg [(4'hc):(1'h0)] forvar29 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar28 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar25 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar24 = (1'h0);
  reg [(5'h10):(1'h0)] forvar20 = (1'h0);
  reg [(4'hb):(1'h0)] forvar15 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar12 = (1'h0);
  reg [(3'h7):(1'h0)] forvar11 = (1'h0);
  assign y = {wire3402,
                 wire1179,
                 wire1040,
                 wire964,
                 wire708,
                 wire707,
                 wire492,
                 reg1176,
                 reg1167,
                 reg1178,
                 reg1177,
                 reg1175,
                 reg1174,
                 reg1173,
                 reg1172,
                 reg1170,
                 reg1169,
                 reg1168,
                 reg1145,
                 reg1165,
                 reg1164,
                 reg1163,
                 reg1161,
                 reg1160,
                 reg1159,
                 reg1158,
                 reg1157,
                 reg1156,
                 reg1155,
                 reg1154,
                 reg1153,
                 reg1152,
                 reg1151,
                 reg1150,
                 reg1149,
                 reg1148,
                 reg1147,
                 reg1146,
                 reg1133,
                 reg1143,
                 reg1142,
                 reg1141,
                 reg1140,
                 reg1138,
                 reg1137,
                 reg1136,
                 reg1135,
                 reg1134,
                 reg1132,
                 reg1125,
                 reg1131,
                 reg1130,
                 reg1129,
                 reg1128,
                 reg1127,
                 reg1126,
                 reg1124,
                 reg1123,
                 reg1122,
                 reg1120,
                 reg1119,
                 reg1118,
                 reg1116,
                 reg1113,
                 reg1115,
                 reg1114,
                 reg1112,
                 reg1111,
                 reg1110,
                 reg1109,
                 reg1108,
                 reg1107,
                 reg1106,
                 reg1105,
                 reg1104,
                 reg1103,
                 reg1102,
                 reg1101,
                 reg1090,
                 reg1099,
                 reg1097,
                 reg1096,
                 reg1095,
                 reg1094,
                 reg1093,
                 reg1092,
                 reg1091,
                 reg1089,
                 reg1088,
                 reg1087,
                 reg1086,
                 reg1085,
                 reg1084,
                 reg1082,
                 reg1081,
                 reg1080,
                 reg1079,
                 reg1076,
                 reg1075,
                 reg1073,
                 reg1072,
                 reg1071,
                 reg1070,
                 reg1069,
                 reg1065,
                 reg1064,
                 reg1045,
                 reg1042,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 reg1057,
                 reg1056,
                 reg1055,
                 reg1053,
                 reg1052,
                 reg1051,
                 reg1046,
                 reg1050,
                 reg1049,
                 reg1048,
                 reg1047,
                 reg1044,
                 reg1043,
                 reg1041,
                 reg1039,
                 reg1037,
                 reg1036,
                 reg1035,
                 reg1034,
                 reg1031,
                 reg1030,
                 reg1029,
                 reg1027,
                 reg1026,
                 reg1025,
                 reg1024,
                 reg1023,
                 reg1022,
                 reg1021,
                 reg1020,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1011,
                 reg1016,
                 reg1015,
                 reg1013,
                 reg1012,
                 reg1010,
                 reg1009,
                 reg1008,
                 reg1007,
                 reg993,
                 reg1004,
                 reg1003,
                 reg1002,
                 reg1001,
                 reg1000,
                 reg999,
                 reg998,
                 reg997,
                 reg995,
                 reg994,
                 reg992,
                 reg991,
                 reg979,
                 reg986,
                 reg981,
                 reg974,
                 reg990,
                 reg989,
                 reg988,
                 reg987,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 reg980,
                 reg969,
                 reg978,
                 reg977,
                 reg976,
                 reg975,
                 reg973,
                 reg972,
                 reg971,
                 reg970,
                 reg968,
                 reg967,
                 reg966,
                 reg965,
                 reg963,
                 reg962,
                 reg961,
                 reg960,
                 reg959,
                 reg958,
                 reg956,
                 reg953,
                 reg952,
                 reg949,
                 reg947,
                 reg946,
                 reg945,
                 reg943,
                 reg942,
                 reg932,
                 reg930,
                 reg940,
                 reg939,
                 reg938,
                 reg937,
                 reg935,
                 reg934,
                 reg933,
                 reg931,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 reg925,
                 reg924,
                 reg923,
                 reg922,
                 reg921,
                 reg920,
                 reg919,
                 reg918,
                 reg917,
                 reg916,
                 reg915,
                 reg913,
                 reg912,
                 reg908,
                 reg907,
                 reg906,
                 reg905,
                 reg903,
                 reg902,
                 reg901,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg893,
                 reg892,
                 reg890,
                 reg891,
                 reg889,
                 reg888,
                 reg887,
                 reg883,
                 reg882,
                 reg881,
                 reg880,
                 reg879,
                 reg877,
                 reg875,
                 reg874,
                 reg873,
                 reg872,
                 reg871,
                 reg868,
                 reg867,
                 reg866,
                 reg865,
                 reg864,
                 reg862,
                 reg861,
                 reg860,
                 reg859,
                 reg851,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 reg852,
                 reg850,
                 reg849,
                 reg847,
                 reg846,
                 reg845,
                 reg843,
                 reg842,
                 reg841,
                 reg840,
                 reg839,
                 reg838,
                 reg837,
                 reg836,
                 reg835,
                 reg834,
                 reg833,
                 reg832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg783,
                 reg824,
                 reg823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 reg818,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 reg793,
                 reg798,
                 reg796,
                 reg811,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 reg797,
                 reg795,
                 reg794,
                 reg792,
                 reg791,
                 reg790,
                 reg789,
                 reg788,
                 reg785,
                 reg787,
                 reg786,
                 reg784,
                 reg782,
                 reg781,
                 reg780,
                 reg779,
                 reg775,
                 reg774,
                 reg773,
                 reg772,
                 reg768,
                 reg771,
                 reg770,
                 reg769,
                 reg762,
                 reg756,
                 reg767,
                 reg766,
                 reg765,
                 reg764,
                 reg763,
                 reg761,
                 reg760,
                 reg759,
                 reg758,
                 reg757,
                 reg753,
                 reg748,
                 reg746,
                 reg745,
                 reg737,
                 reg732,
                 reg714,
                 reg755,
                 reg754,
                 reg752,
                 reg751,
                 reg750,
                 reg749,
                 reg747,
                 reg744,
                 reg743,
                 reg742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 reg735,
                 reg734,
                 reg733,
                 reg731,
                 reg730,
                 reg729,
                 reg728,
                 reg727,
                 reg720,
                 reg722,
                 reg726,
                 reg725,
                 reg724,
                 reg723,
                 reg721,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg713,
                 reg712,
                 reg711,
                 reg710,
                 reg709,
                 reg706,
                 reg705,
                 reg704,
                 reg701,
                 reg698,
                 reg697,
                 reg685,
                 reg702,
                 reg700,
                 reg699,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg689,
                 reg688,
                 reg687,
                 reg686,
                 reg684,
                 reg683,
                 reg682,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg675,
                 reg674,
                 reg673,
                 reg668,
                 reg672,
                 reg671,
                 reg670,
                 reg669,
                 reg667,
                 reg666,
                 reg665,
                 reg660,
                 reg655,
                 reg664,
                 reg663,
                 reg662,
                 reg661,
                 reg659,
                 reg658,
                 reg657,
                 reg656,
                 reg651,
                 reg636,
                 reg654,
                 reg653,
                 reg652,
                 reg650,
                 reg649,
                 reg648,
                 reg647,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 reg642,
                 reg641,
                 reg639,
                 reg638,
                 reg637,
                 reg635,
                 reg614,
                 reg634,
                 reg633,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 reg618,
                 reg617,
                 reg616,
                 reg615,
                 reg587,
                 reg598,
                 reg613,
                 reg612,
                 reg610,
                 reg609,
                 reg608,
                 reg606,
                 reg599,
                 reg586,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg585,
                 reg584,
                 reg583,
                 reg578,
                 reg573,
                 reg582,
                 reg581,
                 reg580,
                 reg579,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 reg571,
                 reg525,
                 reg516,
                 reg514,
                 reg526,
                 reg517,
                 reg509,
                 reg501,
                 reg500,
                 reg545,
                 reg542,
                 reg541,
                 reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 reg551,
                 reg548,
                 reg547,
                 reg546,
                 reg544,
                 reg543,
                 reg540,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg505,
                 reg515,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg508,
                 reg507,
                 reg506,
                 reg504,
                 reg503,
                 reg502,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg10,
                 reg13,
                 reg14,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg21,
                 reg22,
                 reg23,
                 reg26,
                 reg27,
                 reg30,
                 reg32,
                 reg33,
                 reg34,
                 reg36,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 reg42,
                 reg43,
                 reg44,
                 reg45,
                 reg41,
                 reg47,
                 reg48,
                 reg50,
                 reg51,
                 reg52,
                 reg54,
                 reg55,
                 reg56,
                 reg57,
                 reg59,
                 reg60,
                 reg64,
                 reg65,
                 reg66,
                 reg68,
                 reg69,
                 reg70,
                 reg73,
                 reg75,
                 reg76,
                 reg78,
                 reg79,
                 reg80,
                 reg81,
                 reg83,
                 reg74,
                 reg77,
                 reg82,
                 reg84,
                 reg85,
                 reg88,
                 reg89,
                 reg90,
                 reg92,
                 reg93,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 reg100,
                 reg102,
                 reg104,
                 reg105,
                 reg106,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg113,
                 reg114,
                 reg115,
                 reg107,
                 reg112,
                 reg101,
                 reg103,
                 reg118,
                 reg119,
                 reg120,
                 reg121,
                 reg124,
                 reg125,
                 reg126,
                 reg127,
                 reg128,
                 reg99,
                 reg117,
                 reg122,
                 reg123,
                 reg129,
                 reg130,
                 reg131,
                 reg132,
                 reg133,
                 reg134,
                 reg135,
                 reg116,
                 reg139,
                 reg140,
                 reg141,
                 reg142,
                 reg143,
                 reg144,
                 reg146,
                 reg147,
                 reg148,
                 reg149,
                 reg150,
                 reg151,
                 reg152,
                 reg154,
                 reg155,
                 reg156,
                 reg157,
                 reg145,
                 reg159,
                 reg160,
                 reg161,
                 reg164,
                 reg165,
                 reg166,
                 reg168,
                 reg169,
                 reg170,
                 reg171,
                 reg173,
                 reg174,
                 reg175,
                 reg177,
                 reg178,
                 reg179,
                 reg180,
                 reg182,
                 reg183,
                 reg184,
                 reg186,
                 reg187,
                 reg188,
                 reg190,
                 reg191,
                 reg162,
                 reg163,
                 reg167,
                 reg172,
                 reg176,
                 reg185,
                 reg189,
                 reg192,
                 reg193,
                 reg195,
                 reg194,
                 reg196,
                 reg198,
                 reg199,
                 reg200,
                 reg201,
                 reg197,
                 reg203,
                 reg204,
                 reg205,
                 reg206,
                 reg208,
                 reg209,
                 reg210,
                 reg211,
                 reg212,
                 reg213,
                 reg207,
                 reg214,
                 reg216,
                 reg217,
                 reg218,
                 reg219,
                 reg215,
                 reg220,
                 reg221,
                 reg222,
                 reg223,
                 reg225,
                 forvar1176,
                 forvar1171,
                 forvar1167,
                 forvar1166,
                 forvar1151,
                 forvar1146,
                 forvar1162,
                 forvar1145,
                 forvar1144,
                 forvar1139,
                 forvar1133,
                 forvar1125,
                 forvar1121,
                 forvar1117,
                 forvar1113,
                 forvar1110,
                 forvar1103,
                 forvar1100,
                 forvar1098,
                 forvar1090,
                 forvar1083,
                 forvar1078,
                 forvar1077,
                 forvar1074,
                 forvar1068,
                 forvar1067,
                 forvar1066,
                 forvar1063,
                 forvar1058,
                 forvar1056,
                 forvar1044,
                 forvar1043,
                 forvar1060,
                 forvar1054,
                 forvar1050,
                 forvar1046,
                 forvar1045,
                 forvar1042,
                 forvar1038,
                 forvar1033,
                 forvar1032,
                 forvar1028,
                 forvar1024,
                 forvar1009,
                 forvar1014,
                 forvar1011,
                 forvar1006,
                 forvar1005,
                 forvar996,
                 forvar993,
                 forvar982,
                 forvar978,
                 forvar968,
                 forvar966,
                 forvar973,
                 forvar975,
                 forvar965,
                 forvar986,
                 forvar981,
                 forvar979,
                 forvar974,
                 forvar969,
                 forvar957,
                 forvar955,
                 forvar954,
                 forvar951,
                 forvar950,
                 forvar948,
                 forvar944,
                 forvar941,
                 forvar936,
                 forvar932,
                 forvar930,
                 forvar914,
                 forvar911,
                 forvar910,
                 forvar909,
                 forvar904,
                 forvar900,
                 forvar899,
                 forvar894,
                 forvar890,
                 forvar886,
                 forvar885,
                 forvar884,
                 forvar878,
                 forvar876,
                 forvar870,
                 forvar869,
                 forvar863,
                 forvar851,
                 forvar848,
                 forvar844,
                 forvar827,
                 forvar826,
                 forvar825,
                 forvar792,
                 forvar786,
                 forvar784,
                 forvar819,
                 forvar818,
                 forvar812,
                 forvar797,
                 forvar810,
                 forvar809,
                 forvar803,
                 forvar798,
                 forvar796,
                 forvar793,
                 forvar787,
                 forvar785,
                 forvar783,
                 forvar778,
                 forvar777,
                 forvar776,
                 forvar769,
                 forvar768,
                 forvar763,
                 forvar760,
                 forvar762,
                 forvar756,
                 forvar749,
                 forvar744,
                 forvar743,
                 forvar738,
                 forvar729,
                 forvar727,
                 forvar719,
                 forvar717,
                 forvar711,
                 forvar710,
                 forvar753,
                 forvar748,
                 forvar746,
                 forvar745,
                 forvar737,
                 forvar736,
                 forvar730,
                 forvar732,
                 forvar724,
                 forvar722,
                 forvar720,
                 forvar714,
                 forvar709,
                 forvar661,
                 forvar658,
                 forvar656,
                 forvar703,
                 forvar700,
                 forvar696,
                 forvar692,
                 forvar684,
                 forvar701,
                 forvar698,
                 forvar697,
                 forvar685,
                 forvar678,
                 forvar676,
                 forvar669,
                 forvar668,
                 forvar660,
                 forvar655,
                 forvar652,
                 forvar647,
                 forvar639,
                 forvar635,
                 forvar651,
                 forvar640,
                 forvar636,
                 forvar632,
                 forvar625,
                 forvar620,
                 forvar619,
                 forvar614,
                 forvar591,
                 forvar611,
                 forvar607,
                 forvar604,
                 forvar601,
                 forvar597,
                 forvar590,
                 forvar571,
                 forvar599,
                 forvar598,
                 forvar587,
                 forvar586,
                 forvar582,
                 forvar578,
                 forvar573,
                 forvar572,
                 forvar512,
                 forvar519,
                 forvar511,
                 forvar524,
                 forvar520,
                 forvar510,
                 forvar508,
                 forvar499,
                 forvar496,
                 forvar502,
                 forvar536,
                 forvar531,
                 forvar530,
                 forvar550,
                 forvar549,
                 forvar545,
                 forvar542,
                 forvar541,
                 forvar526,
                 forvar525,
                 forvar495,
                 forvar517,
                 forvar516,
                 forvar514,
                 forvar509,
                 forvar505,
                 forvar501,
                 forvar500,
                 forvar497,
                 forvar494,
                 forvar209,
                 forvar224,
                 forvar219,
                 forvar214,
                 forvar215,
                 forvar205,
                 forvar207,
                 forvar202,
                 forvar195,
                 forvar192,
                 forvar197,
                 forvar193,
                 forvar191,
                 forvar187,
                 forvar194,
                 forvar186,
                 forvar166,
                 forvar174,
                 forvar169,
                 forvar164,
                 forvar189,
                 forvar185,
                 forvar181,
                 forvar176,
                 forvar172,
                 forvar167,
                 forvar163,
                 forvar162,
                 forvar158,
                 forvar153,
                 forvar145,
                 forvar138,
                 forvar137,
                 forvar136,
                 forvar125,
                 forvar121,
                 forvar114,
                 forvar131,
                 forvar127,
                 forvar115,
                 forvar108,
                 forvar109,
                 forvar123,
                 forvar122,
                 forvar117,
                 forvar116,
                 forvar104,
                 forvar105,
                 forvar112,
                 forvar107,
                 forvar103,
                 forvar101,
                 forvar99,
                 forvar94,
                 forvar91,
                 forvar87,
                 forvar86,
                 forvar78,
                 forvar82,
                 forvar77,
                 forvar74,
                 forvar72,
                 forvar71,
                 forvar67,
                 forvar63,
                 forvar62,
                 forvar61,
                 forvar58,
                 forvar53,
                 forvar49,
                 forvar46,
                 forvar40,
                 forvar41,
                 forvar35,
                 forvar31,
                 forvar29,
                 forvar28,
                 forvar25,
                 forvar24,
                 forvar20,
                 forvar15,
                 forvar12,
                 forvar11,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned({wire8[(2'h3):(1'h0)]}))
        begin
          reg10 <= wire7[(4'ha):(1'h1)];
          for (forvar11 = (1'h0); (forvar11 < (2'h2)); forvar11 = (forvar11 + (1'h1)))
            begin
              for (forvar12 = (1'h0); (forvar12 < (1'h0)); forvar12 = (forvar12 + (1'h1)))
                begin
                  reg13 <= {wire7};
                  reg14 <= wire6[(2'h2):(2'h2)];
                end
              for (forvar15 = (1'h0); (forvar15 < (2'h3)); forvar15 = (forvar15 + (1'h1)))
                begin
                  if ((!forvar12[(4'h8):(1'h0)]))
                    begin
                      reg16 <= $unsigned($unsigned({(wire8 < reg10)}));
                      reg17 <= reg13[(1'h1):(1'h1)];
                      reg18 <= $unsigned(forvar12[(3'h6):(1'h1)]);
                      reg19 <= ((wire6 * (~&wire8[(1'h0):(1'h0)])) + forvar12);
                    end
                  else
                    begin
                      reg16 <= $unsigned(reg19);
                      reg17 <= (~(^reg19[(3'h5):(3'h4)]));
                    end
                  for (forvar20 = (1'h0); (forvar20 < (2'h3)); forvar20 = (forvar20 + (1'h1)))
                    begin
                      reg21 <= $unsigned($unsigned($unsigned((forvar15 * reg17))));
                    end
                  if (reg14)
                    begin
                      reg22 <= $unsigned({($unsigned(reg13) - reg17[(3'h5):(2'h2)])});
                    end
                  else
                    begin
                      reg22 <= $unsigned($unsigned($signed($signed(forvar20))));
                      reg23 <= $unsigned((((reg17 == reg22) & (reg13 ^~ reg13)) <= $unsigned((~&forvar12))));
                    end
                end
            end
          for (forvar24 = (1'h0); (forvar24 < (1'h1)); forvar24 = (forvar24 + (1'h1)))
            begin
              for (forvar25 = (1'h0); (forvar25 < (2'h3)); forvar25 = (forvar25 + (1'h1)))
                begin
                  if ((forvar15[(1'h0):(1'h0)] - wire7[(4'h8):(1'h0)]))
                    begin
                      reg26 <= (reg21[(3'h6):(3'h6)] ?
                          (+((wire6 > forvar25) == (forvar24 ?
                              wire8 : reg23))) : {((&(8'hb8)) > forvar25[(4'hc):(4'h8)])});
                      reg27 <= forvar24[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg26 <= ((|((reg27 ? reg18 : (8'hb9)) ?
                          (reg26 ?
                              wire6 : reg16) : $unsigned(wire8))) == (((8'ha2) >= (reg23 ?
                              (8'ha4) : (8'hb7))) ?
                          $signed(((8'h9c) ?
                              reg22 : forvar20)) : ($signed(reg27) ?
                              (-(8'ha0)) : {reg16})));
                    end
                end
              for (forvar28 = (1'h0); (forvar28 < (2'h2)); forvar28 = (forvar28 + (1'h1)))
                begin
                  for (forvar29 = (1'h0); (forvar29 < (2'h2)); forvar29 = (forvar29 + (1'h1)))
                    begin
                      reg30 <= {forvar12};
                    end
                  for (forvar31 = (1'h0); (forvar31 < (2'h3)); forvar31 = (forvar31 + (1'h1)))
                    begin
                      reg32 <= {$unsigned(((forvar11 ^~ reg16) >>> (forvar24 ?
                              (8'haf) : (8'had))))};
                      reg33 <= reg13;
                      reg34 <= reg16[(1'h1):(1'h1)];
                    end
                end
              if (forvar31[(2'h2):(2'h2)])
                begin
                  for (forvar35 = (1'h0); (forvar35 < (1'h0)); forvar35 = (forvar35 + (1'h1)))
                    begin
                      reg36 <= (reg19 > $unsigned($unsigned((-wire6))));
                      reg37 <= {$signed($unsigned((reg27 ^ reg22)))};
                      reg38 <= {{reg34[(2'h3):(2'h3)]}};
                    end
                  if (forvar35[(2'h2):(1'h1)])
                    begin
                      reg39 <= (($unsigned($unsigned(forvar28)) ?
                              (!(reg13 ? reg16 : forvar35)) : (+(~forvar25))) ?
                          {(reg32[(3'h5):(1'h1)] ?
                                  ((8'ha3) > forvar25) : (^reg17))} : $unsigned({(forvar35 <<< forvar24)}));
                      reg40 <= (($unsigned($signed(forvar31)) || (8'hb9)) != ((reg34 ?
                          {forvar31} : reg19) ^ $signed((reg38 ?
                          reg30 : wire7))));
                    end
                  else
                    begin
                      reg39 <= {forvar15};
                      reg40 <= {($signed((reg10 == reg26)) ?
                              reg22[(1'h1):(1'h1)] : reg21[(2'h3):(1'h1)])};
                    end
                  for (forvar41 = (1'h0); (forvar41 < (1'h0)); forvar41 = (forvar41 + (1'h1)))
                    begin
                      reg42 <= (-(+(reg40 ^ $unsigned((8'hab)))));
                      reg43 <= forvar41[(2'h2):(1'h1)];
                      reg44 <= $unsigned({(reg33[(2'h2):(2'h2)] == (reg17 && reg33))});
                      reg45 <= ($unsigned($signed($signed(wire9))) ?
                          ($signed((^reg23)) ?
                              (~&(forvar28 < reg43)) : (~|(|reg26))) : ({reg27} ^~ $signed((~reg34))));
                    end
                end
              else
                begin
                  for (forvar35 = (1'h0); (forvar35 < (1'h0)); forvar35 = (forvar35 + (1'h1)))
                    begin
                      reg36 <= (reg32[(3'h7):(3'h6)] + (wire6[(4'ha):(3'h7)] ?
                          $unsigned((^reg26)) : reg19));
                      reg37 <= $unsigned($unsigned(forvar24));
                      reg38 <= {$unsigned((reg14 ?
                              $signed(reg37) : $signed(reg21)))};
                      reg39 <= $signed($signed($unsigned($unsigned((8'ha4)))));
                    end
                  for (forvar40 = (1'h0); (forvar40 < (1'h0)); forvar40 = (forvar40 + (1'h1)))
                    begin
                      reg41 <= reg17[(2'h2):(2'h2)];
                    end
                end
              for (forvar46 = (1'h0); (forvar46 < (2'h2)); forvar46 = (forvar46 + (1'h1)))
                begin
                  if (wire8[(2'h3):(1'h1)])
                    begin
                      reg47 <= ($unsigned({((8'hb3) ?
                              forvar29 : forvar31)}) <<< {forvar25});
                      reg48 <= $unsigned(reg27[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg47 <= $unsigned(wire8[(3'h4):(2'h2)]);
                      reg48 <= (~reg47[(3'h5):(1'h1)]);
                    end
                  for (forvar49 = (1'h0); (forvar49 < (2'h3)); forvar49 = (forvar49 + (1'h1)))
                    begin
                      reg50 <= $unsigned(reg14[(2'h2):(2'h2)]);
                      reg51 <= $unsigned(wire6[(3'h6):(3'h6)]);
                      reg52 <= reg42;
                    end
                  for (forvar53 = (1'h0); (forvar53 < (1'h0)); forvar53 = (forvar53 + (1'h1)))
                    begin
                      reg54 <= forvar49;
                      reg55 <= (reg40[(3'h7):(2'h2)] <<< $signed(reg23));
                      reg56 <= reg54;
                      reg57 <= $unsigned(forvar31[(3'h4):(2'h2)]);
                    end
                  for (forvar58 = (1'h0); (forvar58 < (2'h2)); forvar58 = (forvar58 + (1'h1)))
                    begin
                      reg59 <= forvar58[(4'ha):(4'h8)];
                      reg60 <= ($unsigned(forvar11) ?
                          ($unsigned(reg19) || forvar53) : reg56[(2'h3):(1'h0)]);
                    end
                end
            end
          for (forvar61 = (1'h0); (forvar61 < (1'h1)); forvar61 = (forvar61 + (1'h1)))
            begin
              for (forvar62 = (1'h0); (forvar62 < (1'h0)); forvar62 = (forvar62 + (1'h1)))
                begin
                  for (forvar63 = (1'h0); (forvar63 < (2'h3)); forvar63 = (forvar63 + (1'h1)))
                    begin
                      reg64 <= (8'ha0);
                      reg65 <= (((((8'hb7) ?
                              forvar46 : wire6) * $unsigned(reg52)) ^~ (((8'ha9) ?
                                  wire8 : (8'ha8)) ?
                              (reg50 - reg50) : (forvar12 ? reg48 : reg51))) ?
                          ((~(reg34 ? (8'hb2) : (8'hba))) ?
                              ($signed(reg57) ?
                                  reg60 : $signed(reg36)) : forvar25) : reg47);
                      reg66 <= (&$unsigned({{reg43}}));
                    end
                  for (forvar67 = (1'h0); (forvar67 < (2'h3)); forvar67 = (forvar67 + (1'h1)))
                    begin
                      reg68 <= wire7;
                      reg69 <= reg59[(3'h7):(2'h3)];
                      reg70 <= $unsigned(reg44);
                    end
                end
            end
        end
      else
        begin
          reg10 <= reg36;
        end
      for (forvar71 = (1'h0); (forvar71 < (2'h3)); forvar71 = (forvar71 + (1'h1)))
        begin
          for (forvar72 = (1'h0); (forvar72 < (1'h1)); forvar72 = (forvar72 + (1'h1)))
            begin
              reg73 <= forvar49[(3'h4):(3'h4)];
              if ($unsigned(($unsigned(reg69) ?
                  (reg23[(4'h8):(3'h6)] ?
                      reg69[(3'h6):(3'h6)] : wire8) : reg34)))
                begin
                  for (forvar74 = (1'h0); (forvar74 < (2'h3)); forvar74 = (forvar74 + (1'h1)))
                    begin
                      reg75 <= ((!(((8'ha8) == reg52) ~^ (reg65 ^~ reg52))) ?
                          (wire8 << $signed((reg64 ?
                              (8'haa) : (8'ha6)))) : reg48[(3'h6):(3'h6)]);
                    end
                  reg76 <= ((!(^{reg10})) * ((reg18 && (forvar28 ?
                      reg23 : reg34)) << {forvar12}));
                  for (forvar77 = (1'h0); (forvar77 < (2'h2)); forvar77 = (forvar77 + (1'h1)))
                    begin
                      reg78 <= (((reg55[(2'h2):(2'h2)] > (&forvar35)) & $signed($unsigned(reg44))) ^~ $unsigned((-reg50)));
                      reg79 <= $unsigned({reg75[(2'h3):(1'h1)]});
                      reg80 <= ((|reg59[(3'h6):(1'h1)]) ~^ ($unsigned((reg78 <= (8'hab))) ?
                          reg39 : {$unsigned(forvar72)}));
                      reg81 <= $unsigned(forvar72[(1'h1):(1'h1)]);
                    end
                  for (forvar82 = (1'h0); (forvar82 < (1'h1)); forvar82 = (forvar82 + (1'h1)))
                    begin
                      reg83 <= $signed(reg43);
                    end
                end
              else
                begin
                  if ((reg39[(2'h3):(1'h0)] ?
                      {(reg33[(3'h6):(1'h0)] >>> (reg68 != reg36))} : wire6[(2'h3):(1'h1)]))
                    begin
                      reg74 <= $unsigned($unsigned($signed(forvar77[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg74 <= (($signed((forvar58 ? reg41 : forvar24)) ?
                          reg45[(4'hb):(4'h9)] : $signed($signed(reg73))) << forvar11);
                      reg75 <= (forvar61 ?
                          ($unsigned(reg55[(2'h2):(2'h2)]) ~^ $signed(reg75[(1'h0):(1'h0)])) : $signed($unsigned(reg65)));
                      reg76 <= $unsigned(reg43);
                      reg77 <= $signed(reg51[(2'h2):(2'h2)]);
                    end
                  for (forvar78 = (1'h0); (forvar78 < (2'h3)); forvar78 = (forvar78 + (1'h1)))
                    begin
                      reg79 <= $signed(((~|(~&(8'ha4))) ?
                          $signed($unsigned(reg30)) : (|$unsigned(forvar74))));
                      reg80 <= ($signed({reg60}) ?
                          $unsigned($unsigned({reg38})) : ($signed($unsigned(reg18)) ?
                              (~|$unsigned(forvar63)) : forvar67[(3'h6):(1'h1)]));
                    end
                  reg81 <= ((~^(^(8'hb0))) ?
                      (|((&reg22) * $signed(reg38))) : (reg26 ?
                          $unsigned((reg79 & (8'hab))) : {reg75}));
                  if (reg47)
                    begin
                      reg82 <= $unsigned(reg52);
                    end
                  else
                    begin
                      reg82 <= $signed($unsigned($signed($signed(forvar20))));
                      reg83 <= (~&forvar49[(1'h0):(1'h0)]);
                      reg84 <= (($unsigned(reg81) ?
                              (wire9 | wire7[(1'h1):(1'h1)]) : reg73[(2'h2):(1'h0)]) ?
                          (^~($signed(forvar15) ?
                              reg36[(3'h6):(2'h3)] : forvar58)) : reg21[(1'h0):(1'h0)]);
                      reg85 <= reg33[(2'h3):(1'h1)];
                    end
                end
              for (forvar86 = (1'h0); (forvar86 < (2'h2)); forvar86 = (forvar86 + (1'h1)))
                begin
                  for (forvar87 = (1'h0); (forvar87 < (1'h1)); forvar87 = (forvar87 + (1'h1)))
                    begin
                      reg88 <= {{$signed($signed(reg65))}};
                      reg89 <= $signed(reg70[(2'h3):(1'h1)]);
                      reg90 <= (~&(((reg68 == forvar11) <<< $unsigned(reg55)) || forvar41[(2'h2):(2'h2)]));
                    end
                  for (forvar91 = (1'h0); (forvar91 < (2'h3)); forvar91 = (forvar91 + (1'h1)))
                    begin
                      reg92 <= ($unsigned((8'ha8)) >>> $unsigned((^~((8'ha5) ?
                          reg66 : reg75))));
                    end
                  reg93 <= forvar71;
                  for (forvar94 = (1'h0); (forvar94 < (1'h0)); forvar94 = (forvar94 + (1'h1)))
                    begin
                      reg95 <= (forvar72 && {((!(8'hb0)) ?
                              (|forvar63) : {forvar58})});
                      reg96 <= (reg92[(4'h8):(2'h2)] ?
                          $signed(($signed(forvar77) ?
                              (reg47 << (8'haa)) : ((8'haf) != (8'ha5)))) : ((~reg41[(3'h5):(3'h5)]) + $unsigned((8'hb9))));
                      reg97 <= $signed(reg36[(3'h7):(2'h3)]);
                      reg98 <= $unsigned((8'ha3));
                    end
                end
            end
        end
      if (((($unsigned(reg27) & (reg70 & reg44)) ?
          forvar35[(1'h0):(1'h0)] : (&$signed(forvar78))) >> $signed(reg18)))
        begin
          if ((8'h9c))
            begin
              for (forvar99 = (1'h0); (forvar99 < (2'h2)); forvar99 = (forvar99 + (1'h1)))
                begin
                  reg100 <= (-reg66[(4'hc):(4'ha)]);
                  for (forvar101 = (1'h0); (forvar101 < (2'h2)); forvar101 = (forvar101 + (1'h1)))
                    begin
                      reg102 <= ($signed($unsigned((reg40 > reg90))) >>> $signed(({reg57} ?
                          $unsigned((8'hb2)) : (-reg90))));
                    end
                  for (forvar103 = (1'h0); (forvar103 < (2'h3)); forvar103 = (forvar103 + (1'h1)))
                    begin
                      reg104 <= (8'hb6);
                    end
                end
              if ($signed($signed(($signed(forvar49) ?
                  reg39[(2'h3):(2'h3)] : ((8'ha0) <<< reg104)))))
                begin
                  if ($signed((((reg76 ? reg22 : reg26) ?
                          {forvar53} : $signed(forvar25)) ?
                      $signed(reg95[(3'h5):(2'h3)]) : ($unsigned(reg80) << ((8'hb3) <<< reg34)))))
                    begin
                      reg105 <= {((reg83[(1'h0):(1'h0)] ?
                                  reg89[(3'h7):(1'h1)] : (~&(8'hab))) ?
                              $signed(forvar20[(2'h3):(2'h2)]) : ((reg44 ?
                                  reg51 : reg17) >> (-reg44)))};
                      reg106 <= (!forvar82);
                    end
                  else
                    begin
                      reg105 <= (|$signed((reg43 <<< reg93)));
                    end
                  for (forvar107 = (1'h0); (forvar107 < (2'h2)); forvar107 = (forvar107 + (1'h1)))
                    begin
                      reg108 <= (reg34[(3'h7):(1'h1)] != (forvar67 ^~ reg82));
                      reg109 <= $signed(reg92);
                      reg110 <= ($signed((~^forvar107)) ?
                          (reg108 ?
                              reg73 : ((reg33 ? reg40 : reg104) + (reg105 ?
                                  reg38 : (8'hb5)))) : $unsigned($unsigned($signed(reg18))));
                      reg111 <= $unsigned({((|forvar31) ?
                              $signed((8'hb1)) : $unsigned(forvar40))});
                    end
                  for (forvar112 = (1'h0); (forvar112 < (1'h1)); forvar112 = (forvar112 + (1'h1)))
                    begin
                      reg113 <= $unsigned($unsigned($signed((8'h9c))));
                      reg114 <= reg79[(3'h4):(1'h1)];
                      reg115 <= reg39[(3'h4):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar105 = (1'h0); (forvar105 < (2'h3)); forvar105 = (forvar105 + (1'h1)))
                    begin
                      reg106 <= (~^forvar25[(3'h7):(2'h3)]);
                      reg107 <= (~|($unsigned((reg88 >> reg102)) << reg13[(3'h5):(1'h1)]));
                      reg108 <= $unsigned(reg26[(4'h8):(3'h4)]);
                      reg109 <= $unsigned(((forvar77 != (&reg17)) ~^ {forvar15}));
                    end
                  if (reg84[(2'h2):(2'h2)])
                    begin
                      reg110 <= $unsigned($unsigned((8'h9e)));
                      reg111 <= (((&((8'had) ?
                              (8'hba) : (8'h9c))) & reg33[(1'h1):(1'h0)]) ?
                          $signed(reg97) : $signed((^(reg26 * reg108))));
                      reg112 <= reg47;
                    end
                  else
                    begin
                      reg110 <= $unsigned((reg105 ?
                          $unsigned(reg70[(2'h2):(2'h2)]) : (8'hb6)));
                      reg111 <= forvar20[(3'h4):(3'h4)];
                    end
                end
            end
          else
            begin
              for (forvar99 = (1'h0); (forvar99 < (1'h0)); forvar99 = (forvar99 + (1'h1)))
                begin
                  if ($unsigned(forvar58))
                    begin
                      reg100 <= reg32;
                      reg101 <= $unsigned($unsigned((^$unsigned(reg47))));
                      reg102 <= ((reg78[(3'h6):(2'h2)] <= ((reg78 ?
                              forvar71 : reg109) << reg90)) ?
                          forvar11[(3'h6):(1'h1)] : ((&reg74) >= reg23));
                      reg103 <= reg70;
                    end
                  else
                    begin
                      reg100 <= $signed(forvar63);
                      reg101 <= $signed((forvar28 ~^ ((!forvar112) ^ (reg102 ?
                          reg88 : (8'hab)))));
                    end
                end
              for (forvar104 = (1'h0); (forvar104 < (2'h2)); forvar104 = (forvar104 + (1'h1)))
                begin
                  for (forvar105 = (1'h0); (forvar105 < (2'h3)); forvar105 = (forvar105 + (1'h1)))
                    begin
                      reg106 <= (~|({$signed((8'h9e))} == (forvar86[(4'h8):(3'h7)] | (reg114 ~^ (8'h9d)))));
                      reg107 <= reg98[(2'h3):(2'h2)];
                      reg108 <= (!(~|{(reg45 >>> reg102)}));
                    end
                  reg109 <= forvar99;
                  reg110 <= $unsigned((reg41[(2'h3):(1'h0)] ?
                      $signed((forvar53 << forvar74)) : ($signed(forvar71) != (^~forvar24))));
                end
            end
          for (forvar116 = (1'h0); (forvar116 < (2'h3)); forvar116 = (forvar116 + (1'h1)))
            begin
              if ($signed($signed(($unsigned(forvar103) | (forvar74 && reg70)))))
                begin
                  for (forvar117 = (1'h0); (forvar117 < (2'h3)); forvar117 = (forvar117 + (1'h1)))
                    begin
                      reg118 <= (8'hb2);
                      reg119 <= $unsigned(reg75[(2'h2):(1'h0)]);
                      reg120 <= ((~|((reg41 + reg60) >> ((8'ha8) ?
                          forvar28 : reg40))) >>> {reg70});
                      reg121 <= (8'hba);
                    end
                end
              else
                begin
                  for (forvar117 = (1'h0); (forvar117 < (1'h1)); forvar117 = (forvar117 + (1'h1)))
                    begin
                      reg118 <= reg19[(2'h3):(1'h0)];
                      reg119 <= {$unsigned($signed({reg39}))};
                      reg120 <= $signed((($unsigned(forvar62) ?
                          (reg85 ?
                              forvar82 : (8'hb5)) : (!reg102)) + $unsigned({(8'ha8)})));
                      reg121 <= ($signed($signed(reg52)) <= $signed({$unsigned(forvar112)}));
                    end
                end
              for (forvar122 = (1'h0); (forvar122 < (1'h0)); forvar122 = (forvar122 + (1'h1)))
                begin
                  for (forvar123 = (1'h0); (forvar123 < (2'h2)); forvar123 = (forvar123 + (1'h1)))
                    begin
                      reg124 <= (((^~(!reg23)) ?
                              (!reg16[(3'h7):(2'h3)]) : {$signed(reg27)}) ?
                          $unsigned((&(~|forvar78))) : ($unsigned(((8'hac) ?
                                  reg121 : reg52)) ?
                              $signed((forvar46 * reg54)) : (reg45[(3'h7):(1'h1)] ^~ forvar105)));
                    end
                  if (reg109[(1'h1):(1'h0)])
                    begin
                      reg125 <= $unsigned((~|{forvar20}));
                    end
                  else
                    begin
                      reg125 <= reg48[(4'ha):(4'ha)];
                      reg126 <= (&($unsigned($unsigned(reg36)) | (~^$signed(reg30))));
                      reg127 <= ((forvar53[(3'h4):(1'h1)] & {$unsigned(forvar46)}) ?
                          (forvar62[(2'h3):(2'h3)] < ({forvar31} ?
                              reg89[(4'h9):(3'h7)] : forvar91)) : reg42);
                    end
                end
              reg128 <= (reg26 ?
                  forvar41[(2'h2):(1'h0)] : reg103[(4'h8):(2'h2)]);
            end
        end
      else
        begin
          if ((forvar11 ~^ $signed(reg48[(3'h5):(3'h4)])))
            begin
              for (forvar99 = (1'h0); (forvar99 < (1'h0)); forvar99 = (forvar99 + (1'h1)))
                begin
                  if (reg32[(3'h6):(3'h5)])
                    begin
                      reg100 <= {reg120};
                      reg101 <= reg90[(3'h6):(3'h6)];
                      reg102 <= forvar61;
                      reg103 <= (forvar94[(1'h1):(1'h0)] << ((8'h9d) ?
                          $unsigned((forvar31 ?
                              reg93 : reg45)) : (~&$unsigned(forvar62))));
                    end
                  else
                    begin
                      reg100 <= ({$unsigned((8'ha4))} ^ ($unsigned((reg96 ?
                              forvar24 : (8'h9f))) ?
                          ($unsigned(reg111) <<< forvar117[(3'h4):(2'h3)]) : (|(|(8'ha5)))));
                      reg101 <= $signed(((forvar87[(2'h3):(2'h2)] <= (8'haf)) >= ((reg113 << reg79) > $unsigned(forvar62))));
                    end
                  reg104 <= (!$unsigned(reg127[(3'h4):(2'h2)]));
                  if (((&{(reg21 ? reg44 : forvar87)}) >= reg64))
                    begin
                      reg105 <= {reg13};
                      reg106 <= reg51;
                      reg107 <= $unsigned((^~$signed({(8'hb6)})));
                      reg108 <= (!forvar24[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg105 <= reg16[(4'ha):(4'ha)];
                      reg106 <= ((8'h9f) >>> $unsigned((forvar103[(3'h6):(3'h4)] ?
                          reg96 : reg64[(4'hb):(4'h8)])));
                      reg107 <= (^(8'hb9));
                      reg108 <= {forvar29[(2'h3):(2'h2)]};
                    end
                  for (forvar109 = (1'h0); (forvar109 < (2'h3)); forvar109 = (forvar109 + (1'h1)))
                    begin
                      reg110 <= ((forvar35 ?
                              reg124[(1'h0):(1'h0)] : {$signed(reg84)}) ?
                          reg27[(1'h1):(1'h0)] : reg124);
                      reg111 <= reg68;
                    end
                end
              for (forvar112 = (1'h0); (forvar112 < (2'h3)); forvar112 = (forvar112 + (1'h1)))
                begin
                  reg113 <= $signed($unsigned((((8'hac) ?
                      reg110 : reg18) | reg16)));
                end
            end
          else
            begin
              reg99 <= (reg89 >= reg43[(4'ha):(2'h3)]);
              if ((8'ha5))
                begin
                  if (($signed(reg118) << (8'ha0)))
                    begin
                      reg100 <= forvar40[(1'h0):(1'h0)];
                      reg101 <= $signed((forvar123[(1'h0):(1'h0)] >> {forvar29}));
                    end
                  else
                    begin
                      reg100 <= ({reg37[(3'h5):(2'h2)]} < forvar86);
                      reg101 <= ((((reg43 ? reg107 : reg36) > (reg104 ?
                          forvar104 : forvar107)) | (reg52 <<< {wire6})) & (~^((reg14 ?
                          reg82 : (8'hb5)) * (reg68 ? forvar40 : reg42))));
                      reg102 <= reg70[(2'h2):(2'h2)];
                      reg103 <= forvar41[(3'h7):(1'h1)];
                    end
                  reg104 <= $signed((8'hac));
                  if ({reg81[(4'h9):(3'h6)]})
                    begin
                      reg105 <= ((reg99[(3'h6):(2'h2)] >= forvar101) ?
                          {(~|(forvar20 ?
                                  reg111 : forvar53))} : $signed($signed(forvar86[(4'h9):(3'h7)])));
                      reg106 <= (^reg109[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg105 <= (!{{{reg103}}});
                    end
                end
              else
                begin
                  if (reg56)
                    begin
                      reg100 <= reg101[(1'h0):(1'h0)];
                      reg101 <= $unsigned(forvar78);
                      reg102 <= ((reg108 ?
                          reg56 : $signed($unsigned(forvar104))) << {$unsigned((forvar86 >= reg81))});
                    end
                  else
                    begin
                      reg100 <= ((^(8'hb2)) ? (~^reg100) : (!(~(!reg65))));
                      reg101 <= $unsigned((+$signed((reg54 ?
                          forvar116 : forvar20))));
                      reg102 <= reg40;
                    end
                  for (forvar103 = (1'h0); (forvar103 < (2'h3)); forvar103 = (forvar103 + (1'h1)))
                    begin
                      reg104 <= {(reg102[(2'h3):(2'h2)] >= (^~$unsigned(reg17)))};
                      reg105 <= $signed($unsigned(((reg36 <<< reg16) + (reg126 ?
                          forvar40 : forvar35))));
                      reg106 <= ((forvar94[(1'h1):(1'h1)] & $signed($unsigned((8'hb1)))) - reg51[(3'h7):(1'h1)]);
                    end
                end
              for (forvar107 = (1'h0); (forvar107 < (2'h2)); forvar107 = (forvar107 + (1'h1)))
                begin
                  for (forvar108 = (1'h0); (forvar108 < (1'h0)); forvar108 = (forvar108 + (1'h1)))
                    begin
                      reg109 <= (forvar58 ?
                          $unsigned($unsigned($unsigned(reg68))) : (reg21[(1'h0):(1'h0)] != $signed($unsigned(forvar107))));
                    end
                end
            end
          if ((+($signed($signed(reg90)) * $signed(reg68[(1'h0):(1'h0)]))))
            begin
              reg114 <= $unsigned($signed($signed((&reg60))));
              for (forvar115 = (1'h0); (forvar115 < (2'h2)); forvar115 = (forvar115 + (1'h1)))
                begin
                  for (forvar116 = (1'h0); (forvar116 < (1'h1)); forvar116 = (forvar116 + (1'h1)))
                    begin
                      reg117 <= ((^reg125) < {{(~^reg100)}});
                    end
                  reg118 <= ((reg77 ?
                          (reg85[(1'h1):(1'h1)] >> $signed(reg70)) : reg119) ?
                      $signed(reg57) : $unsigned(({forvar12} <= $unsigned(forvar123))));
                  if ({(8'had)})
                    begin
                      reg119 <= reg89[(1'h1):(1'h1)];
                      reg120 <= (8'ha6);
                      reg121 <= ((forvar101[(1'h1):(1'h1)] >> reg127) ?
                          {reg76[(2'h2):(1'h1)]} : forvar104[(4'hb):(4'h8)]);
                    end
                  else
                    begin
                      reg119 <= (~^reg66[(3'h4):(1'h1)]);
                      reg120 <= (~|((-reg120) == ($signed(reg98) ?
                          reg126 : $unsigned((8'haf)))));
                      reg121 <= (reg112[(2'h2):(1'h1)] ?
                          (($signed(forvar123) ?
                                  {forvar78} : (reg13 == (8'h9f))) ?
                              forvar24 : (reg54 ?
                                  $unsigned(reg54) : reg82)) : forvar29[(3'h5):(3'h4)]);
                    end
                  if ((forvar71 ?
                      $signed($unsigned(reg84)) : (~^(~^$unsigned(reg127)))))
                    begin
                      reg122 <= ((reg109 ?
                          $unsigned($unsigned(reg27)) : (+forvar117[(1'h0):(1'h0)])) <= (-{$unsigned(forvar101)}));
                      reg123 <= forvar78[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg122 <= (!reg69);
                      reg123 <= (|reg52[(3'h5):(2'h3)]);
                      reg124 <= (&$unsigned({(reg55 ? forvar40 : reg102)}));
                      reg125 <= ($unsigned($signed((|reg16))) ?
                          (^{((8'h9d) ?
                                  (8'had) : reg104)}) : $unsigned($signed((wire7 ^~ forvar49))));
                    end
                end
              if ($unsigned((8'h9c)))
                begin
                  reg126 <= reg102[(3'h4):(2'h2)];
                end
              else
                begin
                  reg126 <= reg102[(3'h7):(1'h1)];
                end
              if (($unsigned((~((8'hac) >> forvar11))) ?
                  {reg83[(1'h0):(1'h0)]} : ((forvar77 < (forvar72 ?
                          reg68 : reg106)) ?
                      (&forvar105[(1'h1):(1'h0)]) : ($unsigned(reg69) < reg70))))
                begin
                  for (forvar127 = (1'h0); (forvar127 < (1'h1)); forvar127 = (forvar127 + (1'h1)))
                    begin
                      reg128 <= ($unsigned((-$signed(reg54))) ?
                          ($signed($signed((8'ha9))) <<< $signed((^forvar72))) : $unsigned(((^~(8'hb5)) ?
                              $unsigned(reg13) : $unsigned(reg115))));
                      reg129 <= (reg123 ^ (~&((reg70 > reg51) ?
                          {reg69} : (8'ha0))));
                      reg130 <= $signed(forvar58[(1'h1):(1'h0)]);
                    end
                  reg131 <= $unsigned(forvar117[(1'h1):(1'h0)]);
                  if ({($unsigned({forvar11}) < (reg88[(3'h4):(1'h1)] ?
                          forvar116 : $signed((8'ha1))))})
                    begin
                      reg132 <= $unsigned($signed(reg76[(3'h4):(2'h2)]));
                      reg133 <= (!wire6[(2'h2):(2'h2)]);
                      reg134 <= wire9;
                      reg135 <= (^forvar58);
                    end
                  else
                    begin
                      reg132 <= reg114[(2'h3):(1'h0)];
                      reg133 <= (&reg90);
                    end
                end
              else
                begin
                  for (forvar127 = (1'h0); (forvar127 < (2'h2)); forvar127 = (forvar127 + (1'h1)))
                    begin
                      reg128 <= {{forvar86[(3'h4):(3'h4)]}};
                      reg129 <= (reg73[(1'h1):(1'h1)] < ((reg19[(1'h0):(1'h0)] != (forvar72 > (8'hb0))) != reg133[(4'hc):(4'h9)]));
                      reg130 <= (~|($unsigned({forvar31}) * (forvar41[(3'h4):(2'h2)] ?
                          {(8'hb0)} : $unsigned(reg93))));
                    end
                  for (forvar131 = (1'h0); (forvar131 < (2'h2)); forvar131 = (forvar131 + (1'h1)))
                    begin
                      reg132 <= reg22;
                      reg133 <= {((((8'h9d) + reg112) + reg54[(4'h9):(4'h9)]) * {$signed(forvar71)})};
                      reg134 <= reg90;
                      reg135 <= $unsigned((|$unsigned((reg131 ?
                          reg95 : forvar131))));
                    end
                end
            end
          else
            begin
              for (forvar114 = (1'h0); (forvar114 < (2'h3)); forvar114 = (forvar114 + (1'h1)))
                begin
                  for (forvar115 = (1'h0); (forvar115 < (2'h3)); forvar115 = (forvar115 + (1'h1)))
                    begin
                      reg116 <= (^{((8'ha5) ?
                              (reg98 ? forvar20 : reg105) : ((8'h9f) ?
                                  reg51 : forvar107))});
                      reg117 <= $signed((|(^$signed(reg21))));
                      reg118 <= reg56[(4'h8):(3'h7)];
                      reg119 <= $signed((((reg96 ? reg76 : reg30) ?
                          ((8'haa) ?
                              forvar104 : reg108) : reg60[(4'h9):(4'h9)]) >>> $signed((8'h9c))));
                    end
                  reg120 <= (-(forvar105[(1'h1):(1'h1)] ?
                      reg42[(2'h3):(2'h2)] : (8'ha8)));
                  for (forvar121 = (1'h0); (forvar121 < (1'h0)); forvar121 = (forvar121 + (1'h1)))
                    begin
                      reg122 <= ((reg122 <= $signed($signed(reg57))) ?
                          forvar12[(1'h0):(1'h0)] : ((reg75 <= reg80) ?
                              reg10 : ((forvar29 ?
                                  (8'ha7) : (8'hb1)) >> (forvar99 - forvar87))));
                      reg123 <= reg88[(3'h5):(1'h0)];
                      reg124 <= (forvar71 == (((&reg55) + forvar122[(4'he):(4'h8)]) || forvar29[(3'h6):(2'h2)]));
                    end
                end
              for (forvar125 = (1'h0); (forvar125 < (2'h2)); forvar125 = (forvar125 + (1'h1)))
                begin
                  if (reg21[(3'h5):(3'h5)])
                    begin
                      reg126 <= reg84;
                      reg127 <= forvar63[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg126 <= (8'hb2);
                      reg127 <= $unsigned(({reg43} ?
                          (+reg23[(2'h3):(1'h0)]) : forvar46[(1'h0):(1'h0)]));
                      reg128 <= ((forvar123 ?
                              (reg66 ?
                                  (~wire9) : forvar63) : ((reg127 <<< reg105) && (reg123 >> forvar117))) ?
                          {(~|(reg17 ?
                                  forvar107 : forvar105))} : $unsigned(reg52[(1'h0):(1'h0)]));
                    end
                  reg129 <= (~&$unsigned(reg108));
                  reg130 <= $unsigned($signed((!$signed((8'ha6)))));
                end
            end
          for (forvar136 = (1'h0); (forvar136 < (2'h2)); forvar136 = (forvar136 + (1'h1)))
            begin
              for (forvar137 = (1'h0); (forvar137 < (2'h2)); forvar137 = (forvar137 + (1'h1)))
                begin
                  for (forvar138 = (1'h0); (forvar138 < (2'h2)); forvar138 = (forvar138 + (1'h1)))
                    begin
                      reg139 <= reg42[(1'h0):(1'h0)];
                      reg140 <= $signed((~&$signed($signed(reg70))));
                      reg141 <= (($signed({reg115}) ?
                          $signed(reg89) : (&reg112[(1'h1):(1'h0)])) * $signed($unsigned(forvar63)));
                    end
                  reg142 <= reg48;
                  if ((~|$unsigned(((reg82 << reg109) >> $unsigned(forvar107)))))
                    begin
                      reg143 <= ($signed(($unsigned(reg142) ?
                              forvar12 : {(8'ha0)})) ?
                          forvar86[(2'h3):(2'h2)] : $signed(reg133[(4'ha):(2'h2)]));
                    end
                  else
                    begin
                      reg143 <= reg82;
                      reg144 <= $signed($unsigned(reg132[(2'h2):(1'h1)]));
                    end
                end
              if ($signed($signed(((|forvar82) ?
                  reg130[(1'h1):(1'h1)] : (&reg36)))))
                begin
                  for (forvar145 = (1'h0); (forvar145 < (2'h3)); forvar145 = (forvar145 + (1'h1)))
                    begin
                      reg146 <= {forvar29[(1'h1):(1'h0)]};
                      reg147 <= ($unsigned(reg18) >> reg124[(2'h3):(2'h2)]);
                      reg148 <= $signed({{reg75[(2'h2):(2'h2)]}});
                      reg149 <= ($unsigned($unsigned((forvar28 ?
                          forvar94 : reg65))) < forvar71);
                    end
                  if (((((~^forvar121) != (forvar35 >= forvar131)) << ((reg142 ?
                      reg140 : reg139) ^ (reg93 ? reg111 : wire9))) ^ (((reg17 ?
                          reg59 : forvar31) >= (reg14 <<< reg84)) ?
                      (((8'ha8) <= reg77) ?
                          (reg133 << reg126) : {reg105}) : reg90)))
                    begin
                      reg150 <= (-$unsigned($signed($unsigned(reg70))));
                      reg151 <= reg32;
                      reg152 <= ((~^reg22[(1'h1):(1'h1)]) ?
                          reg133[(4'h9):(1'h0)] : reg128[(3'h5):(2'h2)]);
                    end
                  else
                    begin
                      reg150 <= ({(^(reg148 + reg122))} ?
                          $unsigned(reg68) : forvar109);
                    end
                  for (forvar153 = (1'h0); (forvar153 < (1'h0)); forvar153 = (forvar153 + (1'h1)))
                    begin
                      reg154 <= $signed(reg65);
                      reg155 <= reg17;
                      reg156 <= $signed((8'ha7));
                      reg157 <= (forvar40[(1'h1):(1'h0)] > reg115[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  reg145 <= (|(~^(|$signed((8'hb2)))));
                  reg146 <= $unsigned(reg69[(3'h6):(3'h6)]);
                end
              for (forvar158 = (1'h0); (forvar158 < (2'h2)); forvar158 = (forvar158 + (1'h1)))
                begin
                  if (reg111)
                    begin
                      reg159 <= $unsigned((~forvar108));
                      reg160 <= $signed($unsigned({reg57[(4'h8):(2'h3)]}));
                      reg161 <= (reg133 + $signed((~|(forvar58 * reg41))));
                    end
                  else
                    begin
                      reg159 <= reg66;
                      reg160 <= reg41[(4'hb):(1'h1)];
                      reg161 <= ((($signed(forvar71) ?
                              $signed(reg122) : forvar138[(1'h0):(1'h0)]) ?
                          reg129 : $signed($unsigned(forvar153))) ^~ $signed((^~(forvar104 ?
                          reg97 : (8'hb1)))));
                    end
                end
            end
        end
      if ({({(~^(8'ha9))} + ((-wire6) || $unsigned(reg142)))})
        begin
          if ($signed($unsigned(((forvar20 >= reg18) ?
              forvar153[(1'h1):(1'h1)] : reg22))))
            begin
              for (forvar162 = (1'h0); (forvar162 < (2'h3)); forvar162 = (forvar162 + (1'h1)))
                begin
                  for (forvar163 = (1'h0); (forvar163 < (2'h2)); forvar163 = (forvar163 + (1'h1)))
                    begin
                      reg164 <= ((~^reg124) == forvar101);
                      reg165 <= reg65[(3'h7):(1'h1)];
                      reg166 <= reg146[(2'h3):(2'h3)];
                    end
                  for (forvar167 = (1'h0); (forvar167 < (1'h0)); forvar167 = (forvar167 + (1'h1)))
                    begin
                      reg168 <= ((((reg45 ?
                          (8'ha7) : reg134) >>> {forvar138}) ^~ forvar145[(2'h2):(1'h0)]) > reg128[(2'h2):(1'h0)]);
                      reg169 <= ($signed(($signed(reg101) ?
                          (reg99 >= reg154) : (reg39 | forvar103))) - (reg126[(3'h5):(3'h4)] != forvar78));
                      reg170 <= (&(~&$unsigned((~^reg157))));
                      reg171 <= (!($signed($unsigned(reg34)) ?
                          (reg54 >> (reg107 ? (8'hae) : (8'hb1))) : ((8'haf) ?
                              reg164 : (-wire6))));
                    end
                  for (forvar172 = (1'h0); (forvar172 < (1'h1)); forvar172 = (forvar172 + (1'h1)))
                    begin
                      reg173 <= (~|$signed($unsigned((forvar41 ?
                          reg103 : reg47))));
                      reg174 <= {(({(8'hab)} ? reg82 : $unsigned((8'hac))) ?
                              $unsigned($signed((8'hae))) : (reg68 ?
                                  {forvar20} : (^~reg157)))};
                    end
                end
              reg175 <= $signed($signed(forvar11[(3'h6):(2'h3)]));
              if ((~^(reg60[(1'h0):(1'h0)] & ($signed(wire7) ?
                  $signed((8'ha1)) : {reg68}))))
                begin
                  for (forvar176 = (1'h0); (forvar176 < (1'h0)); forvar176 = (forvar176 + (1'h1)))
                    begin
                      reg177 <= $unsigned(({reg69[(3'h5):(2'h2)]} ?
                          {reg106[(4'hd):(3'h6)]} : {reg154}));
                      reg178 <= (^~(($unsigned(reg19) <= {(8'ha3)}) + (reg36[(1'h0):(1'h0)] ?
                          (forvar77 ? reg70 : forvar122) : (^~reg154))));
                    end
                end
              else
                begin
                  for (forvar176 = (1'h0); (forvar176 < (2'h3)); forvar176 = (forvar176 + (1'h1)))
                    begin
                      reg177 <= (reg26 ? reg178 : forvar108[(3'h7):(1'h0)]);
                      reg178 <= ($signed(({reg38} ?
                          $signed(reg34) : $unsigned((8'hac)))) + ($unsigned(reg40[(1'h0):(1'h0)]) ?
                          reg106[(4'hc):(4'ha)] : $signed(reg151[(2'h3):(2'h2)])));
                      reg179 <= $signed({reg102});
                      reg180 <= (reg120[(1'h1):(1'h1)] != $signed(((-reg151) | {reg105})));
                    end
                  for (forvar181 = (1'h0); (forvar181 < (2'h2)); forvar181 = (forvar181 + (1'h1)))
                    begin
                      reg182 <= ($signed(reg14) ?
                          (reg100[(3'h7):(3'h6)] >> {(reg109 == forvar109)}) : {(reg139 ?
                                  $unsigned(reg88) : (~^forvar121))});
                      reg183 <= {(!$signed((reg39 ? reg166 : reg145)))};
                      reg184 <= ((+$signed(reg66[(4'hb):(3'h4)])) | forvar72[(1'h0):(1'h0)]);
                    end
                  for (forvar185 = (1'h0); (forvar185 < (1'h0)); forvar185 = (forvar185 + (1'h1)))
                    begin
                      reg186 <= ((forvar131 ?
                          (~^{reg112}) : forvar116) | {$unsigned(((8'hb4) > reg54))});
                      reg187 <= $signed(reg124);
                      reg188 <= (+$unsigned(($signed(reg78) ?
                          {forvar62} : reg113[(2'h2):(1'h0)])));
                    end
                  for (forvar189 = (1'h0); (forvar189 < (2'h2)); forvar189 = (forvar189 + (1'h1)))
                    begin
                      reg190 <= forvar137[(3'h6):(2'h3)];
                      reg191 <= ((reg183 ?
                          (forvar145[(1'h0):(1'h0)] * $signed(forvar11)) : reg146) == ((~(reg22 ?
                              (8'hb5) : (8'had))) ?
                          (8'ha9) : ($signed(reg13) ?
                              forvar71[(4'h8):(2'h2)] : (&reg146))));
                    end
                end
            end
          else
            begin
              if ($unsigned($unsigned(forvar181)))
                begin
                  if ($signed($unsigned(reg39[(3'h4):(1'h1)])))
                    begin
                      reg162 <= {((8'ha5) ? forvar53 : reg84[(3'h7):(3'h4)])};
                      reg163 <= reg128[(3'h5):(2'h2)];
                      reg164 <= reg76[(2'h2):(1'h1)];
                      reg165 <= $unsigned((((reg161 ?
                              (8'ha2) : reg106) != $signed((8'hba))) ?
                          $signed((~|reg23)) : $unsigned($unsigned(reg170))));
                    end
                  else
                    begin
                      reg162 <= $unsigned($unsigned($unsigned({forvar53})));
                    end
                  if (($signed(((reg134 ^~ forvar138) << ((8'hb1) ?
                      (8'h9f) : reg22))) > reg107[(4'he):(1'h0)]))
                    begin
                      reg166 <= reg129[(1'h0):(1'h0)];
                      reg167 <= $unsigned($signed((^$unsigned(reg42))));
                    end
                  else
                    begin
                      reg166 <= reg70;
                      reg167 <= (reg160 ^ reg19[(2'h2):(1'h1)]);
                    end
                  if ($unsigned((reg45[(2'h3):(2'h2)] ?
                      reg103 : ($unsigned(reg173) & {reg131}))))
                    begin
                      reg168 <= reg142;
                      reg169 <= ((reg143[(2'h2):(1'h1)] ?
                          reg179[(4'h8):(2'h2)] : $signed($unsigned((8'ha5)))) >= reg26[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg168 <= reg42;
                    end
                  reg170 <= ($unsigned($unsigned((!(8'ha5)))) <= $signed({$signed(reg120)}));
                end
              else
                begin
                  for (forvar162 = (1'h0); (forvar162 < (2'h3)); forvar162 = (forvar162 + (1'h1)))
                    begin
                      reg163 <= (!$signed(forvar61[(2'h2):(1'h1)]));
                    end
                end
            end
        end
      else
        begin
          if (((((reg76 || reg179) ? reg80 : $unsigned(reg188)) ?
              ((&(8'haa)) > forvar112) : $signed((forvar31 < (8'h9f)))) == ({reg97} ?
              $unsigned(reg123) : reg127[(2'h3):(1'h1)])))
            begin
              if (forvar40[(4'hc):(3'h5)])
                begin
                  if ($unsigned((reg106 ?
                      (reg131[(4'h8):(2'h2)] ?
                          (&forvar71) : (&reg65)) : (forvar137[(4'hd):(1'h0)] << (reg146 ?
                          reg57 : forvar189)))))
                    begin
                      reg162 <= (reg152 >= $signed(forvar116[(3'h6):(1'h0)]));
                    end
                  else
                    begin
                      reg162 <= ($unsigned($unsigned((reg51 >= reg48))) & $signed($signed(reg40[(2'h3):(1'h0)])));
                      reg163 <= $signed(reg113);
                    end
                  for (forvar164 = (1'h0); (forvar164 < (1'h1)); forvar164 = (forvar164 + (1'h1)))
                    begin
                      reg165 <= {(((reg54 ? reg147 : reg96) ?
                              ((8'ha2) ?
                                  reg41 : (8'h9e)) : $unsigned(reg68)) + {(forvar101 ~^ reg174)})};
                      reg166 <= (~|(reg169[(2'h2):(2'h2)] ^~ (reg69 ?
                          forvar12[(3'h7):(3'h4)] : reg64[(1'h0):(1'h0)])));
                    end
                  reg167 <= forvar24;
                end
              else
                begin
                  if ($unsigned(($signed((8'h9e)) >> (~&(reg128 ?
                      forvar136 : reg179)))))
                    begin
                      reg162 <= (~reg163);
                    end
                  else
                    begin
                      reg162 <= forvar72[(3'h4):(2'h3)];
                      reg163 <= ((~|{(|reg80)}) <= $unsigned((~(8'hb6))));
                      reg164 <= reg68;
                    end
                  if ((!reg10))
                    begin
                      reg165 <= ((((8'ha5) | (reg161 ? reg10 : (8'had))) ?
                          (forvar117 <<< (reg124 & (8'ha0))) : ({(8'h9d)} & $signed(forvar87))) ^ ((~|reg126[(2'h3):(1'h1)]) ?
                          $signed(reg119) : (reg178[(1'h1):(1'h0)] ?
                              forvar49 : (~^reg174))));
                      reg166 <= reg128;
                    end
                  else
                    begin
                      reg165 <= $signed((forvar109 - ((&reg52) >= reg182[(1'h0):(1'h0)])));
                      reg166 <= $unsigned($signed(reg108));
                      reg167 <= $signed($unsigned($signed((reg32 ?
                          forvar137 : reg45))));
                      reg168 <= $signed(reg74);
                    end
                  for (forvar169 = (1'h0); (forvar169 < (1'h1)); forvar169 = (forvar169 + (1'h1)))
                    begin
                      reg170 <= $unsigned(forvar169[(2'h2):(1'h0)]);
                      reg171 <= $unsigned($unsigned((((8'ha7) ?
                          reg110 : reg156) + {forvar185})));
                      reg172 <= $unsigned($signed($signed(((8'hae) ?
                          reg155 : reg151))));
                      reg173 <= (!(((+(8'hab)) == {reg182}) ?
                          $unsigned(reg169) : ((reg82 ? reg109 : reg97) ?
                              reg154[(2'h3):(2'h3)] : (-reg89))));
                    end
                  for (forvar174 = (1'h0); (forvar174 < (2'h2)); forvar174 = (forvar174 + (1'h1)))
                    begin
                      reg175 <= reg140;
                      reg176 <= $signed(reg47);
                    end
                end
            end
          else
            begin
              for (forvar162 = (1'h0); (forvar162 < (2'h3)); forvar162 = (forvar162 + (1'h1)))
                begin
                  for (forvar163 = (1'h0); (forvar163 < (2'h3)); forvar163 = (forvar163 + (1'h1)))
                    begin
                      reg164 <= $signed(reg17);
                      reg165 <= reg45;
                    end
                  for (forvar166 = (1'h0); (forvar166 < (2'h3)); forvar166 = (forvar166 + (1'h1)))
                    begin
                      reg167 <= ($unsigned($unsigned((&(8'h9f)))) ?
                          $signed((8'hb0)) : reg166[(1'h1):(1'h1)]);
                      reg168 <= reg120;
                      reg169 <= $unsigned($signed({reg64}));
                      reg170 <= $signed((8'ha8));
                    end
                  if (reg79[(4'hb):(2'h2)])
                    begin
                      reg171 <= $unsigned($signed(((reg142 ?
                          wire9 : forvar158) < (+forvar174))));
                      reg172 <= {reg140[(1'h0):(1'h0)]};
                      reg173 <= (~^{($signed(reg114) ?
                              forvar31[(3'h5):(1'h0)] : (reg125 ?
                                  reg54 : reg51))});
                    end
                  else
                    begin
                      reg171 <= (+$unsigned((((8'hab) ?
                          (8'hb3) : reg107) == reg147)));
                      reg172 <= (|reg145);
                      reg173 <= $signed(($signed({forvar82}) ?
                          $signed((~(8'hb6))) : $unsigned((reg80 + reg18))));
                    end
                end
              if (reg190[(4'ha):(1'h0)])
                begin
                  reg174 <= reg108[(1'h0):(1'h0)];
                  if (reg73[(2'h3):(2'h3)])
                    begin
                      reg175 <= (8'hb3);
                    end
                  else
                    begin
                      reg175 <= ((+(|reg120)) ~^ (8'hb9));
                      reg176 <= {$signed($unsigned((reg144 && forvar25)))};
                      reg177 <= reg171[(2'h3):(2'h3)];
                    end
                  if (reg159)
                    begin
                      reg178 <= forvar86;
                      reg179 <= ($signed((8'hb0)) ?
                          ($signed($unsigned((8'h9f))) ?
                              ((reg119 ? reg44 : (8'ha0)) ?
                                  (reg26 ?
                                      reg131 : reg80) : reg160) : $signed(forvar136[(4'h9):(2'h3)])) : reg33[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg178 <= {($unsigned(reg73) >>> reg85[(3'h5):(2'h3)])};
                      reg179 <= {(reg156 >>> ((reg191 ? forvar11 : reg184) ?
                              reg66 : reg54[(4'ha):(1'h1)]))};
                      reg180 <= $signed(reg187[(3'h6):(2'h3)]);
                    end
                end
              else
                begin
                  for (forvar174 = (1'h0); (forvar174 < (1'h1)); forvar174 = (forvar174 + (1'h1)))
                    begin
                      reg175 <= reg178;
                      reg176 <= (reg111 >= {$unsigned(forvar174)});
                      reg177 <= (8'hb0);
                    end
                end
              if ($signed($unsigned(reg19[(3'h5):(1'h0)])))
                begin
                  for (forvar181 = (1'h0); (forvar181 < (1'h0)); forvar181 = (forvar181 + (1'h1)))
                    begin
                      reg182 <= $unsigned(reg177[(2'h3):(2'h2)]);
                    end
                  reg183 <= (&$unsigned($unsigned($signed(reg184))));
                  reg184 <= reg152[(3'h4):(2'h2)];
                end
              else
                begin
                  for (forvar181 = (1'h0); (forvar181 < (1'h0)); forvar181 = (forvar181 + (1'h1)))
                    begin
                      reg182 <= ((forvar174 == reg44[(3'h5):(3'h4)]) ?
                          reg150[(1'h1):(1'h0)] : $unsigned(forvar105[(3'h5):(1'h1)]));
                    end
                end
            end
          reg185 <= (!{{$signed(reg98)}});
          if ((8'hb1))
            begin
              if ({((~^reg111[(1'h0):(1'h0)]) <<< (-(reg188 ^ (8'ha0))))})
                begin
                  for (forvar186 = (1'h0); (forvar186 < (1'h0)); forvar186 = (forvar186 + (1'h1)))
                    begin
                      reg187 <= (8'hb8);
                    end
                  if ($signed($signed(((&reg115) ?
                      (reg64 & forvar107) : reg160[(4'h9):(3'h6)]))))
                    begin
                      reg188 <= reg103[(3'h7):(2'h2)];
                    end
                  else
                    begin
                      reg188 <= (reg26[(4'he):(4'h8)] || {$unsigned((forvar116 ?
                              wire6 : (8'hb3)))});
                      reg189 <= forvar176;
                      reg190 <= ($unsigned($signed((reg117 ?
                          forvar46 : (8'haf)))) <= (8'had));
                    end
                  if (($unsigned($signed(reg167[(1'h1):(1'h0)])) * $signed(((forvar25 <<< forvar105) ?
                      (reg147 ^ reg107) : $unsigned(reg57)))))
                    begin
                      reg191 <= ((|{$signed(reg172)}) && (^~{$unsigned(forvar103)}));
                      reg192 <= (|((-$signed(forvar11)) <= $unsigned((+(8'ha7)))));
                      reg193 <= reg80[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg191 <= reg48[(2'h2):(2'h2)];
                      reg192 <= (&((8'h9e) >= $signed(reg51[(4'h9):(4'h9)])));
                    end
                  for (forvar194 = (1'h0); (forvar194 < (2'h2)); forvar194 = (forvar194 + (1'h1)))
                    begin
                      reg195 <= (^~(((!reg23) ?
                              (|forvar115) : (forvar31 ~^ reg163)) ?
                          forvar91 : {reg96}));
                    end
                end
              else
                begin
                  reg186 <= {((reg42 ? reg97 : $signed((8'had))) <<< forvar62)};
                end
            end
          else
            begin
              for (forvar186 = (1'h0); (forvar186 < (1'h0)); forvar186 = (forvar186 + (1'h1)))
                begin
                  for (forvar187 = (1'h0); (forvar187 < (2'h2)); forvar187 = (forvar187 + (1'h1)))
                    begin
                      reg188 <= reg119[(1'h1):(1'h1)];
                      reg189 <= reg100;
                      reg190 <= ((((!forvar107) & $signed(reg40)) ?
                              reg111[(3'h7):(1'h0)] : $unsigned(forvar99[(2'h2):(1'h0)])) ?
                          $unsigned(wire6[(3'h6):(2'h2)]) : reg13);
                    end
                end
              if (reg154[(3'h6):(3'h4)])
                begin
                  for (forvar191 = (1'h0); (forvar191 < (2'h3)); forvar191 = (forvar191 + (1'h1)))
                    begin
                      reg192 <= {$signed(((~&forvar186) ?
                              reg57[(4'h9):(4'h9)] : $signed(reg21)))};
                    end
                  for (forvar193 = (1'h0); (forvar193 < (2'h3)); forvar193 = (forvar193 + (1'h1)))
                    begin
                      reg194 <= forvar176;
                      reg195 <= $unsigned($signed(reg68[(3'h4):(1'h0)]));
                      reg196 <= reg13;
                    end
                  for (forvar197 = (1'h0); (forvar197 < (1'h1)); forvar197 = (forvar197 + (1'h1)))
                    begin
                      reg198 <= (($signed({reg142}) ?
                          (reg118[(2'h3):(1'h1)] ?
                              (reg23 ?
                                  (8'hba) : forvar72) : $unsigned(reg30)) : {(reg76 - reg41)}) * {forvar123[(1'h0):(1'h0)]});
                      reg199 <= (wire7[(3'h5):(3'h5)] ^ forvar35);
                      reg200 <= (($unsigned($signed(forvar194)) >= reg174) ?
                          $unsigned(((reg122 < wire9) ^ $signed(reg82))) : (8'hb4));
                      reg201 <= $signed($unsigned($unsigned({wire7})));
                    end
                end
              else
                begin
                  reg191 <= $unsigned(forvar67[(2'h3):(2'h3)]);
                  for (forvar192 = (1'h0); (forvar192 < (1'h1)); forvar192 = (forvar192 + (1'h1)))
                    begin
                      reg193 <= (reg192 ?
                          reg37 : $unsigned(reg43[(3'h6):(3'h6)]));
                      reg194 <= (forvar25 ?
                          {({forvar127} ?
                                  reg34 : (|reg196))} : reg111[(3'h6):(2'h3)]);
                    end
                  for (forvar195 = (1'h0); (forvar195 < (2'h2)); forvar195 = (forvar195 + (1'h1)))
                    begin
                      reg196 <= {$unsigned({reg168})};
                      reg197 <= ((~&($unsigned(forvar29) ?
                              $unsigned(reg93) : (forvar105 == reg178))) ?
                          ((reg142[(2'h3):(2'h3)] == reg159) ?
                              (&{reg23}) : $signed((forvar174 ?
                                  reg179 : reg160))) : $unsigned(reg162));
                      reg198 <= reg131;
                    end
                end
            end
          if ($signed((($signed(forvar91) << $unsigned(forvar29)) ?
              ((-reg54) ?
                  (reg90 ?
                      forvar11 : reg116) : forvar103[(1'h0):(1'h0)]) : {reg75})))
            begin
              if ((~&(((reg83 ^ reg113) ?
                  (reg165 & reg161) : (-reg93)) != {$unsigned(forvar122)})))
                begin
                  for (forvar202 = (1'h0); (forvar202 < (1'h0)); forvar202 = (forvar202 + (1'h1)))
                    begin
                      reg203 <= reg55;
                      reg204 <= $signed($signed(($unsigned(reg93) ^ forvar185[(3'h5):(3'h5)])));
                      reg205 <= reg142[(1'h1):(1'h1)];
                      reg206 <= (wire6 ~^ $signed(($signed(reg134) ?
                          (~^reg167) : (forvar35 ? reg121 : (8'ha1)))));
                    end
                  for (forvar207 = (1'h0); (forvar207 < (1'h1)); forvar207 = (forvar207 + (1'h1)))
                    begin
                      reg208 <= {(~$unsigned(reg13))};
                      reg209 <= (~^(8'hb5));
                      reg210 <= forvar103[(4'h8):(2'h3)];
                    end
                  reg211 <= reg84[(2'h2):(1'h1)];
                  if (reg191[(1'h0):(1'h0)])
                    begin
                      reg212 <= ((({reg21} ?
                              (~reg161) : reg157) * (~&reg81[(4'hd):(3'h5)])) ?
                          (&(^reg210)) : $unsigned(reg54));
                    end
                  else
                    begin
                      reg212 <= ({(reg132[(1'h1):(1'h0)] || reg156[(4'h8):(3'h5)])} ?
                          ({reg163[(1'h1):(1'h0)]} ?
                              ((reg163 ?
                                  reg114 : (8'hb3)) ~^ {reg102}) : (+{reg75})) : $signed($unsigned(reg182)));
                      reg213 <= $signed($signed(reg204));
                    end
                end
              else
                begin
                  for (forvar202 = (1'h0); (forvar202 < (1'h1)); forvar202 = (forvar202 + (1'h1)))
                    begin
                      reg203 <= (($unsigned((reg127 ? forvar185 : (8'hb0))) ?
                          $unsigned({reg188}) : ((^reg48) ?
                              $signed(forvar158) : (reg84 ?
                                  reg109 : forvar104))) >>> ((~&{forvar99}) ^ reg76));
                      reg204 <= $signed({reg155[(4'h9):(1'h1)]});
                    end
                  for (forvar205 = (1'h0); (forvar205 < (1'h1)); forvar205 = (forvar205 + (1'h1)))
                    begin
                      reg206 <= reg143;
                      reg207 <= reg60[(2'h2):(2'h2)];
                      reg208 <= (&(+(reg134 <<< reg32[(3'h5):(2'h3)])));
                      reg209 <= ((forvar122[(4'ha):(3'h6)] ?
                              reg207 : ((8'hb8) ^ {reg89})) ?
                          reg69[(2'h2):(2'h2)] : ((~|((8'hb5) ?
                              reg211 : reg135)) <= forvar94[(2'h2):(1'h0)]));
                    end
                end
              if ((reg123[(1'h0):(1'h0)] ?
                  reg54[(3'h7):(1'h0)] : (~^forvar24[(3'h4):(2'h2)])))
                begin
                  reg214 <= $unsigned({$signed((forvar138 ? reg39 : reg169))});
                  for (forvar215 = (1'h0); (forvar215 < (2'h3)); forvar215 = (forvar215 + (1'h1)))
                    begin
                      reg216 <= reg107;
                      reg217 <= (+reg70);
                      reg218 <= $unsigned($unsigned((reg109[(2'h2):(1'h1)] ?
                          (forvar99 && (8'hb1)) : $unsigned(reg133))));
                      reg219 <= $signed(reg117[(4'h8):(3'h4)]);
                    end
                end
              else
                begin
                  for (forvar214 = (1'h0); (forvar214 < (2'h3)); forvar214 = (forvar214 + (1'h1)))
                    begin
                      reg215 <= (&$unsigned({(~&reg211)}));
                      reg216 <= $signed(forvar117[(3'h4):(3'h4)]);
                      reg217 <= $unsigned($signed({(^forvar71)}));
                      reg218 <= reg120[(1'h1):(1'h1)];
                    end
                  for (forvar219 = (1'h0); (forvar219 < (2'h3)); forvar219 = (forvar219 + (1'h1)))
                    begin
                      reg220 <= reg219;
                      reg221 <= $signed(($unsigned($signed(reg148)) ?
                          (~^reg104[(1'h1):(1'h0)]) : (reg48[(4'h9):(1'h1)] - $signed(reg132))));
                      reg222 <= reg176;
                      reg223 <= $signed({reg145});
                    end
                  for (forvar224 = (1'h0); (forvar224 < (1'h0)); forvar224 = (forvar224 + (1'h1)))
                    begin
                      reg225 <= (reg26[(4'hd):(4'h8)] ?
                          (($unsigned((8'hb2)) ?
                              wire9[(1'h1):(1'h1)] : $signed(reg147)) & (reg197[(1'h0):(1'h0)] ?
                              reg42 : $unsigned(reg84))) : (reg111 ^ reg185));
                    end
                end
            end
          else
            begin
              if (reg195)
                begin
                  for (forvar202 = (1'h0); (forvar202 < (2'h3)); forvar202 = (forvar202 + (1'h1)))
                    begin
                      reg203 <= $unsigned(($signed(reg60) ^ {reg148}));
                      reg204 <= forvar41;
                      reg205 <= (|$unsigned((|$unsigned(forvar15))));
                      reg206 <= reg167[(3'h4):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar202 = (1'h0); (forvar202 < (1'h1)); forvar202 = (forvar202 + (1'h1)))
                    begin
                      reg203 <= forvar145[(2'h2):(1'h1)];
                      reg204 <= forvar121;
                    end
                  if (reg218[(1'h1):(1'h0)])
                    begin
                      reg205 <= ((8'hb4) + $unsigned($signed(forvar61[(3'h6):(3'h5)])));
                      reg206 <= (reg213 >>> (~&{$unsigned(reg169)}));
                      reg207 <= reg207;
                      reg208 <= (~(reg222[(4'h9):(2'h2)] == $signed((!forvar49))));
                    end
                  else
                    begin
                      reg205 <= $unsigned((((&reg69) || ((8'h9e) ?
                          (8'h9f) : reg111)) <<< reg152));
                    end
                  for (forvar209 = (1'h0); (forvar209 < (1'h0)); forvar209 = (forvar209 + (1'h1)))
                    begin
                      reg210 <= reg171;
                      reg211 <= $signed(($unsigned(reg218) ?
                          ((reg55 <<< reg69) != reg26[(3'h4):(3'h4)]) : $signed((reg184 | forvar193))));
                      reg212 <= ($signed({(!(8'hb9))}) > (reg45[(3'h4):(1'h0)] ?
                          ({reg54} ?
                              $signed(forvar181) : (reg22 - reg75)) : (~reg80[(4'hb):(2'h2)])));
                      reg213 <= forvar103[(4'h9):(4'h9)];
                    end
                end
              reg214 <= (+(reg192 << $signed($signed(forvar202))));
            end
        end
    end
  module226 #() modinst493 (.wire228(reg178), .y(wire492), .wire227(reg220), .wire231(reg13), .wire229(reg26), .clk(clk), .wire230(reg106));
  always
    @(posedge clk) begin
      if (reg77[(3'h6):(1'h0)])
        begin
          if (reg189)
            begin
              if ((((reg180 ^ $signed(reg102)) >> ($unsigned((8'h9c)) - reg113[(3'h7):(2'h3)])) ?
                  reg190[(1'h1):(1'h0)] : $unsigned((!$signed(reg73)))))
                begin
                  if (reg185[(2'h2):(1'h0)])
                    begin
                      reg494 <= reg162[(1'h1):(1'h0)];
                      reg495 <= (~^(&reg114));
                      reg496 <= (reg219[(3'h4):(3'h4)] < ($unsigned((&reg159)) >= $unsigned($signed(reg190))));
                      reg497 <= ($unsigned(reg219) >= $signed(reg179));
                    end
                  else
                    begin
                      reg494 <= (reg39 ?
                          (~|$unsigned((reg199 ?
                              (8'h9d) : reg200))) : (reg175[(3'h7):(1'h1)] <<< {(reg52 ?
                                  reg22 : reg211)}));
                    end
                end
              else
                begin
                  for (forvar494 = (1'h0); (forvar494 < (2'h3)); forvar494 = (forvar494 + (1'h1)))
                    begin
                      reg495 <= {{(~|reg198)}};
                      reg496 <= ($signed((|reg145)) != {($signed(reg92) ?
                              (reg80 * reg84) : reg159[(3'h4):(1'h1)])});
                    end
                  for (forvar497 = (1'h0); (forvar497 < (2'h2)); forvar497 = (forvar497 + (1'h1)))
                    begin
                      reg498 <= $unsigned((~^{(8'h9d)}));
                      reg499 <= reg144;
                    end
                end
              for (forvar500 = (1'h0); (forvar500 < (1'h0)); forvar500 = (forvar500 + (1'h1)))
                begin
                  for (forvar501 = (1'h0); (forvar501 < (2'h2)); forvar501 = (forvar501 + (1'h1)))
                    begin
                      reg502 <= reg130;
                      reg503 <= $signed(($signed({(8'hb2)}) <= ((reg144 ?
                              (8'hb2) : (8'haf)) ?
                          (reg221 || reg123) : $signed(reg177))));
                      reg504 <= reg502;
                    end
                end
              if ($signed((8'hb0)))
                begin
                  for (forvar505 = (1'h0); (forvar505 < (1'h1)); forvar505 = (forvar505 + (1'h1)))
                    begin
                      reg506 <= reg168;
                      reg507 <= $unsigned((reg502[(3'h4):(1'h1)] ?
                          (reg191[(4'hb):(4'ha)] ?
                              $unsigned(reg127) : $signed(reg40)) : $unsigned(forvar500)));
                      reg508 <= ($signed((|((8'haf) ? reg32 : (8'h9e)))) ?
                          $signed(reg104[(1'h0):(1'h0)]) : reg81);
                    end
                  for (forvar509 = (1'h0); (forvar509 < (2'h3)); forvar509 = (forvar509 + (1'h1)))
                    begin
                      reg510 <= (($signed(reg124[(2'h2):(1'h1)]) * reg56) - ((~^(reg76 ?
                              reg201 : reg177)) ?
                          (!(reg108 * reg195)) : reg199[(2'h2):(2'h2)]));
                      reg511 <= forvar501[(4'hd):(3'h7)];
                      reg512 <= reg185;
                      reg513 <= ($unsigned((~$signed(forvar505))) ?
                          $unsigned($signed((reg47 - reg186))) : ($unsigned($unsigned((8'hb7))) ?
                              reg131[(2'h3):(1'h1)] : $signed({reg503})));
                    end
                  for (forvar514 = (1'h0); (forvar514 < (2'h3)); forvar514 = (forvar514 + (1'h1)))
                    begin
                      reg515 <= $unsigned($unsigned((8'hb3)));
                    end
                end
              else
                begin
                  if ((!$signed($unsigned($unsigned(reg494)))))
                    begin
                      reg505 <= $signed((((reg32 ^ reg199) | reg52[(2'h2):(2'h2)]) - (8'h9d)));
                      reg506 <= $signed(wire8[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg505 <= (^~(-reg183[(4'h8):(1'h0)]));
                      reg506 <= ($unsigned((((8'ha1) ? reg73 : reg85) ?
                              $signed((8'ha7)) : $unsigned(reg52))) ?
                          (^$unsigned(((8'haa) - (8'hb4)))) : reg198[(1'h0):(1'h0)]);
                    end
                end
              for (forvar516 = (1'h0); (forvar516 < (1'h0)); forvar516 = (forvar516 + (1'h1)))
                begin
                  for (forvar517 = (1'h0); (forvar517 < (1'h1)); forvar517 = (forvar517 + (1'h1)))
                    begin
                      reg518 <= reg507;
                      reg519 <= (reg129[(3'h5):(2'h3)] == $unsigned(((-reg209) != $unsigned(reg145))));
                      reg520 <= (forvar494 ?
                          $unsigned((((8'ha0) << reg119) <= reg180)) : $signed(reg515[(3'h7):(3'h4)]));
                    end
                  if ($unsigned($unsigned(($unsigned(reg150) ?
                      $unsigned(forvar516) : reg142))))
                    begin
                      reg521 <= (reg195 ?
                          $unsigned((8'h9d)) : $unsigned($unsigned((~^reg64))));
                      reg522 <= {reg10};
                      reg523 <= reg70;
                      reg524 <= $signed($unsigned(reg161));
                    end
                  else
                    begin
                      reg521 <= (~|((reg218[(1'h1):(1'h0)] && $signed(reg109)) ~^ ($signed(reg70) ?
                          (reg151 ^~ reg155) : {reg511})));
                      reg522 <= $unsigned(reg511[(4'hd):(3'h4)]);
                    end
                end
            end
          else
            begin
              for (forvar494 = (1'h0); (forvar494 < (1'h1)); forvar494 = (forvar494 + (1'h1)))
                begin
                  for (forvar495 = (1'h0); (forvar495 < (1'h0)); forvar495 = (forvar495 + (1'h1)))
                    begin
                      reg496 <= $unsigned((($signed(reg33) ?
                              (reg82 ? forvar509 : reg148) : ((8'ha3) ?
                                  reg497 : reg521)) ?
                          {(reg47 ? reg194 : reg114)} : reg51));
                      reg497 <= reg185[(3'h7):(3'h4)];
                    end
                end
            end
          for (forvar525 = (1'h0); (forvar525 < (2'h3)); forvar525 = (forvar525 + (1'h1)))
            begin
              for (forvar526 = (1'h0); (forvar526 < (2'h3)); forvar526 = (forvar526 + (1'h1)))
                begin
                  if (((8'hae) ?
                      $signed((((8'h9f) ^ reg51) * reg17[(4'hd):(3'h5)])) : reg93))
                    begin
                      reg527 <= $unsigned((((reg99 ? reg101 : (8'hb8)) ?
                          $signed((8'ha9)) : (reg495 == reg70)) < $signed($unsigned(reg217))));
                      reg528 <= reg69;
                    end
                  else
                    begin
                      reg527 <= ($unsigned(((reg119 ~^ reg518) != reg38[(1'h0):(1'h0)])) ?
                          ((~&(reg75 ^ reg156)) && $unsigned((reg220 - reg77))) : reg126);
                      reg528 <= (+reg98);
                    end
                  reg529 <= (((&{reg96}) ?
                          {(^~reg167)} : ($signed(reg76) && (reg173 < forvar516))) ?
                      {((reg54 ? reg499 : reg37) ?
                              (reg125 ?
                                  reg139 : reg19) : (~&reg148))} : (^~({reg22} * forvar501[(2'h3):(2'h2)])));
                end
            end
          if ((~^reg172[(2'h2):(1'h0)]))
            begin
              if ((reg159[(1'h1):(1'h0)] ?
                  reg84[(4'ha):(4'h9)] : reg216[(2'h3):(1'h1)]))
                begin
                  reg530 <= $unsigned((~&$unsigned(reg99)));
                  if ((8'had))
                    begin
                      reg531 <= $signed(reg216);
                      reg532 <= (reg113 ?
                          ($unsigned($unsigned(reg522)) ?
                              $unsigned(reg125) : (reg520[(2'h2):(1'h1)] && $signed(reg148))) : (|$signed((8'h9d))));
                      reg533 <= reg106;
                    end
                  else
                    begin
                      reg531 <= reg215;
                      reg532 <= (-$signed((^~$signed(reg66))));
                      reg533 <= $unsigned($signed((reg193[(2'h3):(1'h0)] + ((8'ha7) ^~ (8'ha5)))));
                    end
                end
              else
                begin
                  if (reg497)
                    begin
                      reg530 <= reg193[(3'h7):(3'h5)];
                      reg531 <= reg171[(2'h3):(2'h3)];
                      reg532 <= reg168[(1'h0):(1'h0)];
                      reg533 <= ((((-reg98) ^~ (reg100 ? (8'hb1) : reg88)) ?
                          $signed($unsigned(reg183)) : reg57) >> reg13[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg530 <= reg206;
                    end
                  if ($unsigned((8'hae)))
                    begin
                      reg534 <= (reg110[(4'h8):(3'h6)] <<< ((|(|reg518)) ?
                          reg148[(3'h7):(2'h2)] : (&reg122[(2'h3):(1'h1)])));
                      reg535 <= (^({(^~reg106)} ?
                          $signed((~^forvar525)) : $unsigned($unsigned(reg93))));
                      reg536 <= $unsigned((((~(8'hb3)) | (!reg171)) < reg180[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg534 <= {reg208};
                      reg535 <= reg104;
                      reg536 <= (($unsigned(reg173[(1'h1):(1'h0)]) ?
                          (~$signed(reg177)) : {$signed((8'h9d))}) >> ((forvar501 == $signed((8'ha5))) == reg44[(4'h9):(4'h9)]));
                    end
                  if (reg150[(3'h5):(1'h0)])
                    begin
                      reg537 <= (~&$signed($signed($unsigned(reg64))));
                      reg538 <= (reg167 ? reg519 : {reg185});
                      reg539 <= ({wire7[(1'h0):(1'h0)]} ?
                          ($unsigned((reg64 | reg165)) ?
                              {{reg105}} : $signed(reg99)) : $unsigned((-(|reg199))));
                      reg540 <= (($unsigned((~^reg508)) < {$signed((8'ha8))}) ?
                          reg95 : reg149[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg537 <= reg219;
                      reg538 <= $unsigned((|reg190));
                      reg539 <= $signed((($signed(reg129) ?
                          (^reg152) : (~|forvar497)) == reg223[(2'h3):(1'h0)]));
                    end
                end
              for (forvar541 = (1'h0); (forvar541 < (2'h3)); forvar541 = (forvar541 + (1'h1)))
                begin
                  for (forvar542 = (1'h0); (forvar542 < (1'h1)); forvar542 = (forvar542 + (1'h1)))
                    begin
                      reg543 <= reg185;
                      reg544 <= $unsigned(reg168);
                    end
                  for (forvar545 = (1'h0); (forvar545 < (1'h1)); forvar545 = (forvar545 + (1'h1)))
                    begin
                      reg546 <= reg27[(1'h0):(1'h0)];
                      reg547 <= $unsigned({{((8'haf) ? reg191 : reg164)}});
                      reg548 <= {reg43[(3'h5):(2'h3)]};
                    end
                end
              for (forvar549 = (1'h0); (forvar549 < (1'h0)); forvar549 = (forvar549 + (1'h1)))
                begin
                  for (forvar550 = (1'h0); (forvar550 < (2'h2)); forvar550 = (forvar550 + (1'h1)))
                    begin
                      reg551 <= $unsigned(((8'hb8) - $signed($signed(reg141))));
                      reg552 <= $signed($signed(reg79[(3'h5):(1'h1)]));
                      reg553 <= reg173;
                      reg554 <= $signed(reg524[(1'h1):(1'h1)]);
                    end
                  if ((reg22 ?
                      $signed(((reg160 ? reg197 : reg190) ?
                          (reg107 ?
                              reg85 : reg19) : reg113)) : reg194[(3'h4):(3'h4)]))
                    begin
                      reg555 <= {{$signed((^reg117))}};
                      reg556 <= (((reg513 + (reg76 ? reg536 : reg82)) ?
                              (-(reg515 * (8'hae))) : $unsigned($unsigned(reg196))) ?
                          $unsigned(reg505) : reg161[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg555 <= $unsigned(reg44);
                      reg556 <= {$signed({(|reg107)})};
                      reg557 <= ({$signed(((8'ha5) & reg129))} != (reg32 ?
                          $signed($signed((8'hba))) : {reg547[(3'h4):(2'h3)]}));
                      reg558 <= $signed($signed(reg92));
                    end
                  if ((reg140 ?
                      {(&((8'ha6) ~^ reg222))} : (($unsigned(wire9) ?
                          $unsigned(reg513) : (reg499 ?
                              reg64 : reg180)) > ({(8'ha8)} ^~ reg203[(4'hb):(2'h3)]))))
                    begin
                      reg559 <= ($signed({{reg39}}) < (~&reg64[(4'hc):(3'h5)]));
                      reg560 <= $unsigned({$signed((~|reg84))});
                    end
                  else
                    begin
                      reg559 <= $signed(reg148);
                      reg560 <= reg556;
                    end
                  if ($signed($signed((~&reg125[(3'h4):(1'h1)]))))
                    begin
                      reg561 <= $unsigned(reg175[(4'h9):(3'h7)]);
                      reg562 <= reg120[(4'hc):(1'h1)];
                      reg563 <= ((((&reg106) != $signed(reg498)) ?
                              (reg82[(4'ha):(3'h7)] << forvar516) : reg529[(1'h1):(1'h0)]) ?
                          $signed(reg14[(4'h9):(2'h3)]) : ((&(&reg205)) ?
                              $signed($unsigned(reg527)) : {reg50[(1'h0):(1'h0)]}));
                      reg564 <= reg209;
                    end
                  else
                    begin
                      reg561 <= $unsigned($signed(($unsigned(reg10) * (reg64 ?
                          reg193 : (8'hb5)))));
                    end
                end
              if (($signed($unsigned($signed(reg209))) ?
                  (($unsigned(reg164) ~^ (~^reg177)) >> $unsigned($unsigned(reg494))) : ((+(reg171 ^ (8'h9c))) >> ((8'h9d) > (reg131 & reg142)))))
                begin
                  if ($signed($unsigned(((-(8'hb9)) << reg519))))
                    begin
                      reg565 <= ($signed($unsigned((forvar495 != reg183))) < reg174[(2'h3):(2'h2)]);
                      reg566 <= $signed(((reg121[(4'h8):(2'h3)] != reg508[(2'h2):(1'h0)]) & $unsigned(reg163)));
                    end
                  else
                    begin
                      reg565 <= ($unsigned($unsigned({reg554})) && (reg52 == $unsigned((~^(8'hac)))));
                      reg566 <= (forvar545[(3'h7):(3'h6)] ?
                          reg165[(2'h3):(1'h0)] : $signed(((!reg162) * $unsigned((8'h9f)))));
                    end
                  if ((8'ha9))
                    begin
                      reg567 <= ((reg80 ?
                          (~^$unsigned(reg546)) : wire8[(2'h2):(2'h2)]) || $signed((reg212[(1'h0):(1'h0)] ?
                          $unsigned(reg43) : (reg213 ? reg537 : reg191))));
                      reg568 <= (~&reg220);
                      reg569 <= ($unsigned(reg540) ? reg83 : (8'h9f));
                      reg570 <= {$unsigned((8'hb5))};
                    end
                  else
                    begin
                      reg567 <= $signed(reg104);
                      reg568 <= reg133[(4'h8):(4'h8)];
                    end
                end
              else
                begin
                  reg565 <= $signed($unsigned((&$unsigned(reg523))));
                end
            end
          else
            begin
              for (forvar530 = (1'h0); (forvar530 < (2'h3)); forvar530 = (forvar530 + (1'h1)))
                begin
                  for (forvar531 = (1'h0); (forvar531 < (2'h2)); forvar531 = (forvar531 + (1'h1)))
                    begin
                      reg532 <= reg149[(3'h7):(1'h0)];
                      reg533 <= (&reg561[(4'hc):(3'h6)]);
                      reg534 <= reg185;
                      reg535 <= $unsigned(reg45);
                    end
                end
              if ((($unsigned(forvar525) && $signed((reg116 ?
                  reg146 : reg557))) != ((8'ha2) * reg192[(2'h3):(2'h2)])))
                begin
                  if ((|$signed({(~(8'h9c))})))
                    begin
                      reg536 <= reg89[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg536 <= (!reg18);
                      reg537 <= $signed(reg174[(1'h0):(1'h0)]);
                      reg538 <= (^reg122);
                    end
                  if ({(^($signed(reg56) == forvar549))})
                    begin
                      reg539 <= ($unsigned(reg150) ?
                          reg80[(1'h0):(1'h0)] : $unsigned((-forvar495)));
                      reg540 <= $unsigned((!{(~reg121)}));
                      reg541 <= reg171;
                    end
                  else
                    begin
                      reg539 <= (reg568[(1'h1):(1'h1)] ?
                          (8'ha1) : ((~(reg141 ? (8'hba) : reg498)) ?
                              $signed($unsigned(reg520)) : (reg178 ?
                                  reg214[(1'h1):(1'h0)] : reg81)));
                      reg540 <= reg532[(1'h1):(1'h1)];
                      reg541 <= reg156[(3'h5):(3'h4)];
                    end
                  if ($signed((~|(~&(^(8'had))))))
                    begin
                      reg542 <= reg23[(4'h8):(2'h2)];
                      reg543 <= (~&reg17);
                    end
                  else
                    begin
                      reg542 <= (((&$signed(reg570)) <<< {$unsigned(reg132)}) >= reg99);
                      reg543 <= (((~&(~|reg510)) ?
                          reg105 : (forvar541 ^ {reg139})) > (reg174[(2'h3):(2'h2)] + ((forvar497 | reg176) ?
                          (~forvar549) : {reg515})));
                      reg544 <= ($unsigned($signed(((8'ha1) >= reg112))) ?
                          reg157 : ($unsigned(((8'ha4) <= reg143)) ^~ reg510));
                    end
                end
              else
                begin
                  for (forvar536 = (1'h0); (forvar536 < (2'h2)); forvar536 = (forvar536 + (1'h1)))
                    begin
                      reg537 <= $unsigned($signed($signed(((8'h9d) ^ reg44))));
                    end
                  if ((8'ha5))
                    begin
                      reg538 <= reg159;
                      reg539 <= reg171;
                      reg540 <= $signed({$unsigned(forvar549)});
                    end
                  else
                    begin
                      reg538 <= $unsigned($signed(((|reg538) ^ wire492)));
                      reg539 <= ((8'h9d) ?
                          (~&((reg192 ? reg180 : reg77) ?
                              reg540[(1'h0):(1'h0)] : reg505[(1'h1):(1'h0)])) : reg197);
                      reg540 <= (reg206[(2'h3):(1'h0)] ?
                          $unsigned($signed((reg512 ?
                              reg184 : forvar497))) : {{$unsigned(reg546)}});
                      reg541 <= reg55[(2'h2):(2'h2)];
                    end
                  if ($unsigned({(+reg103)}))
                    begin
                      reg542 <= $unsigned((reg522 | (^~{reg165})));
                    end
                  else
                    begin
                      reg542 <= ((-reg223) ?
                          (~reg197) : (($unsigned(reg54) ?
                              $unsigned((8'hb7)) : (~reg558)) || reg207));
                      reg543 <= reg174;
                      reg544 <= (reg89[(3'h7):(3'h4)] ?
                          {reg82[(4'hb):(3'h5)]} : ($signed($unsigned(reg495)) ?
                              $signed((!reg37)) : (-reg51)));
                    end
                end
              reg545 <= (forvar509 ?
                  reg13 : $unsigned($unsigned($unsigned(reg568))));
            end
        end
      else
        begin
          for (forvar494 = (1'h0); (forvar494 < (2'h2)); forvar494 = (forvar494 + (1'h1)))
            begin
              reg495 <= (~^(+($signed(reg48) > (reg225 ? forvar509 : reg64))));
              if ($unsigned($signed((8'hb9))))
                begin
                  reg496 <= reg538[(5'h10):(4'hb)];
                  for (forvar497 = (1'h0); (forvar497 < (2'h2)); forvar497 = (forvar497 + (1'h1)))
                    begin
                      reg498 <= reg69[(2'h2):(1'h0)];
                      reg499 <= $unsigned(($signed((forvar500 >> reg563)) ?
                          reg151[(3'h6):(3'h6)] : (reg64 ?
                              (wire7 ? (8'haf) : forvar545) : reg123)));
                      reg500 <= (reg547[(3'h4):(2'h2)] ?
                          ((reg537 ?
                                  $unsigned(reg69) : ((8'hb7) ?
                                      reg503 : reg215)) ?
                              forvar541[(3'h4):(1'h1)] : ($unsigned(reg225) ?
                                  reg111 : $unsigned((8'h9c)))) : reg534);
                      reg501 <= reg82[(3'h6):(1'h0)];
                    end
                  for (forvar502 = (1'h0); (forvar502 < (2'h2)); forvar502 = (forvar502 + (1'h1)))
                    begin
                      reg503 <= (^~(8'hae));
                      reg504 <= {(!((reg80 != reg120) || (+(8'hb5))))};
                      reg505 <= (((&reg105) == $signed((8'hb1))) ?
                          $unsigned(reg184[(3'h4):(1'h0)]) : (reg48[(2'h2):(1'h0)] ^~ $signed(reg134[(3'h5):(3'h4)])));
                    end
                end
              else
                begin
                  for (forvar496 = (1'h0); (forvar496 < (1'h1)); forvar496 = (forvar496 + (1'h1)))
                    begin
                      reg497 <= reg120[(4'hf):(2'h3)];
                      reg498 <= $signed({($signed(reg22) ? (8'haa) : {reg59})});
                    end
                  for (forvar499 = (1'h0); (forvar499 < (2'h3)); forvar499 = (forvar499 + (1'h1)))
                    begin
                      reg500 <= $unsigned((~|((!reg524) - (reg223 >= reg538))));
                    end
                  if ({$signed(reg513[(2'h2):(2'h2)])})
                    begin
                      reg501 <= reg533[(3'h5):(2'h2)];
                      reg502 <= (^~reg70);
                      reg503 <= reg495;
                      reg504 <= $signed(reg547);
                    end
                  else
                    begin
                      reg501 <= (^$unsigned({reg214}));
                      reg502 <= ($signed((reg76 ?
                              reg533 : reg30[(1'h0):(1'h0)])) ?
                          reg205 : ($unsigned(reg14[(4'hd):(4'ha)]) ?
                              reg102 : {$signed(reg133)}));
                      reg503 <= (~^reg139);
                    end
                  for (forvar505 = (1'h0); (forvar505 < (1'h1)); forvar505 = (forvar505 + (1'h1)))
                    begin
                      reg506 <= $signed(reg135[(1'h1):(1'h1)]);
                      reg507 <= (reg527[(1'h0):(1'h0)] ?
                          (((reg208 ? reg496 : reg77) ?
                              $signed(reg558) : reg551) < (~|(reg513 ?
                              reg73 : reg190))) : reg125);
                    end
                end
            end
          for (forvar508 = (1'h0); (forvar508 < (2'h2)); forvar508 = (forvar508 + (1'h1)))
            begin
              reg509 <= (reg201[(1'h0):(1'h0)] ?
                  ($unsigned($unsigned(reg506)) ?
                      (|(!reg162)) : $signed(reg498)) : ({$signed(reg32)} ?
                      $signed(reg77[(4'h8):(1'h1)]) : reg65));
            end
          if (reg102)
            begin
              for (forvar510 = (1'h0); (forvar510 < (2'h3)); forvar510 = (forvar510 + (1'h1)))
                begin
                  if ((~|reg125[(3'h5):(2'h3)]))
                    begin
                      reg511 <= $signed(reg102);
                      reg512 <= $unsigned(({(wire6 < reg191)} >> $signed((reg115 ?
                          reg19 : reg129))));
                      reg513 <= $unsigned(((-$signed(reg552)) >= {$signed(forvar536)}));
                    end
                  else
                    begin
                      reg511 <= $unsigned(reg520);
                    end
                  for (forvar514 = (1'h0); (forvar514 < (2'h2)); forvar514 = (forvar514 + (1'h1)))
                    begin
                      reg515 <= (+($unsigned(reg523[(4'hb):(3'h5)]) ?
                          $unsigned($unsigned(reg155)) : $signed($signed(reg535))));
                    end
                end
              for (forvar516 = (1'h0); (forvar516 < (2'h3)); forvar516 = (forvar516 + (1'h1)))
                begin
                  if ((~&$signed(reg217[(2'h3):(1'h1)])))
                    begin
                      reg517 <= reg100[(4'h9):(3'h4)];
                      reg518 <= reg195[(1'h1):(1'h0)];
                      reg519 <= (reg16[(4'h9):(3'h7)] < $unsigned((reg499 <<< (8'ha8))));
                    end
                  else
                    begin
                      reg517 <= $signed($unsigned($unsigned((8'ha0))));
                      reg518 <= $unsigned(($unsigned(reg541) ?
                          reg541 : reg570));
                      reg519 <= ($unsigned(($unsigned((8'ha6)) & reg116[(3'h4):(3'h4)])) >> reg508[(3'h5):(2'h2)]);
                    end
                  for (forvar520 = (1'h0); (forvar520 < (1'h1)); forvar520 = (forvar520 + (1'h1)))
                    begin
                      reg521 <= (reg77[(4'h8):(1'h1)] ?
                          {reg540[(2'h2):(2'h2)]} : $unsigned(($signed(reg515) ?
                              {(8'hb3)} : reg559[(1'h1):(1'h0)])));
                      reg522 <= (($unsigned(forvar497) <= ({reg148} ?
                              reg515[(2'h3):(2'h3)] : (8'hae))) ?
                          ($unsigned($unsigned(reg122)) != reg116) : (~&reg168[(4'hb):(2'h3)]));
                      reg523 <= reg495[(1'h1):(1'h1)];
                    end
                end
              for (forvar524 = (1'h0); (forvar524 < (2'h3)); forvar524 = (forvar524 + (1'h1)))
                begin
                  for (forvar525 = (1'h0); (forvar525 < (2'h3)); forvar525 = (forvar525 + (1'h1)))
                    begin
                      reg526 <= (forvar549 && reg123);
                      reg527 <= reg211[(4'hd):(1'h0)];
                    end
                  if ($unsigned($signed($unsigned((reg541 ?
                      reg211 : (8'hae))))))
                    begin
                      reg528 <= {$unsigned(reg78[(3'h5):(2'h2)])};
                      reg529 <= $unsigned(reg191[(2'h2):(1'h0)]);
                      reg530 <= reg51[(2'h2):(1'h0)];
                      reg531 <= $signed((8'hac));
                    end
                  else
                    begin
                      reg528 <= $signed((&reg502));
                      reg529 <= reg13;
                      reg530 <= (($signed({(8'hb6)}) <<< (forvar500 ?
                          (8'h9e) : $unsigned(reg507))) << $signed(((8'hb1) + reg85)));
                      reg531 <= $unsigned(reg504);
                    end
                end
            end
          else
            begin
              reg510 <= reg96[(1'h0):(1'h0)];
              if ((($unsigned($signed((8'h9f))) >>> (reg141 >= $unsigned((8'hb8)))) ^ $signed($signed($signed(reg103)))))
                begin
                  for (forvar511 = (1'h0); (forvar511 < (2'h2)); forvar511 = (forvar511 + (1'h1)))
                    begin
                      reg512 <= {$unsigned(reg166[(1'h1):(1'h0)])};
                    end
                  if ((~&($unsigned($unsigned(reg38)) ?
                      {(!reg507)} : ((+reg192) ?
                          $signed(reg73) : (~&(8'ha6))))))
                    begin
                      reg513 <= reg13[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg513 <= (reg212 || $unsigned(($unsigned(reg112) * {(8'hb1)})));
                      reg514 <= ($unsigned($signed($unsigned((8'hae)))) * forvar516);
                      reg515 <= forvar508;
                    end
                  for (forvar516 = (1'h0); (forvar516 < (2'h3)); forvar516 = (forvar516 + (1'h1)))
                    begin
                      reg517 <= ($unsigned(((forvar499 * (8'hb4)) | {reg510})) ^ reg534);
                      reg518 <= $unsigned(reg50[(1'h1):(1'h0)]);
                    end
                  for (forvar519 = (1'h0); (forvar519 < (2'h3)); forvar519 = (forvar519 + (1'h1)))
                    begin
                      reg520 <= reg45[(4'hd):(2'h2)];
                      reg521 <= (^(-((reg174 << reg199) + ((8'h9c) ^ reg552))));
                      reg522 <= (8'hb1);
                      reg523 <= (~&($signed((reg195 ?
                          reg215 : reg89)) | $signed((reg142 ~^ reg192))));
                    end
                end
              else
                begin
                  reg511 <= {$signed($signed((reg569 + (8'ha8))))};
                  for (forvar512 = (1'h0); (forvar512 < (1'h1)); forvar512 = (forvar512 + (1'h1)))
                    begin
                      reg513 <= $unsigned($unsigned((!(reg495 << reg132))));
                      reg514 <= ($unsigned(reg98[(1'h1):(1'h0)]) * wire7[(3'h5):(3'h4)]);
                      reg515 <= $unsigned(reg152[(1'h1):(1'h0)]);
                      reg516 <= ({($signed(reg211) * reg172)} << (($signed(forvar500) ?
                              reg197[(3'h6):(3'h6)] : (reg562 ?
                                  (8'h9c) : (8'hba))) ?
                          reg113 : ((forvar524 ? wire7 : reg495) ?
                              $unsigned((8'hb7)) : $unsigned((8'ha2)))));
                    end
                end
              if ((8'hb9))
                begin
                  for (forvar524 = (1'h0); (forvar524 < (1'h0)); forvar524 = (forvar524 + (1'h1)))
                    begin
                      reg525 <= reg215;
                      reg526 <= ((reg139 >>> (8'ha1)) ?
                          ($unsigned($unsigned(reg535)) ^~ (reg521 ?
                              (wire7 | reg80) : reg562)) : reg78[(3'h4):(2'h3)]);
                      reg527 <= $signed($unsigned($signed(reg22[(3'h6):(3'h6)])));
                      reg528 <= (~&(!(!{reg510})));
                    end
                end
              else
                begin
                  reg524 <= ($unsigned($signed(reg34[(3'h4):(2'h2)])) ?
                      (8'ha6) : ((reg184[(4'h9):(1'h1)] != ((8'ha4) ?
                          reg532 : reg205)) > $unsigned($signed(reg554))));
                  reg525 <= reg79;
                  if (reg543[(4'he):(3'h6)])
                    begin
                      reg526 <= reg542;
                      reg527 <= reg173[(1'h1):(1'h0)];
                      reg528 <= (~$signed((reg37[(1'h1):(1'h0)] - reg188[(2'h3):(1'h0)])));
                    end
                  else
                    begin
                      reg526 <= $unsigned((((8'ha0) != (~&forvar545)) ?
                          {(+(8'ha6))} : (^~$unsigned(reg545))));
                      reg527 <= (reg208 * ($unsigned($unsigned((8'ha5))) ?
                          (!reg51) : reg544));
                      reg528 <= {$unsigned($unsigned((wire7 ?
                              reg536 : reg514)))};
                      reg529 <= reg540;
                    end
                  for (forvar530 = (1'h0); (forvar530 < (2'h3)); forvar530 = (forvar530 + (1'h1)))
                    begin
                      reg531 <= $signed($signed(($signed(reg129) > (reg80 ?
                          (8'h9c) : reg132))));
                    end
                end
            end
        end
      if ((-forvar531[(4'hc):(1'h1)]))
        begin
          reg571 <= ($unsigned((^~$unsigned(reg60))) || reg529);
          for (forvar572 = (1'h0); (forvar572 < (1'h1)); forvar572 = (forvar572 + (1'h1)))
            begin
              if (({reg57} ?
                  ($unsigned((~|forvar508)) ?
                      reg107 : $unsigned((reg538 > reg500))) : $unsigned(({forvar494} ?
                      {reg509} : (reg182 ? reg44 : reg114)))))
                begin
                  for (forvar573 = (1'h0); (forvar573 < (2'h2)); forvar573 = (forvar573 + (1'h1)))
                    begin
                      reg574 <= {(!reg84)};
                      reg575 <= (^$unsigned(($signed((8'hb0)) ?
                          (~reg534) : {reg160})));
                      reg576 <= $signed({$unsigned((reg574 >>> reg571))});
                      reg577 <= {$unsigned(reg33[(1'h0):(1'h0)])};
                    end
                  for (forvar578 = (1'h0); (forvar578 < (1'h0)); forvar578 = (forvar578 + (1'h1)))
                    begin
                      reg579 <= reg543[(4'ha):(3'h4)];
                      reg580 <= {(((reg179 ? reg214 : (8'hb8)) ?
                                  reg503[(3'h4):(2'h2)] : {reg163}) ?
                              forvar549 : (~(+reg37)))};
                      reg581 <= ({reg511[(1'h1):(1'h1)]} ^ reg22);
                    end
                  reg582 <= reg218[(1'h0):(1'h0)];
                end
              else
                begin
                  if (reg571)
                    begin
                      reg573 <= $signed(($unsigned($signed(reg112)) ?
                          (((8'hb2) ?
                              reg497 : reg56) <<< $unsigned(reg18)) : $unsigned($signed((8'ha4)))));
                    end
                  else
                    begin
                      reg573 <= {$unsigned((~&reg504))};
                      reg574 <= (^reg156);
                    end
                  if (($signed(reg84[(4'h8):(3'h6)]) ?
                      reg148 : ($signed((8'ha5)) ?
                          $unsigned((8'hb6)) : (!$unsigned(reg139)))))
                    begin
                      reg575 <= $unsigned(($unsigned((reg127 ?
                              reg518 : reg177)) ?
                          $unsigned((!reg82)) : {(reg522 ? reg146 : reg154)}));
                    end
                  else
                    begin
                      reg575 <= (8'ha1);
                      reg576 <= ($signed(reg167[(2'h2):(1'h0)]) && reg174);
                      reg577 <= (({reg14[(2'h2):(1'h0)]} ?
                              reg200 : ($signed(reg203) < (forvar509 > reg168))) ?
                          ($signed($unsigned(reg59)) ?
                              ((reg130 & reg210) & (reg144 ?
                                  (8'h9c) : (8'hb2))) : $signed(reg13[(1'h1):(1'h0)])) : reg69[(3'h4):(1'h1)]);
                    end
                  if ((^~forvar520[(2'h2):(1'h0)]))
                    begin
                      reg578 <= $signed(reg508[(1'h0):(1'h0)]);
                      reg579 <= ($signed({reg151[(3'h6):(3'h5)]}) >>> (&(~(~^reg44))));
                      reg580 <= reg10;
                      reg581 <= (reg74[(1'h0):(1'h0)] != ($unsigned((-reg14)) ?
                          {(|reg558)} : (-reg553[(2'h3):(1'h0)])));
                    end
                  else
                    begin
                      reg578 <= $signed(reg82);
                      reg579 <= forvar495[(1'h1):(1'h0)];
                    end
                  for (forvar582 = (1'h0); (forvar582 < (2'h3)); forvar582 = (forvar582 + (1'h1)))
                    begin
                      reg583 <= $unsigned($signed((-$signed((8'h9e)))));
                      reg584 <= $unsigned(reg179[(4'hf):(3'h6)]);
                      reg585 <= $signed($signed((^reg508)));
                    end
                end
              for (forvar586 = (1'h0); (forvar586 < (2'h3)); forvar586 = (forvar586 + (1'h1)))
                begin
                  for (forvar587 = (1'h0); (forvar587 < (1'h1)); forvar587 = (forvar587 + (1'h1)))
                    begin
                      reg588 <= reg208[(1'h0):(1'h0)];
                      reg589 <= reg139[(2'h2):(2'h2)];
                      reg590 <= $unsigned($unsigned(((reg141 <= (8'hb4)) ?
                          reg588[(3'h4):(2'h3)] : (reg187 >>> reg16))));
                    end
                  if (reg584[(3'h4):(2'h3)])
                    begin
                      reg591 <= $signed({(reg219 >> {(8'ha1)})});
                      reg592 <= $signed($unsigned(reg142));
                      reg593 <= reg117;
                    end
                  else
                    begin
                      reg591 <= ($unsigned(reg183[(4'he):(1'h1)]) ?
                          {((8'hac) ?
                                  (reg156 ?
                                      reg204 : reg163) : $signed(reg593))} : reg519[(1'h1):(1'h0)]);
                      reg592 <= reg57;
                      reg593 <= ($signed($unsigned((reg539 ?
                          reg543 : reg188))) && {$unsigned((8'hb5))});
                      reg594 <= {((reg568 ?
                                  (reg70 - reg215) : reg192[(3'h6):(2'h3)]) ?
                              (reg152 ?
                                  (wire7 ?
                                      reg198 : reg205) : (reg526 <<< reg536)) : $unsigned(((8'ha1) ?
                                  reg106 : forvar578)))};
                    end
                  if (((+($signed(reg546) ?
                          (-reg103) : reg220[(4'h8):(2'h2)])) ?
                      $signed(reg130[(2'h3):(2'h2)]) : $unsigned(reg39[(3'h5):(2'h3)])))
                    begin
                      reg595 <= $unsigned((reg547 ?
                          reg198[(3'h6):(3'h5)] : $unsigned(reg121)));
                    end
                  else
                    begin
                      reg595 <= forvar501[(4'hc):(4'hb)];
                      reg596 <= $unsigned($unsigned(wire8[(1'h0):(1'h0)]));
                    end
                  reg597 <= reg169[(2'h3):(2'h2)];
                end
              for (forvar598 = (1'h0); (forvar598 < (1'h1)); forvar598 = (forvar598 + (1'h1)))
                begin
                  for (forvar599 = (1'h0); (forvar599 < (2'h2)); forvar599 = (forvar599 + (1'h1)))
                    begin
                      reg600 <= reg597[(4'h8):(1'h0)];
                    end
                  if ({$signed($unsigned((~|(8'hb1))))})
                    begin
                      reg601 <= reg576[(3'h6):(1'h1)];
                      reg602 <= $unsigned(((~|$unsigned(reg68)) ?
                          (8'h9d) : ($signed(forvar517) ?
                              (~^reg13) : $unsigned(reg27))));
                    end
                  else
                    begin
                      reg601 <= reg577;
                      reg602 <= (~|{$signed($signed(reg99))});
                      reg603 <= (reg110[(3'h4):(1'h1)] << ({reg97} ?
                          $signed((~&reg105)) : (&{(8'hb0)})));
                      reg604 <= reg100;
                    end
                  reg605 <= $unsigned($unsigned($unsigned({reg593})));
                end
            end
        end
      else
        begin
          for (forvar571 = (1'h0); (forvar571 < (1'h0)); forvar571 = (forvar571 + (1'h1)))
            begin
              for (forvar572 = (1'h0); (forvar572 < (2'h2)); forvar572 = (forvar572 + (1'h1)))
                begin
                  for (forvar573 = (1'h0); (forvar573 < (2'h3)); forvar573 = (forvar573 + (1'h1)))
                    begin
                      reg574 <= $signed(reg205);
                    end
                  if ($unsigned(reg591))
                    begin
                      reg575 <= $signed($unsigned(reg92[(1'h1):(1'h1)]));
                      reg576 <= (^$unsigned(((reg199 ?
                          reg163 : reg534) < (!reg194))));
                      reg577 <= $signed($unsigned(forvar573[(1'h0):(1'h0)]));
                      reg578 <= reg223;
                    end
                  else
                    begin
                      reg575 <= ((~^{$unsigned(reg534)}) ?
                          $signed($unsigned($unsigned(reg41))) : reg34[(1'h1):(1'h1)]);
                    end
                  if (($signed(({reg148} != (reg187 || reg495))) ?
                      reg536 : $unsigned(((^~(8'hb7)) ?
                          $unsigned(reg109) : (!reg526)))))
                    begin
                      reg579 <= ($unsigned($signed((reg177 ?
                          (8'hb8) : reg13))) ^ (~|reg517));
                      reg580 <= ((reg510 >> reg121) || $unsigned($unsigned($signed(reg560))));
                      reg581 <= (~|($unsigned($signed(reg13)) * (reg160 + reg105[(1'h0):(1'h0)])));
                      reg582 <= $signed(reg217);
                    end
                  else
                    begin
                      reg579 <= reg495[(3'h4):(1'h0)];
                      reg580 <= $signed($unsigned($signed({wire8})));
                    end
                  if (({((reg141 ? reg174 : reg517) ?
                          (~&reg18) : (forvar495 || reg44))} >>> ({$unsigned(reg183)} || reg569[(1'h0):(1'h0)])))
                    begin
                      reg583 <= (~^{((reg604 & reg26) - (^reg171))});
                    end
                  else
                    begin
                      reg583 <= ((^{reg535}) ?
                          (reg110[(3'h5):(1'h1)] ?
                              reg195 : ($signed(reg118) ?
                                  reg511 : forvar525)) : $signed($unsigned(reg604[(1'h1):(1'h1)])));
                      reg584 <= $unsigned((reg23 ?
                          {(reg503 ?
                                  reg187 : (8'hb0))} : forvar501[(4'ha):(2'h2)]));
                      reg585 <= $signed($signed($signed(reg36)));
                    end
                end
            end
          if ((({reg163} ?
              ((~|(8'had)) ~^ $signed(reg113)) : reg208) + $unsigned($signed((|reg185)))))
            begin
              reg586 <= reg183;
              for (forvar587 = (1'h0); (forvar587 < (2'h3)); forvar587 = (forvar587 + (1'h1)))
                begin
                  if ($signed(reg559[(1'h0):(1'h0)]))
                    begin
                      reg588 <= (reg539[(2'h3):(2'h2)] ?
                          reg10 : $unsigned($signed((reg597 <<< reg167))));
                      reg589 <= $unsigned($signed(((reg563 ? reg583 : reg205) ?
                          (~&(8'ha0)) : {reg193})));
                    end
                  else
                    begin
                      reg588 <= (-reg131[(4'h8):(3'h6)]);
                      reg589 <= (&reg514[(1'h0):(1'h0)]);
                    end
                  for (forvar590 = (1'h0); (forvar590 < (2'h3)); forvar590 = (forvar590 + (1'h1)))
                    begin
                      reg591 <= $signed((|$unsigned(reg43)));
                      reg592 <= ((8'hb1) + (~&reg30[(1'h1):(1'h1)]));
                      reg593 <= $signed(((^reg193) ?
                          (~|(reg557 >= reg513)) : ((~|reg188) ?
                              (wire7 ? reg33 : wire7) : reg145)));
                      reg594 <= {({reg592[(1'h1):(1'h0)]} ?
                              reg145 : (reg571 * {reg220}))};
                    end
                  reg595 <= {$unsigned(reg208)};
                  reg596 <= {$unsigned($signed(reg96[(1'h0):(1'h0)]))};
                end
              for (forvar597 = (1'h0); (forvar597 < (1'h1)); forvar597 = (forvar597 + (1'h1)))
                begin
                  for (forvar598 = (1'h0); (forvar598 < (1'h1)); forvar598 = (forvar598 + (1'h1)))
                    begin
                      reg599 <= reg543;
                      reg600 <= (-(&(((8'hb7) ? reg585 : (8'hb0)) ?
                          (reg220 ? reg160 : reg601) : (!reg171))));
                    end
                  for (forvar601 = (1'h0); (forvar601 < (1'h0)); forvar601 = (forvar601 + (1'h1)))
                    begin
                      reg602 <= $signed($unsigned(((forvar530 >= reg538) ?
                          (~|(8'hb6)) : $unsigned(reg36))));
                      reg603 <= (~&reg159[(4'h8):(4'h8)]);
                    end
                  for (forvar604 = (1'h0); (forvar604 < (2'h3)); forvar604 = (forvar604 + (1'h1)))
                    begin
                      reg605 <= reg66[(1'h0):(1'h0)];
                      reg606 <= $signed((8'ha8));
                    end
                end
              for (forvar607 = (1'h0); (forvar607 < (2'h3)); forvar607 = (forvar607 + (1'h1)))
                begin
                  if (reg117[(4'he):(3'h5)])
                    begin
                      reg608 <= (|((reg564 ?
                          (!reg162) : (&reg140)) >> $unsigned(reg174[(2'h3):(2'h3)])));
                      reg609 <= ((|($unsigned(reg546) << (~reg102))) + (~^reg99));
                      reg610 <= {{(8'hb9)}};
                    end
                  else
                    begin
                      reg608 <= reg170[(2'h2):(1'h0)];
                      reg609 <= (reg88[(4'hb):(4'ha)] < (reg130 ?
                          {(reg214 ?
                                  reg602 : reg179)} : forvar607[(2'h2):(1'h0)]));
                    end
                  for (forvar611 = (1'h0); (forvar611 < (1'h0)); forvar611 = (forvar611 + (1'h1)))
                    begin
                      reg612 <= reg110;
                      reg613 <= ((forvar526 ?
                          (~|(forvar517 == reg545)) : (reg214[(1'h1):(1'h0)] | (reg531 ?
                              reg21 : reg90))) * reg125[(3'h7):(3'h6)]);
                    end
                end
            end
          else
            begin
              if (((^$unsigned((reg166 ^~ (8'ha3)))) ?
                  ($signed($unsigned(reg185)) ?
                      $signed(reg585) : ((reg32 ?
                          (8'hba) : reg514) <<< (reg79 < reg30))) : $unsigned($signed(((8'hab) ?
                      reg149 : reg173)))))
                begin
                  reg586 <= reg566[(3'h5):(1'h0)];
                  for (forvar587 = (1'h0); (forvar587 < (1'h1)); forvar587 = (forvar587 + (1'h1)))
                    begin
                      reg588 <= (~^(|$unsigned((-(8'had)))));
                      reg589 <= reg555;
                      reg590 <= $unsigned($unsigned(((~&reg500) ?
                          (reg57 ? (8'ha2) : reg571) : (8'hb2))));
                    end
                  for (forvar591 = (1'h0); (forvar591 < (2'h3)); forvar591 = (forvar591 + (1'h1)))
                    begin
                      reg592 <= (|reg536);
                      reg593 <= reg78[(2'h3):(1'h1)];
                      reg594 <= (forvar520 ?
                          $signed((~|reg74[(1'h0):(1'h0)])) : {($signed((8'ha8)) ?
                                  (-reg160) : $unsigned(reg197))});
                    end
                  if ($unsigned((^~(+$unsigned(reg40)))))
                    begin
                      reg595 <= ((forvar545 != reg52[(2'h3):(1'h0)]) ^ ((~^{reg89}) > $unsigned({(8'h9f)})));
                    end
                  else
                    begin
                      reg595 <= ((reg118 ? $signed((+forvar599)) : reg13) ?
                          reg128 : $signed({forvar582}));
                      reg596 <= (~&((^~reg519[(1'h1):(1'h1)]) ?
                          reg586 : reg164));
                      reg597 <= reg109;
                      reg598 <= $signed(($signed($unsigned((8'hb1))) ?
                          (reg73[(1'h0):(1'h0)] ?
                              $unsigned(reg213) : forvar496[(4'hc):(3'h4)]) : $signed($signed(reg23))));
                    end
                end
              else
                begin
                  if (reg195)
                    begin
                      reg586 <= $unsigned($unsigned(((+reg165) <<< reg78[(3'h5):(3'h5)])));
                      reg587 <= (8'hba);
                      reg588 <= forvar611;
                    end
                  else
                    begin
                      reg586 <= (~^$unsigned(((+(8'hae)) < $unsigned(reg194))));
                      reg587 <= $signed((reg148 << (((8'hb4) & reg499) ^~ (|reg19))));
                      reg588 <= reg605;
                      reg589 <= reg40[(3'h6):(1'h0)];
                    end
                  for (forvar590 = (1'h0); (forvar590 < (1'h1)); forvar590 = (forvar590 + (1'h1)))
                    begin
                      reg591 <= (^$unsigned({(wire7 - reg141)}));
                      reg592 <= {(($signed(reg130) ?
                              (reg166 < reg167) : {reg30}) || reg563[(1'h0):(1'h0)])};
                      reg593 <= (+reg65);
                      reg594 <= $unsigned(forvar591);
                    end
                end
            end
          if (reg186)
            begin
              for (forvar614 = (1'h0); (forvar614 < (2'h3)); forvar614 = (forvar614 + (1'h1)))
                begin
                  if (($unsigned($unsigned((^reg503))) ?
                      (~((reg37 ? reg515 : (8'h9d)) ?
                          $unsigned(reg211) : reg527[(3'h7):(3'h5)])) : $unsigned(forvar520[(2'h2):(1'h0)])))
                    begin
                      reg615 <= forvar614;
                      reg616 <= (~&reg111);
                      reg617 <= $signed($unsigned(reg200));
                      reg618 <= {((8'hb7) << $signed((&reg598)))};
                    end
                  else
                    begin
                      reg615 <= $signed({($signed(reg176) | (forvar530 ?
                              reg52 : reg564))});
                      reg616 <= ($unsigned($signed(reg125[(2'h2):(1'h1)])) ?
                          reg43[(4'h9):(1'h0)] : $unsigned($unsigned(((8'ha0) ?
                              reg191 : reg150))));
                    end
                end
              for (forvar619 = (1'h0); (forvar619 < (2'h3)); forvar619 = (forvar619 + (1'h1)))
                begin
                  for (forvar620 = (1'h0); (forvar620 < (2'h2)); forvar620 = (forvar620 + (1'h1)))
                    begin
                      reg621 <= (($signed(reg16[(2'h3):(1'h0)]) <= (reg18[(3'h7):(3'h4)] ^ {reg557})) >>> reg47[(2'h3):(1'h0)]);
                      reg622 <= {{forvar511[(2'h2):(1'h1)]}};
                      reg623 <= ((reg59 <= reg112[(2'h3):(1'h0)]) || ($signed((reg39 * (8'ha4))) ?
                          ({(8'hb4)} ?
                              reg553[(1'h0):(1'h0)] : (reg192 ~^ (8'h9c))) : ((+reg537) ?
                              reg96 : reg505[(1'h0):(1'h0)])));
                      reg624 <= $signed($signed({(~reg586)}));
                    end
                end
              if (reg172)
                begin
                  for (forvar625 = (1'h0); (forvar625 < (2'h2)); forvar625 = (forvar625 + (1'h1)))
                    begin
                      reg626 <= ((!{$signed((8'hac))}) <= ($unsigned(((8'hb8) <<< forvar614)) ?
                          $unsigned($unsigned(reg623)) : $signed(forvar625[(3'h4):(2'h2)])));
                      reg627 <= $signed($signed((^(-(8'hac)))));
                      reg628 <= $unsigned($signed($unsigned((reg506 ?
                          forvar590 : reg126))));
                    end
                  if ((~^forvar590[(2'h2):(1'h1)]))
                    begin
                      reg629 <= ({reg580} >> reg210[(4'ha):(3'h6)]);
                      reg630 <= reg515[(3'h4):(3'h4)];
                      reg631 <= (reg69[(3'h7):(1'h1)] != $signed((reg113 ?
                          (!reg114) : (reg23 ? (8'hac) : reg508))));
                    end
                  else
                    begin
                      reg629 <= $unsigned((8'hb2));
                    end
                  for (forvar632 = (1'h0); (forvar632 < (2'h3)); forvar632 = (forvar632 + (1'h1)))
                    begin
                      reg633 <= $signed((8'ha6));
                    end
                  reg634 <= $signed((((reg96 ? reg160 : reg225) ?
                          (reg69 >> reg530) : reg608[(3'h6):(1'h1)]) ?
                      (~|reg38[(2'h3):(1'h1)]) : $signed(((8'ha9) >>> reg216))));
                end
              else
                begin
                  for (forvar625 = (1'h0); (forvar625 < (1'h1)); forvar625 = (forvar625 + (1'h1)))
                    begin
                      reg626 <= ($signed((~|$unsigned(reg199))) & reg77);
                      reg627 <= {reg525[(3'h5):(2'h2)]};
                    end
                  if ((reg531[(4'h9):(3'h5)] ? reg531 : reg200[(3'h6):(2'h2)]))
                    begin
                      reg628 <= $signed((forvar542[(4'hc):(3'h5)] ^~ $unsigned((~|reg542))));
                      reg629 <= (reg520[(3'h6):(3'h5)] ?
                          reg618[(2'h3):(2'h2)] : reg575[(3'h7):(3'h4)]);
                    end
                  else
                    begin
                      reg628 <= reg59[(2'h2):(2'h2)];
                      reg629 <= ($signed($unsigned($unsigned(reg525))) ?
                          $signed((!((8'ha2) ?
                              reg502 : reg594))) : ($signed(reg552) ^ ($signed(reg518) || (reg563 | reg56))));
                      reg630 <= $unsigned((!{(forvar572 ? reg48 : forvar598)}));
                      reg631 <= $signed((reg51 <<< (((8'h9e) - reg516) > $signed(forvar499))));
                    end
                  for (forvar632 = (1'h0); (forvar632 < (2'h3)); forvar632 = (forvar632 + (1'h1)))
                    begin
                      reg633 <= (+{forvar620});
                    end
                  reg634 <= $signed($signed($signed((^~reg583))));
                end
            end
          else
            begin
              reg614 <= reg37;
            end
          if ($unsigned(({((8'ha4) ? reg88 : reg626)} ?
              forvar545 : ((reg22 ? reg552 : reg55) ^~ reg627))))
            begin
              reg635 <= reg200;
              for (forvar636 = (1'h0); (forvar636 < (1'h0)); forvar636 = (forvar636 + (1'h1)))
                begin
                  if ({(~&$signed((&reg499)))})
                    begin
                      reg637 <= (reg96[(4'hc):(4'h9)] ?
                          reg594[(1'h0):(1'h0)] : reg84);
                      reg638 <= ($signed({{(8'haa)}}) >= $unsigned($signed((reg614 + reg584))));
                      reg639 <= $unsigned(((~^$signed((8'hb5))) * $unsigned((^reg638))));
                    end
                  else
                    begin
                      reg637 <= $unsigned(({{forvar625}} ?
                          ($signed(reg570) ?
                              {(8'hb4)} : (reg175 & (8'hb1))) : $signed($signed(forvar501))));
                    end
                  for (forvar640 = (1'h0); (forvar640 < (1'h0)); forvar640 = (forvar640 + (1'h1)))
                    begin
                      reg641 <= $signed({{reg92}});
                      reg642 <= (reg589[(4'ha):(3'h6)] ?
                          ((+forvar620[(3'h6):(1'h1)]) > (reg206 ?
                              reg104[(4'ha):(4'ha)] : reg538[(5'h10):(4'ha)])) : ($unsigned((reg101 ?
                                  reg172 : reg174)) ?
                              {{reg522}} : (~|reg205[(4'h8):(3'h7)])));
                      reg643 <= ($unsigned(reg571) ?
                          (~^{$signed(reg165)}) : reg148);
                    end
                  if ((reg145 ? reg129[(3'h5):(1'h0)] : reg566))
                    begin
                      reg644 <= $unsigned(reg107);
                      reg645 <= (^~$signed({reg41}));
                      reg646 <= {$unsigned(reg213)};
                    end
                  else
                    begin
                      reg644 <= (((~(~&forvar619)) ?
                              $unsigned((^reg27)) : reg553) ?
                          $unsigned($signed(reg115)) : (($signed(reg623) <<< $unsigned(forvar601)) ?
                              {reg124[(2'h2):(2'h2)]} : reg513));
                      reg645 <= reg148;
                      reg646 <= (|(($signed(reg642) ^ (&reg581)) ~^ $signed(reg525[(2'h3):(1'h0)])));
                    end
                end
              if ((~|{(reg74 ? (|reg43) : $signed(reg586))}))
                begin
                  if ($signed((reg176 * reg196[(1'h1):(1'h1)])))
                    begin
                      reg647 <= (^reg182[(2'h3):(1'h0)]);
                      reg648 <= (|$signed((~(reg214 ? (8'hb1) : reg540))));
                      reg649 <= reg545;
                      reg650 <= ((reg617 ?
                              $unsigned(reg570[(4'he):(3'h7)]) : $unsigned((reg604 - reg36))) ?
                          {(8'ha6)} : $unsigned(reg100[(2'h3):(2'h3)]));
                    end
                  else
                    begin
                      reg647 <= reg583;
                      reg648 <= reg179[(5'h10):(4'hd)];
                      reg649 <= (^($unsigned({(8'h9e)}) ?
                          {$unsigned(reg132)} : reg200));
                    end
                  for (forvar651 = (1'h0); (forvar651 < (2'h3)); forvar651 = (forvar651 + (1'h1)))
                    begin
                      reg652 <= (^reg189);
                    end
                  reg653 <= (-$signed(((reg588 ? (8'h9e) : reg66) ?
                      (reg556 > reg59) : (reg33 && reg168))));
                  reg654 <= $signed($signed($signed(reg210[(3'h5):(2'h3)])));
                end
              else
                begin
                  if ({reg142[(2'h3):(2'h2)]})
                    begin
                      reg647 <= (((^$unsigned(forvar517)) ?
                          (~^(8'haf)) : $unsigned((reg521 ?
                              reg626 : reg208))) > forvar573[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg647 <= reg652[(4'h9):(1'h1)];
                      reg648 <= (8'ha5);
                      reg649 <= forvar497;
                      reg650 <= (((^$signed(reg518)) ?
                          reg577[(1'h0):(1'h0)] : reg571[(4'h9):(2'h2)]) * reg147[(1'h1):(1'h1)]);
                    end
                  for (forvar651 = (1'h0); (forvar651 < (1'h1)); forvar651 = (forvar651 + (1'h1)))
                    begin
                      reg652 <= reg516[(3'h5):(2'h3)];
                    end
                  reg653 <= {$unsigned(reg631)};
                end
            end
          else
            begin
              for (forvar635 = (1'h0); (forvar635 < (2'h3)); forvar635 = (forvar635 + (1'h1)))
                begin
                  if (((reg56[(4'hc):(3'h5)] ?
                          ((reg22 << reg191) >>> {reg140}) : ($unsigned(reg545) ?
                              (reg219 ? reg546 : (8'hb7)) : reg90)) ?
                      (|reg514) : $unsigned(((reg122 ~^ forvar512) ?
                          (forvar499 ? forvar586 : reg635) : {reg34}))))
                    begin
                      reg636 <= (forvar545 >> $signed((reg545 || $signed(reg113))));
                      reg637 <= reg101;
                    end
                  else
                    begin
                      reg636 <= reg638;
                      reg637 <= $unsigned(reg197[(3'h5):(1'h0)]);
                      reg638 <= $signed($unsigned($signed($unsigned(reg115))));
                    end
                end
              for (forvar639 = (1'h0); (forvar639 < (1'h1)); forvar639 = (forvar639 + (1'h1)))
                begin
                  for (forvar640 = (1'h0); (forvar640 < (2'h3)); forvar640 = (forvar640 + (1'h1)))
                    begin
                      reg641 <= ((forvar500[(1'h0):(1'h0)] ?
                              ((8'hb0) ?
                                  $unsigned(reg149) : reg650) : (~&$signed((8'hb1)))) ?
                          (8'hb6) : ((~^$signed((8'ha2))) & $signed((reg124 == reg117))));
                      reg642 <= (8'h9d);
                    end
                  if ((|$signed($unsigned({(8'ha8)}))))
                    begin
                      reg643 <= (&reg40[(2'h2):(1'h0)]);
                      reg644 <= reg542;
                      reg645 <= (8'ha4);
                      reg646 <= {($unsigned(reg517) ?
                              reg105 : reg134[(3'h7):(2'h2)])};
                    end
                  else
                    begin
                      reg643 <= ((reg216 & {(reg201 || forvar545)}) ^~ $signed($signed({forvar586})));
                      reg644 <= reg539[(1'h1):(1'h1)];
                      reg645 <= (!$unsigned((reg529[(4'hb):(2'h2)] <<< {reg645})));
                    end
                  for (forvar647 = (1'h0); (forvar647 < (2'h2)); forvar647 = (forvar647 + (1'h1)))
                    begin
                      reg648 <= ($unsigned($unsigned((&reg631))) - (~^{reg56}));
                      reg649 <= reg544;
                      reg650 <= reg73;
                      reg651 <= reg502;
                    end
                  for (forvar652 = (1'h0); (forvar652 < (2'h3)); forvar652 = (forvar652 + (1'h1)))
                    begin
                      reg653 <= (^~reg93);
                      reg654 <= {(({reg111} + reg595[(1'h0):(1'h0)]) <= (8'h9d))};
                    end
                end
            end
        end
      if (reg21)
        begin
          if ($unsigned(((forvar571 <= {reg186}) << (reg553[(2'h3):(2'h3)] + {(8'hb8)}))))
            begin
              if ((~reg605))
                begin
                  for (forvar655 = (1'h0); (forvar655 < (2'h3)); forvar655 = (forvar655 + (1'h1)))
                    begin
                      reg656 <= (8'ha2);
                      reg657 <= (|{(~^reg125[(2'h2):(1'h1)])});
                      reg658 <= (~|reg167[(3'h4):(2'h3)]);
                    end
                  reg659 <= reg534[(3'h5):(3'h5)];
                  for (forvar660 = (1'h0); (forvar660 < (2'h3)); forvar660 = (forvar660 + (1'h1)))
                    begin
                      reg661 <= (reg524[(2'h3):(2'h3)] ?
                          (reg145 ?
                              $signed(reg37) : $unsigned((forvar655 >>> reg57))) : ($signed($unsigned(forvar531)) ?
                              reg145[(1'h0):(1'h0)] : reg554[(3'h7):(3'h5)]));
                      reg662 <= (^~(~|$signed((reg124 + reg573))));
                      reg663 <= ((reg518[(4'hc):(4'hb)] == (|(forvar655 > (8'ha6)))) == (^reg628));
                      reg664 <= $unsigned((~^(-$signed(reg564))));
                    end
                end
              else
                begin
                  if ((8'hba))
                    begin
                      reg655 <= $signed($signed($signed($unsigned(forvar636))));
                      reg656 <= (reg643[(1'h0):(1'h0)] ?
                          (|(forvar499 < {reg556})) : ((8'ha8) ?
                              ({reg182} ^ forvar520[(1'h0):(1'h0)]) : $unsigned(reg30)));
                      reg657 <= (~(&$unsigned((~^reg518))));
                    end
                  else
                    begin
                      reg655 <= $signed(($signed($unsigned((8'ha3))) >> {reg545[(4'hb):(1'h0)]}));
                      reg656 <= reg529[(1'h0):(1'h0)];
                      reg657 <= (^~({reg574[(4'he):(2'h3)]} <= ((forvar549 << forvar525) ?
                          reg582 : $signed(reg220))));
                    end
                  if ($unsigned(((+forvar655) ?
                      {$unsigned((8'hb9))} : reg593[(3'h5):(2'h3)])))
                    begin
                      reg658 <= (~(~&(|(~reg182))));
                      reg659 <= $unsigned($signed(reg92));
                      reg660 <= ($unsigned($signed($signed((8'hb1)))) ?
                          forvar590 : $signed($unsigned($signed(reg556))));
                      reg661 <= reg655[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg658 <= {($unsigned((-reg64)) ?
                              (reg27 ?
                                  $signed(reg579) : $signed((8'hac))) : (~&$signed(reg167)))};
                      reg659 <= reg547[(1'h1):(1'h0)];
                      reg660 <= ((($unsigned((8'hb2)) ?
                          (8'ha7) : (reg630 ?
                              reg103 : reg144)) != ($unsigned((8'ha1)) || $signed(reg628))) ^ (($signed(reg205) - $unsigned(forvar510)) ?
                          reg151[(1'h1):(1'h0)] : (~&reg660)));
                      reg661 <= $unsigned(($unsigned($signed((8'hb0))) <= (8'hb1)));
                    end
                  if (reg217)
                    begin
                      reg662 <= $unsigned((~|reg570));
                    end
                  else
                    begin
                      reg662 <= ((8'h9c) ?
                          (reg622 ?
                              (^~(reg13 ?
                                  (8'ha6) : reg206)) : $signed($signed((8'ha4)))) : reg555[(3'h4):(1'h0)]);
                      reg663 <= forvar573;
                      reg664 <= $signed({forvar652});
                    end
                end
            end
          else
            begin
              for (forvar655 = (1'h0); (forvar655 < (1'h1)); forvar655 = (forvar655 + (1'h1)))
                begin
                  if ({(~(reg616[(4'ha):(1'h1)] ?
                          (~^reg150) : (reg501 ? reg504 : reg33)))})
                    begin
                      reg656 <= reg45[(4'hb):(4'ha)];
                      reg657 <= ($signed(((reg116 ? reg518 : reg591) ?
                          $signed(reg189) : (reg175 || (8'h9f)))) >= $unsigned((-$signed(forvar598))));
                      reg658 <= reg548[(3'h6):(3'h6)];
                      reg659 <= $unsigned(reg502);
                    end
                  else
                    begin
                      reg656 <= forvar525[(1'h1):(1'h1)];
                      reg657 <= ({forvar549[(2'h2):(2'h2)]} ^~ (reg41 ?
                          $signed((reg195 ?
                              reg554 : reg103)) : ({reg168} ~^ {(8'had)})));
                      reg658 <= $signed((((-reg545) ?
                              {reg130} : $signed((8'hb5))) ?
                          (8'hae) : ($unsigned(reg612) ?
                              $signed(reg516) : ((8'haa) ?
                                  forvar651 : reg506))));
                      reg659 <= reg548;
                    end
                  for (forvar660 = (1'h0); (forvar660 < (2'h2)); forvar660 = (forvar660 + (1'h1)))
                    begin
                      reg661 <= ({(~^$signed(reg88))} ?
                          ((-(8'hb3)) != (~^reg584)) : $signed((^(+reg215))));
                      reg662 <= reg120;
                    end
                  reg663 <= reg149;
                  if ($signed((~|reg591[(1'h1):(1'h1)])))
                    begin
                      reg664 <= $signed(($unsigned((8'hb6)) >> forvar511[(4'h8):(3'h6)]));
                      reg665 <= ((!{(reg510 ~^ reg162)}) + {{(reg635 & (8'ha2))}});
                      reg666 <= ((($unsigned((8'ha4)) ?
                              (reg564 & reg205) : $signed(reg21)) <<< $signed($signed(forvar519))) ?
                          {(forvar619 + $signed(reg152))} : forvar510[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg664 <= $signed({((forvar587 >> reg221) ?
                              ((8'hac) ? reg579 : reg623) : (^reg184))});
                      reg665 <= forvar512;
                      reg666 <= ((~&$unsigned((reg552 ?
                          reg575 : reg79))) ~^ ((((8'hb4) && reg642) ~^ $signed(reg496)) == (~^$unsigned(reg110))));
                      reg667 <= reg41;
                    end
                end
            end
          if (forvar604)
            begin
              if ({reg634})
                begin
                  for (forvar668 = (1'h0); (forvar668 < (1'h0)); forvar668 = (forvar668 + (1'h1)))
                    begin
                      reg669 <= {reg495};
                      reg670 <= (reg77[(1'h0):(1'h0)] >>> {reg507[(3'h5):(1'h0)]});
                      reg671 <= forvar571[(2'h2):(1'h1)];
                      reg672 <= reg551;
                    end
                end
              else
                begin
                  reg668 <= (reg555[(2'h2):(2'h2)] >>> reg633[(4'h9):(3'h7)]);
                  for (forvar669 = (1'h0); (forvar669 < (1'h1)); forvar669 = (forvar669 + (1'h1)))
                    begin
                      reg670 <= reg197[(2'h3):(1'h1)];
                      reg671 <= (^~$unsigned(reg174));
                    end
                  if (($signed($signed((-reg629))) ^~ reg47[(1'h1):(1'h1)]))
                    begin
                      reg672 <= forvar625;
                    end
                  else
                    begin
                      reg672 <= (reg522 & (8'hb0));
                      reg673 <= reg531[(2'h3):(1'h0)];
                      reg674 <= $unsigned(reg211);
                      reg675 <= reg647;
                    end
                  for (forvar676 = (1'h0); (forvar676 < (2'h3)); forvar676 = (forvar676 + (1'h1)))
                    begin
                      reg677 <= (reg194 ?
                          {($unsigned(reg498) + reg569)} : reg127);
                      reg678 <= reg139[(3'h6):(3'h6)];
                      reg679 <= (^$unsigned($signed((^reg102))));
                      reg680 <= $unsigned(reg585);
                    end
                end
              reg681 <= forvar655;
            end
          else
            begin
              if ($signed($signed(reg96)))
                begin
                  for (forvar668 = (1'h0); (forvar668 < (1'h1)); forvar668 = (forvar668 + (1'h1)))
                    begin
                      reg669 <= $unsigned(reg518);
                      reg670 <= (~&$signed(((reg519 ?
                          (8'h9e) : forvar519) <<< reg622)));
                      reg671 <= ($unsigned($unsigned($signed(reg101))) ?
                          (^reg134[(2'h3):(1'h0)]) : $unsigned(reg110[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar668 = (1'h0); (forvar668 < (2'h3)); forvar668 = (forvar668 + (1'h1)))
                    begin
                      reg669 <= (reg630 - ((|(reg635 && reg96)) != {reg616[(4'h9):(2'h2)]}));
                      reg670 <= reg521;
                      reg671 <= reg571[(4'hc):(4'h9)];
                    end
                  if ((~|forvar639[(3'h7):(3'h5)]))
                    begin
                      reg672 <= ($unsigned((&reg168)) ?
                          (~$signed(reg171[(3'h5):(1'h1)])) : $signed((|$unsigned(reg175))));
                    end
                  else
                    begin
                      reg672 <= {$signed((~&(reg669 ? reg19 : reg50)))};
                    end
                  reg673 <= reg667;
                end
              if (reg577[(1'h0):(1'h0)])
                begin
                  reg674 <= (8'hac);
                end
              else
                begin
                  if ((8'hb9))
                    begin
                      reg674 <= (reg673[(4'hb):(4'h9)] ?
                          (8'haf) : ((|(~|forvar586)) ?
                              {{reg115}} : (|{reg156})));
                      reg675 <= reg92;
                    end
                  else
                    begin
                      reg674 <= reg93[(4'h9):(3'h4)];
                    end
                  for (forvar676 = (1'h0); (forvar676 < (2'h2)); forvar676 = (forvar676 + (1'h1)))
                    begin
                      reg677 <= reg210[(3'h6):(3'h6)];
                    end
                  for (forvar678 = (1'h0); (forvar678 < (2'h2)); forvar678 = (forvar678 + (1'h1)))
                    begin
                      reg679 <= $signed((~|reg64[(1'h0):(1'h0)]));
                      reg680 <= $unsigned($unsigned($unsigned((reg636 ?
                          reg187 : reg612))));
                    end
                  if ({(^~$unsigned(forvar524))})
                    begin
                      reg681 <= reg626[(3'h5):(3'h5)];
                      reg682 <= forvar578;
                      reg683 <= ({reg624} != (+reg122));
                    end
                  else
                    begin
                      reg681 <= reg170;
                      reg682 <= ($signed(reg114) ?
                          reg496 : $signed(((^~(8'hb2)) >= $unsigned(reg210))));
                      reg683 <= reg128;
                    end
                end
            end
          if (({(8'had)} && {$unsigned(reg118[(2'h2):(1'h1)])}))
            begin
              reg684 <= ($unsigned((~^$unsigned(reg514))) != $signed($signed($unsigned(reg55))));
              for (forvar685 = (1'h0); (forvar685 < (2'h2)); forvar685 = (forvar685 + (1'h1)))
                begin
                  reg686 <= reg626[(2'h3):(1'h1)];
                  reg687 <= (reg599 ^ $signed((^~{reg79})));
                  if ($signed({reg27}))
                    begin
                      reg688 <= ($unsigned($unsigned(reg108[(2'h3):(1'h0)])) & (((8'h9f) + (~|(8'hba))) ?
                          ($unsigned((8'hb7)) ?
                              reg197[(3'h7):(3'h7)] : ((8'ha9) ^~ reg634)) : reg643[(3'h4):(2'h3)]));
                    end
                  else
                    begin
                      reg688 <= $unsigned($signed($unsigned((+wire8))));
                      reg689 <= reg109;
                    end
                  if ({(-reg657)})
                    begin
                      reg690 <= ({$signed((~reg206))} ?
                          (reg580 ?
                              reg129 : reg567[(1'h1):(1'h1)]) : $unsigned($unsigned((reg197 ?
                              forvar651 : forvar676))));
                      reg691 <= $unsigned({forvar505[(2'h3):(1'h0)]});
                    end
                  else
                    begin
                      reg690 <= (reg643[(2'h3):(1'h1)] ^~ $signed($signed($signed(reg577))));
                      reg691 <= (($signed((8'hac)) > (reg73 ?
                              reg626[(3'h4):(3'h4)] : reg189[(1'h1):(1'h0)])) ?
                          (8'hb8) : $unsigned(($unsigned(reg656) ?
                              reg40 : reg37[(3'h4):(1'h0)])));
                      reg692 <= reg585[(2'h2):(1'h1)];
                    end
                end
              if ({(~{reg526})})
                begin
                  if ((reg115 <= (^reg117[(5'h10):(4'hf)])))
                    begin
                      reg693 <= ({reg204} ?
                          ((+reg155[(4'hd):(4'hc)]) ?
                              {$signed((8'hb7))} : forvar651[(3'h4):(3'h4)]) : ((-(reg170 ?
                              reg667 : reg668)) >>> ((forvar496 ?
                                  reg199 : reg37) ?
                              reg506[(3'h4):(3'h4)] : reg102[(3'h7):(2'h2)])));
                      reg694 <= forvar495;
                      reg695 <= reg16[(4'h9):(4'h9)];
                      reg696 <= ($unsigned($signed((reg505 | reg154))) ?
                          ((reg48[(1'h0):(1'h0)] != (8'hb1)) | reg124) : (&$signed($signed(wire7))));
                    end
                  else
                    begin
                      reg693 <= (wire7 ?
                          reg531[(4'h9):(3'h6)] : (reg651[(2'h3):(1'h1)] ?
                              reg679[(2'h2):(1'h0)] : reg116[(2'h3):(1'h0)]));
                      reg694 <= ($signed(($unsigned((8'had)) ?
                          $unsigned(reg667) : $signed(reg687))) ~^ ((reg499[(3'h6):(1'h0)] ?
                          forvar517 : (&(8'ha8))) | $signed($signed(reg45))));
                      reg695 <= reg672[(3'h6):(1'h0)];
                      reg696 <= wire6;
                    end
                end
              else
                begin
                  if (reg151[(1'h0):(1'h0)])
                    begin
                      reg693 <= (~(reg536 ?
                          $signed($signed(reg142)) : reg547[(1'h1):(1'h1)]));
                      reg694 <= reg573;
                    end
                  else
                    begin
                      reg693 <= reg60[(3'h4):(1'h1)];
                      reg694 <= $unsigned(reg70);
                      reg695 <= (&($unsigned($signed(reg69)) << (reg145[(2'h2):(2'h2)] ?
                          (reg154 ? reg41 : reg128) : $unsigned(reg674))));
                    end
                end
              for (forvar697 = (1'h0); (forvar697 < (1'h1)); forvar697 = (forvar697 + (1'h1)))
                begin
                  for (forvar698 = (1'h0); (forvar698 < (2'h2)); forvar698 = (forvar698 + (1'h1)))
                    begin
                      reg699 <= (((|(-reg581)) ~^ $signed((8'ha0))) | (|((reg635 ?
                              reg498 : reg659) ?
                          (8'h9f) : $unsigned(reg692))));
                      reg700 <= {reg684[(4'h9):(3'h6)]};
                    end
                  for (forvar701 = (1'h0); (forvar701 < (1'h1)); forvar701 = (forvar701 + (1'h1)))
                    begin
                      reg702 <= (reg176 <= (forvar510 ?
                          ((reg42 ? reg117 : forvar611) != ((8'h9d) ?
                              (8'hb8) : reg594)) : (&$unsigned((8'hb3)))));
                    end
                end
            end
          else
            begin
              if ((|(forvar611 ?
                  $unsigned(reg111) : (reg39[(3'h4):(2'h3)] ^~ {reg678}))))
                begin
                  for (forvar684 = (1'h0); (forvar684 < (1'h0)); forvar684 = (forvar684 + (1'h1)))
                    begin
                      reg685 <= ($signed((~forvar511[(3'h6):(3'h6)])) << $unsigned((^$signed(reg517))));
                      reg686 <= (({(reg21 ? forvar550 : (8'ha8))} ?
                              (^~$unsigned((8'hab))) : $unsigned(reg527)) ?
                          reg127[(2'h2):(1'h0)] : (~|$unsigned((forvar508 ?
                              reg524 : reg10))));
                      reg687 <= ((((&reg38) ? forvar520 : (reg650 ~^ reg530)) ?
                          $unsigned(reg188) : $unsigned($unsigned(forvar639))) > (!((wire492 ^~ forvar590) ?
                          reg33[(3'h5):(2'h3)] : $unsigned(forvar524))));
                    end
                  if (((((reg135 && (8'hac)) ?
                          (reg74 + reg68) : (reg219 ? forvar611 : reg111)) ?
                      $unsigned(forvar505[(2'h3):(1'h1)]) : ($unsigned(forvar619) ?
                          (!reg596) : $unsigned((8'ha9)))) <= ((|$signed(reg90)) > reg57)))
                    begin
                      reg688 <= (^reg175[(4'hf):(3'h4)]);
                      reg689 <= {reg523};
                    end
                  else
                    begin
                      reg688 <= (~^$signed($signed(reg119)));
                      reg689 <= ($unsigned($signed($unsigned((8'hac)))) < (+{reg615[(2'h3):(1'h0)]}));
                      reg690 <= $signed(($unsigned(reg565) - (-(forvar514 | reg680))));
                      reg691 <= forvar591;
                    end
                end
              else
                begin
                  if ((-((reg167 - reg670[(3'h7):(1'h1)]) ?
                      reg596 : reg123[(2'h3):(1'h1)])))
                    begin
                      reg684 <= forvar495[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg684 <= (((^$signed(reg88)) ?
                          {forvar678[(1'h0):(1'h0)]} : reg672[(4'h9):(1'h0)]) < (reg559[(2'h2):(1'h0)] <= {(8'ha1)}));
                    end
                  reg685 <= reg495;
                end
              for (forvar692 = (1'h0); (forvar692 < (1'h0)); forvar692 = (forvar692 + (1'h1)))
                begin
                  if (((~|reg142[(1'h1):(1'h0)]) >= $unsigned(forvar508[(1'h1):(1'h1)])))
                    begin
                      reg693 <= forvar660[(3'h5):(2'h3)];
                      reg694 <= $signed((({reg110} + (|reg512)) ?
                          reg647 : $unsigned($unsigned(forvar601))));
                      reg695 <= reg695;
                    end
                  else
                    begin
                      reg693 <= $signed((|(reg16 & (forvar497 & reg43))));
                    end
                  for (forvar696 = (1'h0); (forvar696 < (2'h3)); forvar696 = (forvar696 + (1'h1)))
                    begin
                      reg697 <= $unsigned({reg209[(3'h5):(2'h2)]});
                      reg698 <= (-($signed((&reg540)) || ($unsigned(reg674) ?
                          (|reg582) : (!reg508))));
                      reg699 <= {(~&$signed($signed(reg193)))};
                    end
                end
              for (forvar700 = (1'h0); (forvar700 < (1'h0)); forvar700 = (forvar700 + (1'h1)))
                begin
                  if ({$unsigned(((~|(8'hb1)) ^~ (reg592 <= (8'hae))))})
                    begin
                      reg701 <= $unsigned(reg667);
                      reg702 <= reg577[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg701 <= (($unsigned((reg148 == forvar655)) >= reg578[(2'h3):(1'h1)]) != ({$unsigned(reg665)} >> (^~(|reg81))));
                    end
                  for (forvar703 = (1'h0); (forvar703 < (2'h3)); forvar703 = (forvar703 + (1'h1)))
                    begin
                      reg704 <= {reg69[(2'h3):(2'h3)]};
                      reg705 <= $signed(reg78);
                      reg706 <= {reg143};
                    end
                end
            end
        end
      else
        begin
          for (forvar655 = (1'h0); (forvar655 < (2'h2)); forvar655 = (forvar655 + (1'h1)))
            begin
              if (reg150)
                begin
                  if (reg183[(3'h4):(2'h2)])
                    begin
                      reg656 <= $unsigned($signed($unsigned((reg677 ?
                          (8'haa) : forvar497))));
                      reg657 <= $signed($unsigned((&reg212[(4'hb):(4'ha)])));
                      reg658 <= reg635[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg656 <= reg661[(1'h1):(1'h1)];
                      reg657 <= {(8'haa)};
                      reg658 <= reg184[(4'hc):(4'h9)];
                      reg659 <= (forvar520[(1'h1):(1'h0)] ?
                          (8'ha1) : forvar697[(4'ha):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar656 = (1'h0); (forvar656 < (1'h1)); forvar656 = (forvar656 + (1'h1)))
                    begin
                      reg657 <= (reg59[(3'h5):(1'h0)] == $signed((+(reg93 >= reg191))));
                    end
                  for (forvar658 = (1'h0); (forvar658 < (1'h1)); forvar658 = (forvar658 + (1'h1)))
                    begin
                      reg659 <= (+(((&reg704) | reg146[(4'h9):(2'h3)]) < (~&$unsigned((8'hae)))));
                      reg660 <= $unsigned(($unsigned($unsigned(reg70)) > ((~reg664) ?
                          (reg223 ? reg65 : (8'ha7)) : (reg209 ?
                              reg222 : reg528))));
                    end
                  for (forvar661 = (1'h0); (forvar661 < (1'h1)); forvar661 = (forvar661 + (1'h1)))
                    begin
                      reg662 <= (8'h9f);
                      reg663 <= reg10;
                    end
                  if (forvar525)
                    begin
                      reg664 <= reg566[(3'h7):(2'h2)];
                      reg665 <= reg132;
                      reg666 <= $unsigned((-((reg512 ?
                          reg123 : reg592) != (forvar587 >>> reg685))));
                      reg667 <= ((reg569 ?
                              $signed((reg568 <= reg658)) : forvar531) ?
                          reg175 : forvar640);
                    end
                  else
                    begin
                      reg664 <= reg563[(2'h3):(1'h0)];
                      reg665 <= {{$signed(reg169)}};
                    end
                end
              for (forvar668 = (1'h0); (forvar668 < (1'h1)); forvar668 = (forvar668 + (1'h1)))
                begin
                  for (forvar669 = (1'h0); (forvar669 < (2'h3)); forvar669 = (forvar669 + (1'h1)))
                    begin
                      reg670 <= $signed(reg40[(3'h5):(2'h2)]);
                      reg671 <= ($unsigned((^$unsigned((8'haa)))) >= $signed($signed($signed((8'h9f)))));
                      reg672 <= {((reg180[(1'h1):(1'h0)] - $signed(reg654)) < (8'ha9))};
                      reg673 <= ($unsigned(({reg168} >= (reg639 <= reg81))) ?
                          $unsigned($signed((reg501 << reg538))) : (^(+(reg507 ^~ (8'hac)))));
                    end
                  reg674 <= ({reg211} & $unsigned((8'ha9)));
                end
            end
        end
    end
  assign wire707 = reg165;
  assign wire708 = (((~^$signed(reg495)) ?
                       (reg159[(1'h0):(1'h0)] ?
                           (&reg144) : (reg97 >>> reg628)) : $unsigned(reg23)) <= ($signed((|reg631)) && reg120));
  always
    @(posedge clk) begin
      if ((reg558[(1'h0):(1'h0)] ?
          {reg66[(4'hb):(1'h0)]} : (|$unsigned(((8'h9e) ? (8'hb7) : reg186)))))
        begin
          if (((reg51[(4'h9):(3'h6)] << $unsigned($unsigned(reg655))) ?
              {$unsigned((^reg37))} : $unsigned($signed((reg595 ^~ reg631)))))
            begin
              reg709 <= reg184[(3'h7):(1'h0)];
            end
          else
            begin
              for (forvar709 = (1'h0); (forvar709 < (1'h0)); forvar709 = (forvar709 + (1'h1)))
                begin
                  if ((reg571 * (reg82 ?
                      (reg667[(3'h5):(3'h5)] ^~ (reg206 > reg689)) : $unsigned((!reg600)))))
                    begin
                      reg710 <= reg520[(4'h8):(3'h4)];
                      reg711 <= (~^reg132);
                      reg712 <= $signed((wire6 ?
                          reg111[(2'h2):(1'h0)] : (reg679 ?
                              (&reg501) : (reg78 ? reg113 : (8'h9d)))));
                      reg713 <= reg68[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg710 <= {(((+reg645) ?
                              $unsigned(reg673) : reg503[(1'h0):(1'h0)]) < (-(reg106 != reg221)))};
                    end
                  for (forvar714 = (1'h0); (forvar714 < (2'h2)); forvar714 = (forvar714 + (1'h1)))
                    begin
                      reg715 <= reg523[(3'h6):(1'h0)];
                      reg716 <= reg639;
                    end
                  if ((8'h9d))
                    begin
                      reg717 <= {{($unsigned(reg612) ?
                                  (reg139 ? reg85 : (8'ha0)) : (8'hb6))}};
                      reg718 <= ({({(8'hac)} ? {reg99} : ((8'hb8) + reg680))} ?
                          (reg521 ?
                              reg174[(1'h0):(1'h0)] : ($unsigned(reg120) ~^ reg659)) : (^{$unsigned(reg195)}));
                    end
                  else
                    begin
                      reg717 <= reg167[(3'h4):(1'h0)];
                      reg718 <= $unsigned(reg667);
                    end
                  reg719 <= ({$unsigned((reg13 ?
                          reg654 : reg152))} >>> (~^$signed(reg710[(1'h1):(1'h1)])));
                end
            end
          if ({$signed(((&reg690) ? ((8'ha9) & (8'h9d)) : $signed(reg520)))})
            begin
              if ({reg90})
                begin
                  for (forvar720 = (1'h0); (forvar720 < (2'h2)); forvar720 = (forvar720 + (1'h1)))
                    begin
                      reg721 <= $unsigned((&((wire708 ?
                          reg580 : (8'ha2)) > reg164)));
                    end
                  for (forvar722 = (1'h0); (forvar722 < (2'h2)); forvar722 = (forvar722 + (1'h1)))
                    begin
                      reg723 <= reg537[(2'h2):(2'h2)];
                    end
                  if ($signed((!$unsigned((reg610 ? reg555 : wire9)))))
                    begin
                      reg724 <= ((((^~reg563) + {reg666}) <<< ((reg684 ?
                              reg706 : reg203) ?
                          $signed(reg127) : (reg629 || wire7))) >= $signed($unsigned({reg579})));
                      reg725 <= reg684;
                    end
                  else
                    begin
                      reg724 <= $unsigned((+((reg225 ? reg580 : reg145) ?
                          reg684[(3'h6):(3'h6)] : reg570[(2'h2):(1'h0)])));
                      reg725 <= reg160[(4'hd):(4'ha)];
                      reg726 <= {($unsigned($signed(reg542)) || reg196[(1'h0):(1'h0)])};
                    end
                end
              else
                begin
                  for (forvar720 = (1'h0); (forvar720 < (1'h1)); forvar720 = (forvar720 + (1'h1)))
                    begin
                      reg721 <= (($signed((reg102 ? reg713 : reg88)) ?
                          (8'hb4) : reg629[(4'hc):(4'hc)]) >> $unsigned($signed((reg56 > reg706))));
                      reg722 <= (^(~&reg47));
                      reg723 <= $signed($unsigned($unsigned({reg535})));
                    end
                end
            end
          else
            begin
              if (reg695[(2'h3):(1'h0)])
                begin
                  reg720 <= ((^reg645[(3'h5):(2'h3)]) + reg512);
                  if ((-$signed(($unsigned(reg592) ? reg225 : (~^reg548)))))
                    begin
                      reg721 <= (($unsigned($unsigned(reg538)) <<< reg719) * $signed($unsigned(reg225[(1'h0):(1'h0)])));
                      reg722 <= reg511[(1'h1):(1'h0)];
                      reg723 <= ($signed(reg197) ?
                          (&reg534[(2'h2):(2'h2)]) : (+$unsigned((reg603 >>> reg591))));
                    end
                  else
                    begin
                      reg721 <= (|reg715[(3'h5):(2'h2)]);
                      reg722 <= (reg515[(1'h0):(1'h0)] + reg510);
                    end
                  for (forvar724 = (1'h0); (forvar724 < (1'h0)); forvar724 = (forvar724 + (1'h1)))
                    begin
                      reg725 <= wire708[(2'h2):(2'h2)];
                    end
                  if ((reg661 ? (|$signed(reg568)) : reg103))
                    begin
                      reg726 <= reg89[(2'h3):(1'h0)];
                      reg727 <= $unsigned(($signed($unsigned(reg661)) * ($signed(reg14) >= (reg156 ?
                          reg206 : reg148))));
                    end
                  else
                    begin
                      reg726 <= $signed($unsigned(reg696));
                    end
                end
              else
                begin
                  for (forvar720 = (1'h0); (forvar720 < (2'h2)); forvar720 = (forvar720 + (1'h1)))
                    begin
                      reg721 <= reg173[(3'h5):(1'h1)];
                    end
                end
              if ($signed($signed((reg68 && (&reg122)))))
                begin
                  if ((reg517[(3'h4):(2'h3)] ?
                      ((|reg14[(4'h8):(4'h8)]) < $signed(((8'hae) ?
                          reg501 : reg635))) : (({reg96} ?
                              $unsigned(reg535) : $unsigned(reg172)) ?
                          $unsigned((reg96 ?
                              reg225 : reg168)) : (~$signed((8'ha6))))))
                    begin
                      reg728 <= reg616[(3'h5):(1'h0)];
                      reg729 <= $signed((|(reg691 & (~reg175))));
                    end
                  else
                    begin
                      reg728 <= {(($unsigned((8'ha4)) * (reg183 ?
                              reg722 : reg536)) < {$signed(reg99)})};
                      reg729 <= (^$signed(((&(8'h9f)) ?
                          reg160 : $signed(reg581))));
                      reg730 <= ($signed($unsigned((reg33 != (8'hb7)))) ?
                          reg97 : {($unsigned(reg66) != ((8'hac) ?
                                  reg553 : reg127))});
                      reg731 <= $unsigned(($unsigned(reg179[(3'h6):(3'h5)]) && ({reg624} ?
                          $signed((8'hb9)) : (&(8'ha9)))));
                    end
                  for (forvar732 = (1'h0); (forvar732 < (1'h1)); forvar732 = (forvar732 + (1'h1)))
                    begin
                      reg733 <= {(^~$signed((reg141 & reg100)))};
                      reg734 <= $unsigned((|(reg613[(2'h2):(1'h0)] ?
                          (8'ha2) : (reg662 ? reg544 : reg694))));
                    end
                  reg735 <= (reg655[(2'h2):(1'h0)] & {$signed(reg150)});
                end
              else
                begin
                  if (reg562[(3'h4):(2'h3)])
                    begin
                      reg728 <= {$signed((+$unsigned(reg190)))};
                    end
                  else
                    begin
                      reg728 <= $signed(reg219[(3'h4):(2'h2)]);
                      reg729 <= (($signed($signed(reg723)) ?
                          ($signed(reg622) == reg687) : ((reg52 ?
                              reg125 : reg530) <<< reg143)) >> (({reg161} >= (+(8'ha4))) ?
                          $unsigned($unsigned(reg639)) : ($signed(reg208) ?
                              (reg163 | wire492) : $signed(reg103))));
                    end
                  for (forvar730 = (1'h0); (forvar730 < (1'h1)); forvar730 = (forvar730 + (1'h1)))
                    begin
                      reg731 <= ({$signed((|reg170))} ?
                          (~|(reg14 || (reg13 ? reg39 : (8'hba)))) : (reg10 ?
                              $signed((reg16 ?
                                  reg99 : reg89)) : reg528[(3'h5):(3'h4)]));
                    end
                end
              for (forvar736 = (1'h0); (forvar736 < (2'h3)); forvar736 = (forvar736 + (1'h1)))
                begin
                  for (forvar737 = (1'h0); (forvar737 < (2'h2)); forvar737 = (forvar737 + (1'h1)))
                    begin
                      reg738 <= $signed((reg690 ?
                          ($signed(reg115) <<< (reg60 ?
                              reg604 : reg190)) : reg129));
                      reg739 <= ($signed(reg589[(3'h6):(3'h4)]) != $signed($signed((reg544 ?
                          (8'haa) : reg145))));
                      reg740 <= reg13;
                      reg741 <= reg559[(1'h0):(1'h0)];
                    end
                  if (({reg515[(2'h3):(1'h1)]} >> ((((8'hac) || reg212) - $signed(reg171)) <= reg624[(1'h0):(1'h0)])))
                    begin
                      reg742 <= (reg211[(4'h8):(2'h2)] ?
                          {$unsigned({reg30})} : ((~^reg698[(2'h3):(2'h2)]) ?
                              (^~{reg78}) : ($unsigned((8'hb2)) ?
                                  {reg164} : reg583[(3'h5):(2'h3)])));
                      reg743 <= $unsigned($signed((-(~reg617))));
                    end
                  else
                    begin
                      reg742 <= reg660;
                      reg743 <= (~&($signed($signed(reg19)) != ((-reg533) ?
                          (reg662 ? reg139 : reg132) : (reg502 > reg518))));
                      reg744 <= (^~(~($signed(reg605) + (8'had))));
                    end
                end
            end
          for (forvar745 = (1'h0); (forvar745 < (1'h1)); forvar745 = (forvar745 + (1'h1)))
            begin
              for (forvar746 = (1'h0); (forvar746 < (2'h3)); forvar746 = (forvar746 + (1'h1)))
                begin
                  reg747 <= reg728[(2'h2):(1'h0)];
                  for (forvar748 = (1'h0); (forvar748 < (1'h0)); forvar748 = (forvar748 + (1'h1)))
                    begin
                      reg749 <= ({reg534[(2'h3):(1'h0)]} ^~ ({{reg170}} ?
                          $unsigned(reg172[(2'h3):(1'h1)]) : $unsigned((reg616 ?
                              reg735 : reg600))));
                      reg750 <= reg187;
                    end
                  reg751 <= {$unsigned($signed(forvar736))};
                  reg752 <= (((8'h9d) >>> (+reg200)) ?
                      (reg38[(2'h2):(1'h0)] ?
                          $unsigned((reg155 ^~ reg114)) : $signed(reg66)) : reg557[(1'h0):(1'h0)]);
                end
              for (forvar753 = (1'h0); (forvar753 < (1'h1)); forvar753 = (forvar753 + (1'h1)))
                begin
                  if ((reg199[(1'h1):(1'h0)] == (reg675 ^ {(reg589 ?
                          reg564 : reg569)})))
                    begin
                      reg754 <= $signed(reg587);
                    end
                  else
                    begin
                      reg754 <= (!reg143[(1'h1):(1'h1)]);
                    end
                end
            end
          reg755 <= ((~^$unsigned((!reg47))) ?
              $signed({reg193[(3'h5):(3'h5)]}) : (~^(reg641 ?
                  $unsigned(reg700) : (~&reg628))));
        end
      else
        begin
          for (forvar709 = (1'h0); (forvar709 < (2'h3)); forvar709 = (forvar709 + (1'h1)))
            begin
              for (forvar710 = (1'h0); (forvar710 < (2'h2)); forvar710 = (forvar710 + (1'h1)))
                begin
                  for (forvar711 = (1'h0); (forvar711 < (1'h0)); forvar711 = (forvar711 + (1'h1)))
                    begin
                      reg712 <= $signed(reg139);
                    end
                  if ((reg21[(1'h1):(1'h0)] == $signed(($signed(reg651) ?
                      reg188 : $unsigned(reg685)))))
                    begin
                      reg713 <= $signed(reg540[(1'h1):(1'h1)]);
                      reg714 <= {reg547};
                      reg715 <= reg666;
                    end
                  else
                    begin
                      reg713 <= ((~^(reg180[(3'h5):(2'h2)] == (reg613 ?
                          (8'hb4) : reg41))) <<< ($unsigned($unsigned(reg741)) || $unsigned((reg167 ?
                          reg113 : reg90))));
                      reg714 <= ((-reg660) ?
                          reg140 : (reg173[(1'h0):(1'h0)] ?
                              reg590[(4'hd):(4'hd)] : (forvar748 ?
                                  $signed(reg95) : reg194)));
                    end
                  reg716 <= $unsigned($unsigned($unsigned($signed(reg511))));
                end
              for (forvar717 = (1'h0); (forvar717 < (1'h0)); forvar717 = (forvar717 + (1'h1)))
                begin
                  if (reg50)
                    begin
                      reg718 <= ({reg524[(2'h3):(2'h2)]} ?
                          (($signed(reg60) & (+reg116)) >>> reg545) : (((reg551 ?
                                  forvar722 : reg88) ~^ (8'hb7)) ?
                              {$signed(forvar710)} : $signed($unsigned(reg713))));
                    end
                  else
                    begin
                      reg718 <= (reg740 & reg104[(4'hd):(2'h2)]);
                    end
                  for (forvar719 = (1'h0); (forvar719 < (2'h2)); forvar719 = (forvar719 + (1'h1)))
                    begin
                      reg720 <= ($signed({$signed(reg185)}) ?
                          ($unsigned($signed((8'ha7))) ?
                              {(reg710 > reg47)} : $unsigned(reg591)) : reg21[(3'h5):(3'h5)]);
                      reg721 <= $unsigned(reg545[(3'h5):(3'h5)]);
                      reg722 <= reg102;
                    end
                  reg723 <= reg729[(1'h1):(1'h0)];
                  if ({(~(&reg635))})
                    begin
                      reg724 <= $unsigned($signed(((reg40 ?
                          reg188 : reg754) + $unsigned(reg717))));
                      reg725 <= (&$signed(reg655[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg724 <= (8'ha5);
                      reg725 <= reg178;
                    end
                end
              reg726 <= (reg214 ?
                  $signed($signed($unsigned(reg720))) : ($unsigned(reg129[(4'hd):(3'h7)]) ?
                      reg174[(2'h2):(1'h0)] : ((reg542 ^ forvar748) > (8'hb2))));
            end
          if ((8'hba))
            begin
              for (forvar727 = (1'h0); (forvar727 < (1'h1)); forvar727 = (forvar727 + (1'h1)))
                begin
                  reg728 <= $signed((~^(reg553 ? reg596 : (~|reg657))));
                end
              for (forvar729 = (1'h0); (forvar729 < (1'h1)); forvar729 = (forvar729 + (1'h1)))
                begin
                  for (forvar730 = (1'h0); (forvar730 < (1'h1)); forvar730 = (forvar730 + (1'h1)))
                    begin
                      reg731 <= $signed($signed($unsigned((reg545 ?
                          reg217 : reg644))));
                      reg732 <= reg101[(3'h4):(1'h0)];
                      reg733 <= ((({reg17} ? {reg44} : (!forvar737)) ?
                          (+$unsigned((8'hb5))) : $unsigned($signed(reg727))) * {$signed(reg151)});
                      reg734 <= (reg730 ? reg563[(1'h1):(1'h1)] : reg201);
                    end
                  reg735 <= ((((forvar709 ? reg671 : reg147) ?
                      (~&reg174) : (reg172 ?
                          reg45 : (8'haf))) >= $signed(reg730[(2'h3):(1'h1)])) <<< $unsigned($unsigned((+(8'hb8)))));
                  for (forvar736 = (1'h0); (forvar736 < (1'h0)); forvar736 = (forvar736 + (1'h1)))
                    begin
                      reg737 <= ($signed(forvar730) && reg599);
                    end
                  for (forvar738 = (1'h0); (forvar738 < (2'h2)); forvar738 = (forvar738 + (1'h1)))
                    begin
                      reg739 <= ((reg22[(3'h7):(3'h4)] * $signed((reg714 ?
                              reg733 : (8'hba)))) ?
                          reg604 : (8'h9d));
                      reg740 <= $unsigned(($signed({reg23}) << (!reg107)));
                      reg741 <= $unsigned($unsigned($unsigned($unsigned(reg725))));
                      reg742 <= ($unsigned(reg38) | reg752);
                    end
                end
              for (forvar743 = (1'h0); (forvar743 < (1'h1)); forvar743 = (forvar743 + (1'h1)))
                begin
                  for (forvar744 = (1'h0); (forvar744 < (1'h1)); forvar744 = (forvar744 + (1'h1)))
                    begin
                      reg745 <= (reg556[(2'h2):(1'h0)] ?
                          reg643[(1'h1):(1'h1)] : (forvar724 << (~&$signed(reg591))));
                      reg746 <= ((~&$unsigned(reg631[(4'h8):(3'h5)])) ?
                          {$signed(reg693[(1'h1):(1'h0)])} : (^({reg751} ?
                              (reg727 ?
                                  reg548 : (8'ha3)) : reg659[(3'h6):(3'h5)])));
                      reg747 <= {$unsigned((~^(&reg588)))};
                      reg748 <= (!reg159);
                    end
                  for (forvar749 = (1'h0); (forvar749 < (1'h1)); forvar749 = (forvar749 + (1'h1)))
                    begin
                      reg750 <= (reg161 ?
                          $unsigned(($unsigned(wire6) != $unsigned(reg715))) : $signed($signed($unsigned((8'h9f)))));
                      reg751 <= reg82;
                    end
                  if (reg750)
                    begin
                      reg752 <= (~&$signed($signed($signed((8'hb5)))));
                      reg753 <= (reg210[(3'h6):(1'h1)] ?
                          {reg127[(2'h2):(1'h0)]} : ((reg739 != (reg81 | reg746)) ?
                              ($signed(reg683) ?
                                  $unsigned((8'hb6)) : (~reg702)) : {(reg178 ?
                                      reg84 : reg121)}));
                    end
                  else
                    begin
                      reg752 <= $signed(reg526[(1'h0):(1'h0)]);
                      reg753 <= reg537[(1'h1):(1'h0)];
                      reg754 <= reg105[(2'h2):(1'h1)];
                    end
                  if ((reg533 ?
                      (reg637[(2'h3):(2'h2)] ?
                          reg652[(3'h5):(3'h4)] : $signed((reg82 - (8'ha2)))) : (~&$signed((|reg159)))))
                    begin
                      reg755 <= ({($signed(reg90) | (reg554 < reg699))} ?
                          reg683 : (((reg637 ? (8'had) : reg722) > (reg729 ?
                              reg646 : reg210)) && ($signed((8'ha4)) < reg23)));
                    end
                  else
                    begin
                      reg755 <= $unsigned(reg145);
                    end
                end
              if ($unsigned($signed(reg134)))
                begin
                  for (forvar756 = (1'h0); (forvar756 < (1'h0)); forvar756 = (forvar756 + (1'h1)))
                    begin
                      reg757 <= (8'hb3);
                      reg758 <= reg530;
                      reg759 <= ($unsigned(((reg564 ?
                          (8'h9c) : reg64) >> (8'hba))) | reg68[(1'h0):(1'h0)]);
                    end
                  if ((~^$signed(wire8)))
                    begin
                      reg760 <= $unsigned(($unsigned(reg21[(2'h3):(2'h2)]) & (~^(reg141 >> reg514))));
                      reg761 <= reg663[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg760 <= {{($signed(reg720) ?
                                  reg633 : (reg69 ? wire708 : reg41))}};
                      reg761 <= $signed($unsigned(reg114[(3'h4):(1'h0)]));
                    end
                  for (forvar762 = (1'h0); (forvar762 < (1'h1)); forvar762 = (forvar762 + (1'h1)))
                    begin
                      reg763 <= ((reg196 ? reg595 : reg573) ?
                          reg165 : ($unsigned($signed((8'hac))) ?
                              (+(-reg511)) : $signed({(8'hb3)})));
                      reg764 <= {($signed(reg115) ?
                              $unsigned((~^reg77)) : (!reg629[(1'h0):(1'h0)]))};
                    end
                  if (reg190[(3'h5):(3'h4)])
                    begin
                      reg765 <= reg726[(2'h2):(1'h0)];
                      reg766 <= (~|reg590[(4'hd):(3'h6)]);
                    end
                  else
                    begin
                      reg765 <= (!$signed((~(~^reg186))));
                      reg766 <= reg218[(1'h1):(1'h1)];
                      reg767 <= ($unsigned($signed($unsigned(reg145))) ?
                          reg526 : reg177[(2'h3):(1'h1)]);
                    end
                end
              else
                begin
                  if ((!(reg755[(4'he):(2'h3)] ?
                      ((&reg717) ? (~^reg763) : reg554) : $signed((8'had)))))
                    begin
                      reg756 <= $signed(($signed({reg729}) <= reg739));
                      reg757 <= $signed($signed(reg197[(3'h7):(2'h2)]));
                    end
                  else
                    begin
                      reg756 <= (-((8'h9c) ?
                          $signed($signed(reg716)) : ({reg608} ?
                              (^reg681) : (^reg665))));
                      reg757 <= wire9[(4'hd):(3'h4)];
                      reg758 <= $unsigned((~&reg102));
                      reg759 <= $signed(($unsigned(reg535) >> ((reg657 ?
                          reg734 : reg126) | (reg582 >>> reg213))));
                    end
                  for (forvar760 = (1'h0); (forvar760 < (1'h1)); forvar760 = (forvar760 + (1'h1)))
                    begin
                      reg761 <= $unsigned(($signed((reg711 - reg118)) * (reg162 ?
                          ((8'hb8) ? reg537 : reg559) : $unsigned(reg759))));
                    end
                  reg762 <= (({{(8'ha7)}} == ((^~reg503) ~^ (reg503 ?
                          reg666 : reg70))) ?
                      $unsigned({(wire492 ^ reg562)}) : ($unsigned($unsigned(reg104)) ?
                          (8'hb1) : $signed((|(8'ha9)))));
                  for (forvar763 = (1'h0); (forvar763 < (2'h3)); forvar763 = (forvar763 + (1'h1)))
                    begin
                      reg764 <= ((^(8'ha3)) ?
                          (8'hb7) : (((reg18 < reg757) ?
                              (8'hab) : (reg547 ? reg732 : reg184)) >> reg636));
                      reg765 <= reg746[(1'h1):(1'h1)];
                      reg766 <= {(~^(forvar729[(4'h8):(2'h3)] ?
                              (reg538 ? reg636 : reg749) : (8'hb8)))};
                      reg767 <= ($signed((^((8'haa) && reg27))) ?
                          $unsigned((&((8'hb8) ?
                              (8'had) : reg205))) : $unsigned(($unsigned(reg726) ?
                              $signed((8'h9e)) : $signed(reg47))));
                    end
                end
            end
          else
            begin
              if ({(!reg56[(4'hb):(2'h3)])})
                begin
                  reg727 <= (^(~&reg64[(1'h0):(1'h0)]));
                end
              else
                begin
                  for (forvar727 = (1'h0); (forvar727 < (2'h2)); forvar727 = (forvar727 + (1'h1)))
                    begin
                      reg728 <= $unsigned((reg752 == ({reg103} << (reg713 <<< reg678))));
                      reg729 <= (+((~&$signed(reg207)) & forvar711[(3'h5):(1'h0)]));
                      reg730 <= ({((reg636 ^ reg114) && $unsigned(reg50))} == ((^~$unsigned(reg689)) ?
                          $unsigned((reg78 ?
                              (8'had) : (8'ha7))) : $unsigned(reg129)));
                    end
                end
            end
          if ((reg706[(1'h0):(1'h0)] ?
              (&$unsigned(forvar763[(3'h6):(2'h3)])) : reg634))
            begin
              for (forvar768 = (1'h0); (forvar768 < (1'h1)); forvar768 = (forvar768 + (1'h1)))
                begin
                  if ((&(($signed(reg159) ?
                      reg513 : reg529[(4'ha):(3'h7)]) < ($signed(reg671) ?
                      reg516[(1'h0):(1'h0)] : $signed(forvar717)))))
                    begin
                      reg769 <= (reg183[(1'h0):(1'h0)] ?
                          (reg718[(3'h5):(2'h2)] ?
                              (~^reg208) : reg83) : reg565[(1'h1):(1'h1)]);
                      reg770 <= ($unsigned($signed({reg712})) + (~&forvar745));
                      reg771 <= {(|(^reg525[(3'h6):(3'h5)]))};
                    end
                  else
                    begin
                      reg769 <= reg562;
                    end
                end
            end
          else
            begin
              reg768 <= reg758[(4'h8):(2'h2)];
              for (forvar769 = (1'h0); (forvar769 < (1'h0)); forvar769 = (forvar769 + (1'h1)))
                begin
                  reg770 <= ((~|reg687[(4'h9):(1'h1)]) ?
                      $unsigned(($signed(reg173) | (reg724 ?
                          wire6 : reg567))) : $unsigned((reg505 <= (reg670 ?
                          reg673 : reg564))));
                  if ((8'ha3))
                    begin
                      reg771 <= {$signed(({reg765} ?
                              reg201[(2'h3):(2'h2)] : reg655))};
                      reg772 <= (8'ha3);
                      reg773 <= forvar737[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg771 <= (!{$unsigned(reg761[(3'h4):(2'h3)])});
                      reg772 <= (($signed((reg624 != reg143)) ?
                              ($unsigned((8'ha3)) ~^ (reg178 ?
                                  reg114 : reg147)) : ((~reg193) >> $signed((8'h9e)))) ?
                          (reg97[(3'h5):(3'h4)] ?
                              ((reg684 ? reg679 : reg55) <= (reg205 ?
                                  reg710 : reg713)) : reg89) : reg191);
                    end
                end
              reg774 <= $signed($unsigned((8'hae)));
              reg775 <= $signed($unsigned($signed(reg734[(1'h0):(1'h0)])));
            end
          for (forvar776 = (1'h0); (forvar776 < (1'h1)); forvar776 = (forvar776 + (1'h1)))
            begin
              for (forvar777 = (1'h0); (forvar777 < (1'h0)); forvar777 = (forvar777 + (1'h1)))
                begin
                  for (forvar778 = (1'h0); (forvar778 < (2'h3)); forvar778 = (forvar778 + (1'h1)))
                    begin
                      reg779 <= reg79[(2'h3):(2'h3)];
                      reg780 <= $unsigned(($signed((reg169 >> reg142)) ?
                          (reg651 ? {reg107} : $unsigned(reg213)) : reg51));
                      reg781 <= $unsigned(reg92);
                    end
                  reg782 <= (!($signed((!reg734)) && reg174[(1'h0):(1'h0)]));
                end
            end
        end
      if (reg581)
        begin
          for (forvar783 = (1'h0); (forvar783 < (1'h1)); forvar783 = (forvar783 + (1'h1)))
            begin
              if (($unsigned((reg74 ?
                  $signed(forvar743) : $signed(reg749))) * reg686))
                begin
                  reg784 <= ($unsigned($signed($signed(reg675))) ?
                      ((8'ha7) ?
                          (-(^~reg768)) : reg88[(4'h9):(2'h3)]) : reg734[(1'h0):(1'h0)]);
                  for (forvar785 = (1'h0); (forvar785 < (2'h2)); forvar785 = (forvar785 + (1'h1)))
                    begin
                      reg786 <= $signed(((+$unsigned(reg768)) ?
                          {reg743} : $unsigned(((8'hb7) ? reg748 : (8'hb2)))));
                      reg787 <= reg128[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  if ($signed({(reg212 <<< reg715[(1'h0):(1'h0)])}))
                    begin
                      reg784 <= reg732[(4'ha):(3'h5)];
                      reg785 <= reg779[(3'h5):(1'h1)];
                      reg786 <= ($unsigned(((!reg193) ? reg668 : (+reg124))) ?
                          (!($unsigned(reg197) << {(8'hb9)})) : $unsigned(($signed(reg514) ^ $signed(reg705))));
                    end
                  else
                    begin
                      reg784 <= (&$unsigned(reg77[(3'h7):(3'h7)]));
                      reg785 <= (((+$signed(reg47)) - (~(~reg731))) < $unsigned((|$signed(reg566))));
                      reg786 <= $signed(reg755[(4'he):(2'h2)]);
                    end
                  for (forvar787 = (1'h0); (forvar787 < (2'h3)); forvar787 = (forvar787 + (1'h1)))
                    begin
                      reg788 <= $signed((((reg102 - reg656) && (reg526 ?
                              forvar783 : reg196)) ?
                          (reg716[(2'h3):(2'h2)] ?
                              $signed(reg97) : reg583[(1'h1):(1'h1)]) : (-(reg635 ?
                              reg165 : reg177))));
                      reg789 <= reg108;
                    end
                  if ((8'hb0))
                    begin
                      reg790 <= $unsigned(reg710[(1'h1):(1'h0)]);
                      reg791 <= $signed(reg105[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg790 <= reg66[(1'h1):(1'h0)];
                      reg791 <= $unsigned($unsigned(reg32));
                    end
                end
              reg792 <= ($unsigned((~|reg531)) ^~ reg149);
            end
          if ($unsigned($unsigned(reg705[(3'h5):(1'h0)])))
            begin
              for (forvar793 = (1'h0); (forvar793 < (1'h1)); forvar793 = (forvar793 + (1'h1)))
                begin
                  if ($unsigned((($signed((8'h9c)) ^ reg562) ?
                      {reg751} : {$unsigned(reg55)})))
                    begin
                      reg794 <= ($unsigned((8'ha4)) ?
                          reg51[(3'h4):(2'h2)] : $unsigned((-$signed(reg568))));
                      reg795 <= $signed(reg109[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg794 <= $signed((^~reg74[(1'h0):(1'h0)]));
                      reg795 <= ($unsigned(((~reg156) >= (~^reg552))) ?
                          reg37 : $signed({((8'hb4) || reg788)}));
                    end
                  for (forvar796 = (1'h0); (forvar796 < (2'h2)); forvar796 = (forvar796 + (1'h1)))
                    begin
                      reg797 <= (8'hb9);
                    end
                  for (forvar798 = (1'h0); (forvar798 < (1'h0)); forvar798 = (forvar798 + (1'h1)))
                    begin
                      reg799 <= reg757;
                      reg800 <= (8'hb5);
                      reg801 <= $unsigned((~reg514[(2'h3):(1'h0)]));
                      reg802 <= $unsigned(({reg213} ?
                          (reg503[(3'h5):(3'h4)] ^ reg677[(3'h5):(2'h2)]) : (~^reg699)));
                    end
                end
              if ($unsigned((~(reg663[(2'h2):(1'h1)] ?
                  $unsigned((8'ha2)) : $unsigned(reg16)))))
                begin
                  reg803 <= ($signed((((8'hb1) && reg117) ?
                      $signed(reg704) : ((8'ha0) ^ reg225))) ^ reg741);
                  reg804 <= reg200;
                end
              else
                begin
                  for (forvar803 = (1'h0); (forvar803 < (2'h3)); forvar803 = (forvar803 + (1'h1)))
                    begin
                      reg804 <= $unsigned(((reg110 - $signed(reg191)) ?
                          $unsigned(reg505[(4'hb):(3'h6)]) : (|reg660[(4'hf):(2'h2)])));
                    end
                  if ((8'haf))
                    begin
                      reg805 <= forvar746[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg805 <= $unsigned((reg121 <= reg126));
                      reg806 <= (reg759 && {$unsigned(reg204)});
                      reg807 <= $unsigned(reg556[(1'h0):(1'h0)]);
                      reg808 <= reg213;
                    end
                end
              for (forvar809 = (1'h0); (forvar809 < (1'h1)); forvar809 = (forvar809 + (1'h1)))
                begin
                  for (forvar810 = (1'h0); (forvar810 < (2'h2)); forvar810 = (forvar810 + (1'h1)))
                    begin
                      reg811 <= ($unsigned(($unsigned(reg756) ~^ $unsigned(reg506))) ?
                          reg157 : (reg497 < ({reg615} ?
                              reg656[(1'h0):(1'h0)] : reg218)));
                    end
                end
            end
          else
            begin
              if (reg744)
                begin
                  for (forvar793 = (1'h0); (forvar793 < (2'h3)); forvar793 = (forvar793 + (1'h1)))
                    begin
                      reg794 <= (reg789[(2'h3):(2'h2)] * (8'hb5));
                      reg795 <= (reg102 ?
                          {(8'haf)} : $signed(({reg552} ?
                              (^forvar785) : (~|reg562))));
                      reg796 <= ((reg616[(1'h1):(1'h0)] == reg40) <= ($signed($unsigned(reg668)) > $unsigned(reg591)));
                    end
                  for (forvar797 = (1'h0); (forvar797 < (1'h0)); forvar797 = (forvar797 + (1'h1)))
                    begin
                      reg798 <= reg760;
                      reg799 <= $unsigned(reg189[(3'h4):(2'h2)]);
                    end
                end
              else
                begin
                  reg793 <= {reg662};
                  reg794 <= ((reg22[(3'h7):(3'h7)] ^~ reg793) ?
                      $signed($signed((forvar729 ?
                          reg538 : reg194))) : (8'ha5));
                end
            end
          if ((((reg786 * (~^(8'hb3))) >> (-$unsigned(reg686))) ?
              (reg556 ?
                  reg578[(1'h0):(1'h0)] : ($signed(reg662) - forvar724)) : $unsigned($unsigned((reg514 ?
                  reg170 : reg143)))))
            begin
              if ((^~$signed(reg135[(1'h1):(1'h1)])))
                begin
                  for (forvar812 = (1'h0); (forvar812 < (2'h2)); forvar812 = (forvar812 + (1'h1)))
                    begin
                      reg813 <= $signed({(reg45 != reg184)});
                      reg814 <= (~&(($signed(reg656) + $unsigned(reg183)) > reg60));
                    end
                  if ({(|$unsigned((|reg785)))})
                    begin
                      reg815 <= reg544[(4'hb):(4'ha)];
                      reg816 <= $signed(($unsigned($unsigned(reg512)) - $unsigned((!reg647))));
                      reg817 <= $unsigned(reg41[(3'h5):(3'h5)]);
                      reg818 <= (8'ha0);
                    end
                  else
                    begin
                      reg815 <= {(reg175[(2'h2):(2'h2)] ?
                              ({forvar722} ?
                                  $signed(reg742) : (reg18 == reg517)) : reg199[(1'h0):(1'h0)])};
                      reg816 <= $unsigned(((^(reg519 && (8'hb0))) || reg602[(4'ha):(2'h3)]));
                      reg817 <= $signed((((reg526 ^ reg208) != {reg596}) && reg691[(1'h1):(1'h0)]));
                    end
                  reg819 <= reg200[(3'h4):(3'h4)];
                  reg820 <= wire6[(4'h9):(3'h4)];
                end
              else
                begin
                  for (forvar812 = (1'h0); (forvar812 < (1'h0)); forvar812 = (forvar812 + (1'h1)))
                    begin
                      reg813 <= $signed($signed((~reg143)));
                      reg814 <= reg604[(1'h0):(1'h0)];
                      reg815 <= ($signed({(~reg148)}) + reg27[(1'h0):(1'h0)]);
                      reg816 <= $unsigned(reg140);
                    end
                  if ($signed(((~&reg34) ?
                      $unsigned((^reg151)) : (reg508 << (8'hb8)))))
                    begin
                      reg817 <= $unsigned((~$unsigned((reg171 + reg635))));
                      reg818 <= reg215;
                      reg819 <= reg645;
                    end
                  else
                    begin
                      reg817 <= {(+(reg537[(2'h2):(1'h1)] == $signed(reg68)))};
                      reg818 <= $unsigned($unsigned((!(reg733 - reg60))));
                    end
                  if ((8'ha8))
                    begin
                      reg820 <= (~({reg743} + ($unsigned(reg113) || forvar783[(2'h3):(2'h3)])));
                      reg821 <= $unsigned(reg629[(3'h4):(2'h2)]);
                      reg822 <= (-(~^$unsigned(reg528)));
                      reg823 <= ({(reg64[(3'h5):(2'h3)] ?
                              (reg523 >>> (8'hac)) : $unsigned(reg130))} ^~ (((reg88 <<< reg791) * wire708) >= $unsigned($signed(reg674))));
                    end
                  else
                    begin
                      reg820 <= reg216[(1'h1):(1'h0)];
                      reg821 <= {{reg219[(1'h1):(1'h1)]}};
                      reg822 <= reg131;
                      reg823 <= ((~|reg519[(1'h0):(1'h0)]) ^~ $signed((!$signed(reg639))));
                    end
                  reg824 <= ({$signed($unsigned((8'hab)))} ?
                      $signed($unsigned((|forvar738))) : (^~reg699[(2'h3):(1'h1)]));
                end
            end
          else
            begin
              for (forvar812 = (1'h0); (forvar812 < (1'h1)); forvar812 = (forvar812 + (1'h1)))
                begin
                  if (reg162[(2'h2):(2'h2)])
                    begin
                      reg813 <= reg543;
                      reg814 <= $unsigned((+(reg172[(4'hc):(4'h8)] << $signed(reg647))));
                      reg815 <= $signed(($signed((reg681 << reg186)) ?
                          reg651 : reg726[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg813 <= ((8'ha8) ? reg38 : ((8'h9f) - reg590));
                      reg814 <= ((8'had) ?
                          (~|forvar743[(3'h5):(1'h0)]) : reg704[(1'h0):(1'h0)]);
                      reg815 <= reg503;
                    end
                  if (reg741[(3'h5):(3'h4)])
                    begin
                      reg816 <= $signed((~&($signed(reg606) || reg516)));
                    end
                  else
                    begin
                      reg816 <= $unsigned((~|(reg576 ?
                          reg791[(3'h5):(1'h1)] : (reg691 ?
                              forvar709 : reg89))));
                    end
                end
              reg817 <= {$unsigned($signed($unsigned((8'had))))};
              for (forvar818 = (1'h0); (forvar818 < (1'h0)); forvar818 = (forvar818 + (1'h1)))
                begin
                  for (forvar819 = (1'h0); (forvar819 < (1'h1)); forvar819 = (forvar819 + (1'h1)))
                    begin
                      reg820 <= {((~&{(8'hba)}) > $signed($unsigned((8'ha2))))};
                      reg821 <= reg516;
                      reg822 <= reg538[(3'h4):(1'h1)];
                      reg823 <= ($signed((|reg83)) >>> (reg747[(2'h2):(1'h0)] ^ {((8'ha6) << reg799)}));
                    end
                end
            end
        end
      else
        begin
          if ({reg518[(3'h7):(3'h4)]})
            begin
              for (forvar783 = (1'h0); (forvar783 < (1'h1)); forvar783 = (forvar783 + (1'h1)))
                begin
                  for (forvar784 = (1'h0); (forvar784 < (2'h3)); forvar784 = (forvar784 + (1'h1)))
                    begin
                      reg785 <= $signed($signed(((reg114 | reg592) ?
                          (reg564 ? (8'hae) : reg141) : {reg786})));
                    end
                  for (forvar786 = (1'h0); (forvar786 < (1'h1)); forvar786 = (forvar786 + (1'h1)))
                    begin
                      reg787 <= ((~|((reg196 ? (8'hb5) : (8'hac)) * reg125)) ?
                          ($signed($signed(reg90)) ?
                              ((8'hac) ^~ $signed(reg799)) : (reg134[(3'h4):(1'h0)] >> $signed(reg681))) : $signed({(-reg141)}));
                    end
                end
              if (($unsigned($signed((reg97 ? reg802 : reg38))) * reg747))
                begin
                  if ($signed({reg164}))
                    begin
                      reg788 <= reg151[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg788 <= {($unsigned(((8'had) ? (8'h9f) : reg78)) ?
                              $unsigned($signed(reg595)) : reg125[(2'h3):(2'h2)])};
                      reg789 <= ($unsigned(reg162[(2'h2):(1'h1)]) ?
                          $unsigned((&reg198[(1'h1):(1'h0)])) : ($unsigned(reg199[(2'h2):(1'h1)]) + $unsigned({reg117})));
                      reg790 <= reg595;
                      reg791 <= (~$signed((reg558[(2'h2):(1'h0)] >> (reg44 | reg634))));
                    end
                  for (forvar792 = (1'h0); (forvar792 < (1'h1)); forvar792 = (forvar792 + (1'h1)))
                    begin
                      reg793 <= reg88;
                      reg794 <= $unsigned((8'hb6));
                      reg795 <= ((~&$unsigned(reg600[(2'h2):(1'h0)])) ?
                          $unsigned($unsigned((~|reg34))) : reg699[(3'h5):(3'h4)]);
                    end
                  for (forvar796 = (1'h0); (forvar796 < (2'h3)); forvar796 = (forvar796 + (1'h1)))
                    begin
                      reg797 <= {({(reg42 ? reg713 : reg78)} ?
                              {(8'hb9)} : $unsigned($unsigned(reg152)))};
                      reg798 <= $unsigned(wire707[(2'h3):(2'h2)]);
                      reg799 <= reg148;
                      reg800 <= ($unsigned($signed((^~reg216))) ?
                          $signed((reg791[(4'hc):(4'h8)] > {reg75})) : reg654);
                    end
                  if (reg69)
                    begin
                      reg801 <= (8'hb2);
                      reg802 <= ({reg547} * (^~$signed((reg758 ?
                          reg185 : reg763))));
                      reg803 <= reg808[(3'h4):(1'h0)];
                      reg804 <= ($unsigned($unsigned((8'hab))) ?
                          ($unsigned((&reg663)) ^ reg546) : {($signed(reg662) & $signed(reg207))});
                    end
                  else
                    begin
                      reg801 <= reg504[(4'h9):(2'h3)];
                      reg802 <= {({(8'ha4)} >= ($unsigned((8'h9c)) ?
                              (reg118 && reg592) : (reg608 ? reg36 : reg40)))};
                    end
                end
              else
                begin
                  if (reg564)
                    begin
                      reg788 <= (reg605 != $unsigned(forvar719));
                      reg789 <= (reg529[(1'h0):(1'h0)] ?
                          {($signed((8'ha9)) ~^ (reg38 ?
                                  (8'hab) : reg816))} : reg787);
                      reg790 <= {reg186[(3'h7):(2'h2)]};
                    end
                  else
                    begin
                      reg788 <= $signed((!{(reg534 ? (8'hb3) : wire708)}));
                      reg789 <= $signed(reg134);
                      reg790 <= $signed(reg203);
                      reg791 <= $unsigned(((((8'h9d) ? reg597 : reg680) ?
                              (reg811 ? reg215 : reg759) : {reg107}) ?
                          (reg166[(2'h2):(1'h1)] < (reg26 ?
                              reg176 : reg605)) : (reg512 ?
                              $unsigned((8'hb4)) : $signed(reg604))));
                    end
                end
            end
          else
            begin
              reg783 <= ((!$signed(reg547[(1'h0):(1'h0)])) * ($unsigned($signed(reg147)) == (|(reg193 == reg55))));
            end
        end
      for (forvar825 = (1'h0); (forvar825 < (2'h3)); forvar825 = (forvar825 + (1'h1)))
        begin
          for (forvar826 = (1'h0); (forvar826 < (2'h3)); forvar826 = (forvar826 + (1'h1)))
            begin
              for (forvar827 = (1'h0); (forvar827 < (1'h0)); forvar827 = (forvar827 + (1'h1)))
                begin
                  if ({(reg626 ?
                          $signed($signed(reg66)) : $signed(reg162[(1'h0):(1'h0)]))})
                    begin
                      reg828 <= (reg123[(3'h7):(2'h3)] | {$signed((~^reg639))});
                      reg829 <= reg696;
                    end
                  else
                    begin
                      reg828 <= (reg644 > (reg88 ?
                          $unsigned(reg695[(1'h1):(1'h1)]) : (|(reg116 ?
                              reg796 : forvar720))));
                      reg829 <= ($signed({{forvar784}}) + $signed($signed((reg109 ~^ reg36))));
                      reg830 <= ((($signed(reg677) ?
                              reg113[(3'h5):(1'h0)] : (~reg26)) ?
                          reg114 : ($unsigned(reg651) + reg683)) <<< (((reg570 ?
                              reg691 : forvar749) ?
                          $signed(reg529) : $signed(reg706)) >= ((!reg208) ?
                          (&reg784) : {reg688})));
                      reg831 <= $signed($unsigned(reg78[(1'h1):(1'h0)]));
                    end
                  if ($signed({(|(reg578 && reg768))}))
                    begin
                      reg832 <= ($signed((!$signed(reg757))) < (reg185 ?
                          $unsigned((reg728 == reg547)) : (reg616 ?
                              (~reg207) : (+forvar784))));
                      reg833 <= (reg555[(3'h4):(2'h2)] <<< ($unsigned((reg552 * (8'ha3))) >= (^~$signed(reg501))));
                      reg834 <= $signed($signed({(reg131 ? reg645 : (8'hb5))}));
                    end
                  else
                    begin
                      reg832 <= ((reg494 >>> reg692) ^ (reg149[(3'h4):(2'h2)] ?
                          reg103[(4'hc):(3'h6)] : ($unsigned(reg615) > (wire492 ?
                              reg603 : (8'hb3)))));
                      reg833 <= reg528;
                    end
                  reg835 <= reg763[(4'hc):(2'h3)];
                  reg836 <= $unsigned(($signed($signed(reg547)) < $unsigned((reg27 ?
                      reg171 : reg101))));
                end
              reg837 <= ((~&$unsigned(reg583[(4'h8):(2'h2)])) ~^ $signed((-reg89)));
              if (((($unsigned(reg21) | (reg217 <<< reg32)) && {(8'ha1)}) << (8'ha4)))
                begin
                  if ({(reg495 <<< reg643[(2'h2):(1'h0)])})
                    begin
                      reg838 <= $signed((^~(~^reg582)));
                      reg839 <= reg210;
                    end
                  else
                    begin
                      reg838 <= $signed(($signed($signed(reg115)) && $signed({reg646})));
                      reg839 <= {(!(8'haa))};
                      reg840 <= (|$unsigned($signed(forvar777[(3'h6):(2'h3)])));
                      reg841 <= (wire8 >>> (reg598[(1'h1):(1'h0)] ?
                          (reg222 ?
                              $unsigned(reg801) : $signed(reg581)) : (reg191 - $unsigned((8'hb8)))));
                    end
                end
              else
                begin
                  if ({$signed($signed(reg815[(4'hc):(2'h3)]))})
                    begin
                      reg838 <= {$unsigned(((reg98 ?
                              reg702 : reg720) <= (&reg212)))};
                      reg839 <= ((reg533 ~^ reg131) + $unsigned((~^(reg533 ?
                          reg786 : reg77))));
                      reg840 <= reg501;
                      reg841 <= reg615;
                    end
                  else
                    begin
                      reg838 <= reg108;
                      reg839 <= ({(((8'hb9) ? reg583 : reg759) ?
                              (wire6 ?
                                  (8'h9d) : forvar768) : $signed(reg670))} != ($signed(reg189[(2'h3):(1'h0)]) >>> (+$signed(reg785))));
                      reg840 <= (!($signed({reg540}) <<< $signed($signed(reg522))));
                      reg841 <= (forvar803[(2'h3):(2'h3)] ?
                          $unsigned({$signed(reg130)}) : $signed(reg606[(1'h1):(1'h0)]));
                    end
                  if (reg506[(3'h5):(3'h5)])
                    begin
                      reg842 <= $signed($signed((reg213 ?
                          $unsigned(reg124) : reg717[(2'h2):(2'h2)])));
                      reg843 <= ((+((reg83 - forvar753) ?
                          reg45 : (^~forvar746))) ^~ $signed(reg723));
                    end
                  else
                    begin
                      reg842 <= {reg738[(4'hb):(1'h1)]};
                      reg843 <= reg203;
                    end
                  for (forvar844 = (1'h0); (forvar844 < (1'h0)); forvar844 = (forvar844 + (1'h1)))
                    begin
                      reg845 <= $signed(reg752[(4'h8):(2'h3)]);
                      reg846 <= {$signed((~|(-reg222)))};
                      reg847 <= (|$signed($unsigned(((8'hb9) ?
                          (8'haa) : reg534))));
                    end
                  for (forvar848 = (1'h0); (forvar848 < (2'h3)); forvar848 = (forvar848 + (1'h1)))
                    begin
                      reg849 <= (&reg668[(1'h1):(1'h1)]);
                    end
                end
              reg850 <= (~$unsigned(($signed(reg655) << (-(8'hb1)))));
            end
          if ((~&(+((8'hb8) || (forvar784 ? reg157 : reg837)))))
            begin
              if (({{reg573[(1'h0):(1'h0)]}} ?
                  $signed($signed({(8'ha9)})) : (reg19[(1'h1):(1'h1)] ?
                      $unsigned((~^(8'haa))) : {$unsigned(reg738)})))
                begin
                  for (forvar851 = (1'h0); (forvar851 < (1'h0)); forvar851 = (forvar851 + (1'h1)))
                    begin
                      reg852 <= $unsigned(reg688[(1'h1):(1'h1)]);
                    end
                  if (reg763[(4'h8):(4'h8)])
                    begin
                      reg853 <= reg614;
                      reg854 <= ({reg850[(3'h6):(2'h2)]} ? reg689 : reg523);
                      reg855 <= (&reg723);
                    end
                  else
                    begin
                      reg853 <= ((8'hba) ?
                          ((reg107 ^~ reg207) ?
                              (reg750[(3'h4):(1'h0)] ?
                                  forvar753[(2'h2):(1'h0)] : (reg759 != reg539)) : ($signed((8'ha5)) ?
                                  {forvar787} : (reg714 ?
                                      reg599 : reg584))) : ($signed({reg807}) || $unsigned((reg772 ?
                              reg191 : reg822))));
                      reg854 <= (reg615[(2'h3):(1'h0)] ^ reg604[(1'h0):(1'h0)]);
                      reg855 <= reg188[(1'h0):(1'h0)];
                    end
                  if (reg681[(1'h1):(1'h1)])
                    begin
                      reg856 <= (reg648[(4'hb):(4'h8)] ?
                          ((8'ha9) ?
                              reg103 : reg657) : $signed((reg734[(2'h2):(1'h1)] ^~ ((8'hb5) ?
                              reg673 : reg134))));
                      reg857 <= ({reg183} ?
                          $unsigned(reg710) : ({(reg73 << reg837)} && (~^$signed(reg618))));
                      reg858 <= ((((-reg529) ?
                          forvar844[(2'h3):(2'h3)] : $unsigned((8'ha4))) != (!$signed(forvar729))) * (8'h9c));
                    end
                  else
                    begin
                      reg856 <= $unsigned($unsigned((~|$unsigned(reg667))));
                      reg857 <= $signed((({reg692} && reg614) == reg589[(2'h2):(1'h0)]));
                    end
                end
              else
                begin
                  if (($unsigned($unsigned(forvar714)) && (8'hb0)))
                    begin
                      reg851 <= $unsigned(reg89);
                    end
                  else
                    begin
                      reg851 <= {$unsigned((^~reg170[(2'h2):(1'h0)]))};
                      reg852 <= reg83[(1'h0):(1'h0)];
                      reg853 <= (|$signed((8'ha7)));
                    end
                end
            end
          else
            begin
              for (forvar851 = (1'h0); (forvar851 < (2'h3)); forvar851 = (forvar851 + (1'h1)))
                begin
                  if (($signed((~^(+reg506))) ? $signed(reg697) : forvar787))
                    begin
                      reg852 <= $signed($unsigned($unsigned((8'ha1))));
                      reg853 <= reg101;
                      reg854 <= $unsigned((|(^reg540[(2'h2):(2'h2)])));
                    end
                  else
                    begin
                      reg852 <= reg139;
                      reg853 <= reg584[(3'h4):(3'h4)];
                      reg854 <= $unsigned($unsigned($signed({(8'h9d)})));
                      reg855 <= ((+reg746[(5'h10):(4'ha)]) | forvar763);
                    end
                  if (reg794[(4'h9):(3'h6)])
                    begin
                      reg856 <= reg169[(2'h3):(2'h3)];
                      reg857 <= $signed($unsigned(reg596));
                      reg858 <= (!reg598);
                      reg859 <= (reg506 <<< reg688);
                    end
                  else
                    begin
                      reg856 <= $unsigned((|$signed((reg155 > reg770))));
                      reg857 <= (&(!($unsigned(reg828) - (wire492 && reg671))));
                      reg858 <= (reg764[(4'ha):(3'h4)] ?
                          ((reg95 << $unsigned(reg664)) != $unsigned($unsigned(forvar724))) : ({$signed((8'h9c))} && reg102[(2'h2):(1'h1)]));
                      reg859 <= (~^reg732);
                    end
                  reg860 <= reg806;
                  if ((~&$unsigned({$unsigned(reg841)})))
                    begin
                      reg861 <= ((+{reg783[(2'h2):(2'h2)]}) >= ((&(-(8'ha6))) ?
                          ((^~reg129) ?
                              $signed((8'hb7)) : $signed(reg682)) : $unsigned(reg831)));
                    end
                  else
                    begin
                      reg861 <= reg795[(2'h3):(1'h1)];
                      reg862 <= ({$unsigned($signed(reg733))} ?
                          $unsigned({{reg744}}) : ({reg161[(4'h8):(1'h1)]} ?
                              reg517 : reg793));
                    end
                end
              if ($unsigned(reg206))
                begin
                  for (forvar863 = (1'h0); (forvar863 < (2'h3)); forvar863 = (forvar863 + (1'h1)))
                    begin
                      reg864 <= reg766;
                      reg865 <= (~|({$signed(reg721)} >> (8'ha7)));
                      reg866 <= reg193[(3'h7):(1'h0)];
                      reg867 <= ($unsigned($unsigned(reg93[(1'h1):(1'h0)])) ^ (~(+$unsigned(reg513))));
                    end
                  reg868 <= $signed(($signed((!reg66)) ?
                      reg847[(3'h6):(2'h3)] : (reg495 <= {reg858})));
                end
              else
                begin
                  for (forvar863 = (1'h0); (forvar863 < (1'h0)); forvar863 = (forvar863 + (1'h1)))
                    begin
                      reg864 <= ($signed((~^$unsigned(reg134))) ?
                          {((reg818 ~^ reg855) ?
                                  reg124[(3'h4):(3'h4)] : $unsigned(reg143))} : (reg724[(1'h1):(1'h0)] >= ((reg788 ?
                              reg753 : reg799) != (reg569 ? reg727 : reg677))));
                      reg865 <= reg836;
                    end
                end
              for (forvar869 = (1'h0); (forvar869 < (2'h3)); forvar869 = (forvar869 + (1'h1)))
                begin
                  for (forvar870 = (1'h0); (forvar870 < (1'h0)); forvar870 = (forvar870 + (1'h1)))
                    begin
                      reg871 <= (reg149[(1'h1):(1'h1)] * forvar762);
                      reg872 <= (($unsigned($signed(reg627)) ?
                              reg151 : reg716[(2'h2):(1'h1)]) ?
                          $signed((-(-reg851))) : $signed({((8'ha9) + reg150)}));
                      reg873 <= (^~reg199);
                      reg874 <= $unsigned(((reg602 ?
                              reg132[(1'h0):(1'h0)] : reg178) ?
                          $signed((~reg660)) : (^~(reg570 >= reg194))));
                    end
                  reg875 <= $unsigned(forvar778[(3'h7):(2'h2)]);
                end
              for (forvar876 = (1'h0); (forvar876 < (1'h1)); forvar876 = (forvar876 + (1'h1)))
                begin
                  reg877 <= (!({{(8'hae)}} < (-$signed(reg560))));
                  for (forvar878 = (1'h0); (forvar878 < (2'h3)); forvar878 = (forvar878 + (1'h1)))
                    begin
                      reg879 <= (^$signed(((reg560 ?
                          reg645 : reg85) - (reg507 <= reg695))));
                      reg880 <= {(reg79 ?
                              (reg701[(3'h7):(2'h3)] ?
                                  $unsigned(forvar762) : (reg710 <= reg498)) : $unsigned((!reg706)))};
                      reg881 <= reg594[(2'h3):(2'h3)];
                      reg882 <= reg775[(4'hb):(1'h0)];
                    end
                end
            end
          reg883 <= reg194[(4'hc):(1'h0)];
          for (forvar884 = (1'h0); (forvar884 < (2'h3)); forvar884 = (forvar884 + (1'h1)))
            begin
              for (forvar885 = (1'h0); (forvar885 < (2'h3)); forvar885 = (forvar885 + (1'h1)))
                begin
                  for (forvar886 = (1'h0); (forvar886 < (1'h0)); forvar886 = (forvar886 + (1'h1)))
                    begin
                      reg887 <= {(~$unsigned($signed(reg216)))};
                      reg888 <= $signed((8'ha7));
                      reg889 <= forvar793;
                    end
                end
              if ((~(~&((reg728 || reg731) ~^ reg121))))
                begin
                  for (forvar890 = (1'h0); (forvar890 < (1'h1)); forvar890 = (forvar890 + (1'h1)))
                    begin
                      reg891 <= ((((+reg65) ?
                              $unsigned(reg853) : ((8'ha3) ~^ (8'hb2))) ^ $unsigned(reg599)) ?
                          reg92[(1'h0):(1'h0)] : reg792[(2'h3):(2'h2)]);
                    end
                end
              else
                begin
                  if ((&(|(~{reg664}))))
                    begin
                      reg890 <= $unsigned($unsigned(($unsigned(reg44) << reg509[(3'h4):(3'h4)])));
                      reg891 <= reg560;
                      reg892 <= reg151[(2'h3):(1'h1)];
                      reg893 <= reg198;
                    end
                  else
                    begin
                      reg890 <= $signed($signed(($unsigned(reg817) & (+reg790))));
                    end
                  for (forvar894 = (1'h0); (forvar894 < (2'h2)); forvar894 = (forvar894 + (1'h1)))
                    begin
                      reg895 <= (~^(^reg57[(4'hd):(4'hb)]));
                      reg896 <= (~^(~|{$signed(reg797)}));
                      reg897 <= {reg517};
                      reg898 <= forvar710;
                    end
                end
              for (forvar899 = (1'h0); (forvar899 < (2'h3)); forvar899 = (forvar899 + (1'h1)))
                begin
                  for (forvar900 = (1'h0); (forvar900 < (1'h0)); forvar900 = (forvar900 + (1'h1)))
                    begin
                      reg901 <= $unsigned((&$signed($unsigned((8'h9c)))));
                      reg902 <= ($signed((^~$signed(reg557))) ?
                          $signed($signed((|(8'ha6)))) : $unsigned(($unsigned(reg678) <<< reg14[(4'hb):(2'h2)])));
                      reg903 <= reg111[(3'h6):(1'h1)];
                    end
                end
              for (forvar904 = (1'h0); (forvar904 < (2'h2)); forvar904 = (forvar904 + (1'h1)))
                begin
                  if ($unsigned(reg64))
                    begin
                      reg905 <= ($unsigned($unsigned((~^reg169))) > (reg694 << reg647));
                      reg906 <= $signed((((reg677 > reg806) >= $signed(reg519)) | reg688));
                      reg907 <= reg557[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg905 <= forvar819[(4'h9):(3'h5)];
                      reg906 <= ({(8'hac)} & $signed((+$signed((8'ha0)))));
                    end
                  if ((+$signed({$unsigned(reg594)})))
                    begin
                      reg908 <= reg759;
                    end
                  else
                    begin
                      reg908 <= reg859[(4'he):(4'hd)];
                    end
                end
            end
        end
      for (forvar909 = (1'h0); (forvar909 < (1'h0)); forvar909 = (forvar909 + (1'h1)))
        begin
          for (forvar910 = (1'h0); (forvar910 < (2'h2)); forvar910 = (forvar910 + (1'h1)))
            begin
              if (($signed(reg112) || reg220))
                begin
                  for (forvar911 = (1'h0); (forvar911 < (2'h2)); forvar911 = (forvar911 + (1'h1)))
                    begin
                      reg912 <= (reg598[(1'h1):(1'h1)] & ((reg738 ?
                          reg725[(3'h7):(1'h1)] : reg44) || (!(~|reg889))));
                      reg913 <= (reg726[(1'h1):(1'h1)] == ((|$signed(reg97)) ?
                          (^~reg838[(4'hc):(4'hb)]) : reg726[(3'h5):(3'h5)]));
                    end
                  for (forvar914 = (1'h0); (forvar914 < (1'h1)); forvar914 = (forvar914 + (1'h1)))
                    begin
                      reg915 <= reg198[(2'h3):(1'h0)];
                      reg916 <= {$unsigned((forvar784[(4'hb):(3'h5)] > reg901[(2'h2):(2'h2)]))};
                      reg917 <= reg577;
                    end
                  if ({reg115[(2'h2):(1'h1)]})
                    begin
                      reg918 <= (~|($signed($signed(reg117)) & (forvar730 ?
                          ((8'hb3) ? reg200 : reg568) : reg770)));
                      reg919 <= (~&(reg617[(3'h4):(1'h0)] ?
                          ((reg824 < reg570) ?
                              reg498[(1'h1):(1'h1)] : (reg855 ~^ reg163)) : (reg806[(4'h8):(2'h3)] ?
                              $signed(reg139) : $signed(reg791))));
                      reg920 <= $signed(reg642);
                      reg921 <= $unsigned({$unsigned($signed(reg861))});
                    end
                  else
                    begin
                      reg918 <= $unsigned(reg79[(1'h1):(1'h0)]);
                      reg919 <= $signed({reg845});
                    end
                  if ((&($unsigned($signed(reg653)) ?
                      $signed($unsigned(reg684)) : $unsigned((reg804 ?
                          forvar724 : reg709)))))
                    begin
                      reg922 <= (+(&(reg744 - (reg792 ? reg555 : reg123))));
                      reg923 <= {reg494[(1'h0):(1'h0)]};
                      reg924 <= $signed(({$signed(reg149)} ^ ((reg804 ?
                              reg661 : (8'ha9)) ?
                          (reg204 == reg606) : (reg212 > (8'h9d)))));
                      reg925 <= $signed((((reg187 ? reg644 : reg668) ?
                              reg506[(3'h6):(2'h2)] : $signed(reg88)) ?
                          ($signed((8'ha4)) ^~ $signed(reg59)) : (8'ha1)));
                    end
                  else
                    begin
                      reg922 <= reg23;
                      reg923 <= ($signed(({reg734} < (forvar743 + reg792))) ?
                          reg26 : $signed($unsigned(((8'h9f) ?
                              forvar786 : reg690))));
                    end
                end
              else
                begin
                  for (forvar911 = (1'h0); (forvar911 < (1'h0)); forvar911 = (forvar911 + (1'h1)))
                    begin
                      reg912 <= $signed(reg852);
                      reg913 <= $unsigned(reg146[(3'h5):(1'h1)]);
                    end
                  for (forvar914 = (1'h0); (forvar914 < (1'h0)); forvar914 = (forvar914 + (1'h1)))
                    begin
                      reg915 <= (^~$unsigned(((reg868 <= reg764) >= $unsigned((8'hb5)))));
                      reg916 <= wire8[(2'h2):(1'h0)];
                    end
                end
              if (reg552)
                begin
                  if (forvar722[(4'hc):(4'ha)])
                    begin
                      reg926 <= (reg766 ?
                          ({{reg168}} ^~ reg50) : $unsigned((reg173 ^ (reg763 > (8'hb2)))));
                      reg927 <= ((forvar762 | reg170[(1'h1):(1'h0)]) & $signed({(^(8'h9d))}));
                      reg928 <= (!(+(reg906 | (~&reg881))));
                      reg929 <= ($signed(reg504) << reg871[(4'hc):(4'h9)]);
                    end
                  else
                    begin
                      reg926 <= $unsigned($signed(reg143));
                    end
                end
              else
                begin
                  if (reg666[(2'h2):(1'h0)])
                    begin
                      reg926 <= reg142[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg926 <= $signed(reg220);
                      reg927 <= reg805[(2'h3):(2'h2)];
                      reg928 <= $signed($unsigned(forvar885[(2'h3):(2'h2)]));
                      reg929 <= reg902[(2'h2):(1'h1)];
                    end
                end
              if ((~($unsigned((reg126 == reg834)) > ($signed(reg664) ~^ (&reg57)))))
                begin
                  for (forvar930 = (1'h0); (forvar930 < (1'h1)); forvar930 = (forvar930 + (1'h1)))
                    begin
                      reg931 <= (($unsigned((reg742 - reg713)) ?
                          {(^forvar785)} : ($signed(reg821) | reg705)) < $signed($signed((~reg144))));
                    end
                  for (forvar932 = (1'h0); (forvar932 < (2'h2)); forvar932 = (forvar932 + (1'h1)))
                    begin
                      reg933 <= reg537;
                      reg934 <= $unsigned((^reg565[(4'h8):(2'h3)]));
                      reg935 <= {(8'ha0)};
                    end
                  for (forvar936 = (1'h0); (forvar936 < (1'h0)); forvar936 = (forvar936 + (1'h1)))
                    begin
                      reg937 <= ((((reg160 ?
                              forvar900 : reg516) <<< $unsigned(reg797)) == ({(8'hb6)} * (reg770 ?
                              reg30 : (8'ha7)))) ?
                          ({(reg747 ? reg168 : reg557)} > ((+reg751) ?
                              $unsigned(forvar914) : reg892)) : $signed($unsigned((^reg922))));
                      reg938 <= (|reg221);
                      reg939 <= $unsigned((^reg811[(3'h4):(1'h0)]));
                      reg940 <= reg85[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  if ($unsigned(reg52[(1'h1):(1'h0)]))
                    begin
                      reg930 <= $unsigned(((^(reg213 >> reg714)) ^~ (&(forvar819 ?
                          (8'hba) : forvar732))));
                      reg931 <= ((~reg214[(1'h0):(1'h0)]) ?
                          (reg892[(4'ha):(4'ha)] ?
                              ((8'ha4) ?
                                  (reg854 ? reg219 : reg105) : (reg189 ?
                                      reg207 : reg218)) : reg89) : $signed($signed(((8'hab) ^ reg713))));
                    end
                  else
                    begin
                      reg930 <= ({$signed((reg551 ?
                              reg669 : reg215))} || {forvar736[(4'h8):(3'h4)]});
                    end
                  if (reg523[(3'h6):(1'h1)])
                    begin
                      reg932 <= (~&$signed((^~reg149)));
                      reg933 <= (~&(($signed(reg617) | (wire707 & reg841)) > $signed((reg798 * (8'ha7)))));
                      reg934 <= $signed($unsigned(((reg127 ?
                          reg139 : (8'ha2)) > (forvar825 + wire492))));
                      reg935 <= $signed(forvar710);
                    end
                  else
                    begin
                      reg932 <= $signed(reg915);
                      reg933 <= (|(-(~|(-forvar851))));
                      reg934 <= (&(!(!$unsigned(reg888))));
                    end
                end
              for (forvar941 = (1'h0); (forvar941 < (2'h2)); forvar941 = (forvar941 + (1'h1)))
                begin
                  reg942 <= (~^reg543);
                  if (reg525[(3'h6):(1'h0)])
                    begin
                      reg943 <= (($unsigned((reg675 >> forvar792)) ?
                              forvar792 : forvar769) ?
                          $unsigned(($unsigned(reg77) ^ (reg774 ?
                              reg188 : (8'had)))) : ($signed((reg211 + reg515)) >= ((^reg505) < $signed(reg759))));
                    end
                  else
                    begin
                      reg943 <= reg599;
                    end
                  for (forvar944 = (1'h0); (forvar944 < (1'h0)); forvar944 = (forvar944 + (1'h1)))
                    begin
                      reg945 <= ({forvar890} != $unsigned($signed($unsigned(reg710))));
                      reg946 <= $signed(($signed({forvar848}) ?
                          reg206 : $unsigned((reg155 ? reg645 : (8'haa)))));
                      reg947 <= (&(($signed(reg817) || (reg208 ?
                              reg117 : reg119)) ?
                          {(reg208 > reg874)} : reg525));
                    end
                  for (forvar948 = (1'h0); (forvar948 < (2'h3)); forvar948 = (forvar948 + (1'h1)))
                    begin
                      reg949 <= reg880[(1'h1):(1'h0)];
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar950 = (1'h0); (forvar950 < (2'h2)); forvar950 = (forvar950 + (1'h1)))
        begin
          for (forvar951 = (1'h0); (forvar951 < (2'h3)); forvar951 = (forvar951 + (1'h1)))
            begin
              reg952 <= $signed({((|(8'h9f)) ? (reg200 << (8'hb5)) : reg622)});
              reg953 <= reg739[(2'h2):(1'h1)];
              for (forvar954 = (1'h0); (forvar954 < (1'h0)); forvar954 = (forvar954 + (1'h1)))
                begin
                  for (forvar955 = (1'h0); (forvar955 < (2'h2)); forvar955 = (forvar955 + (1'h1)))
                    begin
                      reg956 <= reg795[(1'h1):(1'h0)];
                    end
                  for (forvar957 = (1'h0); (forvar957 < (2'h3)); forvar957 = (forvar957 + (1'h1)))
                    begin
                      reg958 <= $unsigned(($unsigned($unsigned(reg639)) & reg709[(1'h1):(1'h0)]));
                    end
                  if ((reg849[(1'h0):(1'h0)] <= reg105[(1'h0):(1'h0)]))
                    begin
                      reg959 <= (^reg880);
                      reg960 <= (~^$unsigned($unsigned((reg644 ?
                          reg614 : reg785))));
                      reg961 <= $unsigned(($unsigned((reg10 < (8'hb7))) ^ reg693[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg959 <= reg112[(1'h0):(1'h0)];
                      reg960 <= $signed($signed((reg51 ?
                          (reg168 - reg82) : reg554[(3'h5):(3'h5)])));
                    end
                end
            end
        end
      reg962 <= ((($signed(reg150) > forvar950[(4'hb):(4'h8)]) ?
          $signed(reg512) : $unsigned($signed(reg947))) - reg688[(3'h4):(1'h1)]);
      reg963 <= reg524[(3'h4):(3'h4)];
    end
  assign wire964 = reg877[(2'h3):(1'h0)];
  always
    @(posedge clk) begin
      if ((+((~|(reg115 << reg40)) ? (8'ha4) : reg805[(4'ha):(2'h2)])))
        begin
          if (reg193)
            begin
              if ($unsigned(reg766[(3'h4):(1'h1)]))
                begin
                  reg965 <= reg608[(3'h4):(1'h0)];
                  if ((($signed((!reg664)) * (((8'hae) ^ reg765) ?
                      reg89[(3'h5):(1'h0)] : (reg209 ?
                          wire492 : reg829))) || ($unsigned({reg627}) ?
                      {$signed(reg586)} : reg505[(3'h5):(3'h4)])))
                    begin
                      reg966 <= $unsigned(((^(~^reg906)) ?
                          {$signed(reg756)} : (reg714 << (reg675 ?
                              reg78 : (8'ha1)))));
                      reg967 <= ({({reg834} ?
                              $unsigned(reg822) : (^reg913))} < (8'haf));
                      reg968 <= reg804;
                    end
                  else
                    begin
                      reg966 <= (!reg595);
                    end
                  for (forvar969 = (1'h0); (forvar969 < (1'h0)); forvar969 = (forvar969 + (1'h1)))
                    begin
                      reg970 <= (reg222[(4'ha):(4'ha)] <= $signed(reg588[(4'h9):(3'h7)]));
                      reg971 <= reg718;
                      reg972 <= (reg817 + reg545);
                      reg973 <= $signed($unsigned((~^(~&reg760))));
                    end
                  for (forvar974 = (1'h0); (forvar974 < (2'h2)); forvar974 = (forvar974 + (1'h1)))
                    begin
                      reg975 <= (reg89 ?
                          reg630[(4'h8):(3'h6)] : $signed(reg811));
                      reg976 <= {reg538};
                      reg977 <= {reg220[(3'h7):(3'h7)]};
                      reg978 <= (!reg207[(2'h2):(1'h1)]);
                    end
                end
              else
                begin
                  if (reg666)
                    begin
                      reg965 <= $signed({(+(reg615 ? reg874 : (8'ha8)))});
                      reg966 <= $unsigned($unsigned(((reg630 ?
                          reg892 : (8'h9d)) < ((8'hb1) >> reg873))));
                      reg967 <= ($signed({reg711[(4'h8):(1'h0)]}) ?
                          {(+(reg853 ? reg180 : (8'hb7)))} : $signed(reg66));
                    end
                  else
                    begin
                      reg965 <= (($signed($signed(reg718)) ?
                          ((8'ha4) && (reg675 <= reg513)) : ($signed((8'ha9)) ?
                              {reg191} : ((8'ha7) <<< reg709))) >> reg109[(3'h5):(3'h4)]);
                      reg966 <= reg50;
                      reg967 <= (reg169[(1'h1):(1'h1)] ?
                          (((reg26 <<< (8'hb4)) || $unsigned(reg80)) ?
                              reg775[(2'h3):(2'h2)] : ((8'hb6) - $signed(reg515))) : (|(reg221 | $signed(reg140))));
                      reg968 <= reg101;
                    end
                  reg969 <= reg603[(3'h6):(3'h5)];
                  if (reg694[(3'h4):(1'h0)])
                    begin
                      reg970 <= (reg509[(3'h5):(1'h0)] & reg725);
                      reg971 <= $signed($signed((reg644 ?
                          {(8'hab)} : (reg630 << reg503))));
                    end
                  else
                    begin
                      reg970 <= ({{$signed(reg210)}} ?
                          reg720[(3'h4):(1'h1)] : reg563[(1'h1):(1'h1)]);
                      reg971 <= (|((+$unsigned(reg125)) <<< reg728));
                      reg972 <= (reg112 ~^ (~|($signed(reg73) ^~ $signed(reg698))));
                    end
                end
              for (forvar979 = (1'h0); (forvar979 < (1'h0)); forvar979 = (forvar979 + (1'h1)))
                begin
                  reg980 <= ($signed((^(reg40 > reg636))) ?
                      (reg535[(1'h0):(1'h0)] <<< reg47) : (8'ha6));
                  for (forvar981 = (1'h0); (forvar981 < (2'h3)); forvar981 = (forvar981 + (1'h1)))
                    begin
                      reg982 <= {(~&(+reg834))};
                      reg983 <= reg742[(2'h3):(2'h3)];
                      reg984 <= reg769[(4'h9):(1'h0)];
                      reg985 <= reg36[(2'h2):(1'h1)];
                    end
                  for (forvar986 = (1'h0); (forvar986 < (1'h1)); forvar986 = (forvar986 + (1'h1)))
                    begin
                      reg987 <= (reg156 ?
                          reg782 : $signed((+(reg796 ? reg507 : reg43))));
                      reg988 <= reg804[(1'h0):(1'h0)];
                      reg989 <= reg517;
                    end
                end
              reg990 <= reg591;
            end
          else
            begin
              for (forvar965 = (1'h0); (forvar965 < (1'h0)); forvar965 = (forvar965 + (1'h1)))
                begin
                  if (reg140)
                    begin
                      reg966 <= (((((8'had) ?
                              reg646 : wire708) <<< (reg48 & reg148)) ?
                          (8'ha3) : reg889[(4'hb):(3'h5)]) == (8'hb6));
                      reg967 <= (&reg222[(1'h1):(1'h0)]);
                      reg968 <= ((reg956[(4'he):(1'h0)] + (!(reg871 >> (8'ha7)))) ?
                          ($unsigned($signed(reg990)) ?
                              ((reg152 ? reg108 : (8'haf)) ?
                                  (~|reg789) : $signed((8'ha2))) : reg19[(3'h5):(3'h4)]) : reg780);
                    end
                  else
                    begin
                      reg966 <= (-reg943);
                      reg967 <= ({$signed({reg508})} ?
                          $unsigned(reg22[(2'h3):(2'h3)]) : $signed(((reg654 != reg541) * $unsigned(reg581))));
                      reg968 <= $unsigned($unsigned(reg563));
                      reg969 <= (8'ha5);
                    end
                  reg970 <= $unsigned(reg724);
                  if ((+$signed(((!reg45) * $signed(reg942)))))
                    begin
                      reg971 <= ({(~^((8'hb1) ?
                              (8'hba) : reg857))} || (reg647 | reg45));
                    end
                  else
                    begin
                      reg971 <= $signed(({(~|reg532)} ?
                          $unsigned(reg127[(1'h0):(1'h0)]) : ($signed(reg871) * $unsigned(reg616))));
                      reg972 <= $signed(reg663[(1'h1):(1'h0)]);
                      reg973 <= $unsigned($unsigned(reg984[(2'h3):(1'h1)]));
                      reg974 <= reg14[(3'h6):(1'h1)];
                    end
                end
              for (forvar975 = (1'h0); (forvar975 < (2'h3)); forvar975 = (forvar975 + (1'h1)))
                begin
                  reg976 <= {reg523};
                  reg977 <= $signed((+(((8'haf) ? reg110 : reg973) >>> (reg660 ?
                      reg737 : reg191))));
                  reg978 <= $signed($unsigned((^reg892)));
                  for (forvar979 = (1'h0); (forvar979 < (1'h0)); forvar979 = (forvar979 + (1'h1)))
                    begin
                      reg980 <= ($signed($unsigned(((8'hb3) > wire6))) >= $signed($unsigned({(8'hba)})));
                    end
                end
              reg981 <= (reg89[(3'h6):(2'h3)] ?
                  $unsigned(((^reg769) ?
                      (reg978 ?
                          reg47 : (8'h9f)) : $unsigned((8'h9f)))) : ({$unsigned(reg664)} | $unsigned(reg121)));
            end
        end
      else
        begin
          if (reg857[(2'h3):(2'h2)])
            begin
              if ({$unsigned(reg192)})
                begin
                  for (forvar965 = (1'h0); (forvar965 < (1'h1)); forvar965 = (forvar965 + (1'h1)))
                    begin
                      reg966 <= reg559;
                      reg967 <= (~^(~{reg503}));
                      reg968 <= ($unsigned({{(8'haa)}}) >>> reg145);
                      reg969 <= {{$signed($unsigned(reg713))}};
                    end
                  if (reg528)
                    begin
                      reg970 <= (!reg716);
                      reg971 <= reg701;
                      reg972 <= (-$signed(reg68));
                      reg973 <= (reg749[(1'h0):(1'h0)] ?
                          (((reg100 || reg205) ? reg499 : $signed(reg775)) ?
                              $unsigned((8'ha8)) : reg77[(4'h9):(2'h3)]) : reg761);
                    end
                  else
                    begin
                      reg970 <= $unsigned((+$signed(reg862)));
                      reg971 <= reg130;
                      reg972 <= ((8'hb3) ?
                          (($signed(reg888) ~^ $unsigned(reg105)) != ({reg859} ?
                              (reg855 | reg586) : reg578)) : (reg540 ?
                              ($unsigned(reg188) ?
                                  reg915 : (8'h9c)) : (~&(reg699 ?
                                  reg167 : (8'ha5)))));
                      reg973 <= $unsigned($unsigned((~^reg132)));
                    end
                  reg974 <= {$signed($signed($unsigned(reg875)))};
                  if ($signed(((~((8'ha1) > reg983)) ? reg160 : (8'ha4))))
                    begin
                      reg975 <= ($unsigned({(reg576 << (8'hab))}) ?
                          (~&reg47[(2'h2):(2'h2)]) : (reg701[(4'ha):(1'h0)] >= ({reg531} ?
                              $signed(reg175) : (reg946 != reg739))));
                      reg976 <= (-($unsigned(reg105) ?
                          (((8'hac) >> reg527) ?
                              (reg895 ^~ reg198) : (reg857 ?
                                  reg642 : reg45)) : reg599));
                      reg977 <= reg987[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg975 <= (~|(~&(~(!reg195))));
                    end
                end
              else
                begin
                  if ({($unsigned((reg199 ? reg772 : reg75)) != reg621)})
                    begin
                      reg965 <= $signed({(~(reg552 ? reg195 : reg726))});
                      reg966 <= reg763;
                    end
                  else
                    begin
                      reg965 <= ($signed(reg720[(3'h4):(2'h2)]) <<< $unsigned($unsigned(((8'haa) ?
                          reg795 : (8'hb3)))));
                      reg966 <= reg666;
                      reg967 <= ($unsigned(((reg629 ? reg796 : reg54) ?
                          reg536[(1'h1):(1'h1)] : reg963)) >> reg164);
                    end
                  reg968 <= reg605;
                  if (((reg517[(1'h1):(1'h1)] ?
                          $signed(reg64[(1'h1):(1'h0)]) : $signed((reg525 ?
                              reg598 : reg653))) ?
                      $signed($unsigned(reg37)) : $signed($unsigned($unsigned(wire8)))))
                    begin
                      reg969 <= reg671[(3'h6):(3'h6)];
                      reg970 <= (~&(-(^(reg166 & reg156))));
                      reg971 <= ($unsigned($unsigned(reg596)) | reg18);
                      reg972 <= (reg612 ? reg759[(2'h2):(1'h0)] : reg702);
                    end
                  else
                    begin
                      reg969 <= $signed((((8'hb4) ?
                          reg160 : reg110) ^ (((8'hb7) == reg657) << (&reg522))));
                      reg970 <= {$signed({(~^reg201)})};
                      reg971 <= $unsigned(reg773);
                      reg972 <= reg600;
                    end
                  for (forvar973 = (1'h0); (forvar973 < (1'h1)); forvar973 = (forvar973 + (1'h1)))
                    begin
                      reg974 <= (-reg591[(1'h0):(1'h0)]);
                      reg975 <= reg834;
                      reg976 <= $signed(reg790);
                    end
                end
            end
          else
            begin
              reg965 <= reg875;
              for (forvar966 = (1'h0); (forvar966 < (2'h3)); forvar966 = (forvar966 + (1'h1)))
                begin
                  reg967 <= ($signed(((forvar969 >= reg926) < (&reg581))) << (^~(^(reg893 << reg198))));
                  for (forvar968 = (1'h0); (forvar968 < (2'h2)); forvar968 = (forvar968 + (1'h1)))
                    begin
                      reg969 <= (wire8[(2'h2):(1'h0)] ?
                          {{$signed(reg168)}} : reg852);
                      reg970 <= {((~^(reg673 ? reg540 : reg165)) ?
                              $unsigned((^~reg788)) : (!$signed(reg215)))};
                      reg971 <= $unsigned((8'hae));
                    end
                end
            end
          if ((reg195 ?
              (!($unsigned(reg545) ^ reg922)) : (((reg109 ? reg543 : (8'ha4)) ?
                  (reg186 ^ reg690) : (^~reg678)) ^ $unsigned($unsigned(reg654)))))
            begin
              for (forvar978 = (1'h0); (forvar978 < (1'h1)); forvar978 = (forvar978 + (1'h1)))
                begin
                  for (forvar979 = (1'h0); (forvar979 < (1'h1)); forvar979 = (forvar979 + (1'h1)))
                    begin
                      reg980 <= (reg652 && reg150[(2'h2):(2'h2)]);
                    end
                end
              for (forvar981 = (1'h0); (forvar981 < (2'h3)); forvar981 = (forvar981 + (1'h1)))
                begin
                  for (forvar982 = (1'h0); (forvar982 < (2'h2)); forvar982 = (forvar982 + (1'h1)))
                    begin
                      reg983 <= (+($unsigned($signed(reg775)) ?
                          (8'haf) : reg194[(2'h2):(1'h1)]));
                      reg984 <= ((reg907[(2'h2):(2'h2)] ^~ (~(reg953 && reg496))) - reg95);
                      reg985 <= $signed($signed($unsigned((reg929 >> reg616))));
                    end
                end
              reg986 <= (((+$signed(reg760)) ?
                  (8'ha1) : reg22[(1'h0):(1'h0)]) > reg687);
              reg987 <= $unsigned((reg858 ?
                  ($signed(reg110) * reg502[(2'h2):(1'h0)]) : $signed(reg586)));
            end
          else
            begin
              if ({reg727[(2'h2):(1'h0)]})
                begin
                  reg978 <= reg223;
                end
              else
                begin
                  if (($signed({$unsigned(reg187)}) ?
                      {$signed($unsigned(reg925))} : $signed(reg145[(1'h1):(1'h1)])))
                    begin
                      reg978 <= (^~($signed((reg824 ? reg207 : (8'had))) ?
                          $unsigned(((8'ha1) > reg547)) : {$signed(reg930)}));
                    end
                  else
                    begin
                      reg978 <= (reg152 < $unsigned($unsigned($unsigned(reg556))));
                      reg979 <= {($unsigned($signed((8'ha8))) ^ $unsigned(reg98[(2'h3):(2'h3)]))};
                      reg980 <= $unsigned((^reg523[(4'hb):(4'h8)]));
                      reg981 <= ($signed(((forvar978 ? reg581 : reg932) ?
                          (-reg109) : reg849[(1'h0):(1'h0)])) > reg915);
                    end
                  for (forvar982 = (1'h0); (forvar982 < (1'h1)); forvar982 = (forvar982 + (1'h1)))
                    begin
                      reg983 <= reg184[(3'h7):(3'h5)];
                      reg984 <= {$signed(reg745[(1'h0):(1'h0)])};
                      reg985 <= (~&(((reg156 != reg749) & $signed(reg540)) ?
                          reg927 : reg800[(3'h4):(3'h4)]));
                    end
                  if ({($unsigned($signed(reg867)) ?
                          {(reg962 ? (8'ha3) : reg657)} : $signed((~reg768)))})
                    begin
                      reg986 <= wire707[(3'h4):(1'h0)];
                      reg987 <= $unsigned(reg114);
                      reg988 <= {reg747[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg986 <= (8'ha2);
                      reg987 <= ((+(8'ha1)) ?
                          {((^reg657) || $signed(reg981))} : {reg755});
                      reg988 <= reg650;
                      reg989 <= $unsigned($signed($signed($unsigned(reg590))));
                    end
                  if ($signed((reg971 ?
                      reg693[(2'h3):(1'h0)] : (~reg930[(3'h5):(1'h1)]))))
                    begin
                      reg990 <= ({(8'hb8)} >>> ($signed($unsigned(reg819)) ?
                          (-reg919[(1'h1):(1'h1)]) : $unsigned((forvar969 | reg791))));
                      reg991 <= ($unsigned((reg498 ?
                              $unsigned((8'hb7)) : reg567[(2'h2):(2'h2)])) ?
                          (!{(^~reg818)}) : (^reg850[(2'h2):(1'h1)]));
                      reg992 <= {($signed((reg680 ?
                              (8'h9d) : reg84)) || $unsigned($signed(reg626)))};
                    end
                  else
                    begin
                      reg990 <= {reg502};
                      reg991 <= (!(8'ha1));
                    end
                end
              if ($unsigned($unsigned($signed(wire492[(4'hd):(4'h9)]))))
                begin
                  for (forvar993 = (1'h0); (forvar993 < (2'h3)); forvar993 = (forvar993 + (1'h1)))
                    begin
                      reg994 <= (reg898[(4'hd):(4'ha)] ?
                          (reg122 <= $unsigned((+reg800))) : (~|reg665));
                      reg995 <= (({$signed(reg529)} & reg633[(4'h8):(4'h8)]) ?
                          $unsigned({(~^reg875)}) : reg596);
                    end
                  for (forvar996 = (1'h0); (forvar996 < (1'h0)); forvar996 = (forvar996 + (1'h1)))
                    begin
                      reg997 <= (8'hb2);
                      reg998 <= reg853;
                      reg999 <= $unsigned((reg204 ?
                          $unsigned(reg763[(4'h9):(2'h3)]) : $signed((~^(8'haa)))));
                      reg1000 <= $unsigned($unsigned(reg790[(4'h9):(3'h7)]));
                    end
                  if (($unsigned(reg116[(3'h6):(1'h1)]) ?
                      (~^$unsigned($signed(reg895))) : reg637))
                    begin
                      reg1001 <= $unsigned(((reg784[(3'h5):(3'h4)] ?
                              $unsigned(reg813) : $signed(reg586)) ?
                          reg109[(1'h0):(1'h0)] : $signed(reg931)));
                      reg1002 <= $unsigned((reg842[(4'he):(2'h2)] & ($signed(reg157) + reg664[(2'h3):(1'h0)])));
                      reg1003 <= reg519;
                      reg1004 <= ($signed($signed((!reg746))) ?
                          $signed({{reg121}}) : reg913[(3'h7):(2'h2)]);
                    end
                  else
                    begin
                      reg1001 <= $unsigned($signed((reg637[(3'h7):(3'h4)] <<< $signed(reg16))));
                      reg1002 <= reg976;
                    end
                end
              else
                begin
                  reg993 <= ((8'hb7) ? (~^{$unsigned(reg39)}) : {reg145});
                  reg994 <= (~^($signed((+forvar965)) ?
                      $signed($signed(forvar966)) : (((8'hba) ?
                              reg570 : reg650) ?
                          $unsigned((8'h9d)) : $unsigned(reg135))));
                end
            end
          for (forvar1005 = (1'h0); (forvar1005 < (1'h0)); forvar1005 = (forvar1005 + (1'h1)))
            begin
              if (((reg737 ?
                      $unsigned($unsigned(reg200)) : ($unsigned(reg989) ?
                          reg81 : ((8'hb8) ^ (8'h9d)))) ?
                  reg836[(4'hf):(4'h8)] : reg835[(2'h2):(2'h2)]))
                begin
                  for (forvar1006 = (1'h0); (forvar1006 < (2'h2)); forvar1006 = (forvar1006 + (1'h1)))
                    begin
                      reg1007 <= ($unsigned(reg98) >> (8'ha1));
                      reg1008 <= (reg82[(3'h6):(1'h1)] ?
                          (~|reg207) : $unsigned((-((8'ha0) ?
                              reg675 : reg1000))));
                      reg1009 <= $signed(reg774);
                      reg1010 <= reg134[(3'h5):(1'h0)];
                    end
                  for (forvar1011 = (1'h0); (forvar1011 < (2'h3)); forvar1011 = (forvar1011 + (1'h1)))
                    begin
                      reg1012 <= $unsigned($unsigned($unsigned((reg190 ?
                          reg659 : reg834))));
                      reg1013 <= reg780;
                    end
                  for (forvar1014 = (1'h0); (forvar1014 < (2'h2)); forvar1014 = (forvar1014 + (1'h1)))
                    begin
                      reg1015 <= ({((reg674 ? (8'hb2) : reg36) >> ((8'hb8) ?
                                  reg82 : reg712))} ?
                          {reg542[(1'h0):(1'h0)]} : reg805[(3'h7):(1'h0)]);
                    end
                  reg1016 <= $signed(reg512);
                end
              else
                begin
                  for (forvar1006 = (1'h0); (forvar1006 < (1'h1)); forvar1006 = (forvar1006 + (1'h1)))
                    begin
                      reg1007 <= (^~$unsigned(reg80));
                      reg1008 <= ($unsigned((!$unsigned(reg839))) >= $signed($unsigned($signed(reg636))));
                    end
                  for (forvar1009 = (1'h0); (forvar1009 < (2'h3)); forvar1009 = (forvar1009 + (1'h1)))
                    begin
                      reg1010 <= forvar973;
                    end
                  reg1011 <= {{$signed((^wire9))}};
                end
              if (reg976[(3'h6):(2'h3)])
                begin
                  if ((8'ha4))
                    begin
                      reg1017 <= reg637[(4'ha):(1'h0)];
                      reg1018 <= reg719;
                      reg1019 <= (($signed($signed(reg610)) ?
                          (!{reg557}) : $signed((!(8'hba)))) * reg805);
                      reg1020 <= reg56[(4'h9):(2'h3)];
                    end
                  else
                    begin
                      reg1017 <= reg102[(2'h3):(2'h2)];
                      reg1018 <= (({reg178[(2'h2):(1'h0)]} >>> reg781) ?
                          $unsigned($signed((reg976 ?
                              reg44 : reg594))) : {forvar996[(4'hb):(4'ha)]});
                    end
                  reg1021 <= reg734[(3'h4):(1'h0)];
                end
              else
                begin
                  if ((reg681[(1'h0):(1'h0)] && reg164[(1'h1):(1'h0)]))
                    begin
                      reg1017 <= (reg34 ?
                          ({(reg985 > reg960)} ?
                              (reg570[(4'ha):(3'h5)] ?
                                  (~|reg213) : (~|reg515)) : ((reg760 ?
                                  reg879 : reg119) & $unsigned(reg679))) : {reg626[(3'h5):(3'h5)]});
                      reg1018 <= $signed(reg772[(3'h6):(2'h2)]);
                      reg1019 <= reg80[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1017 <= reg107;
                    end
                end
              if ((^(~&((reg142 ? forvar978 : reg1019) ?
                  (reg182 ? reg860 : reg210) : reg553))))
                begin
                  if ($unsigned((($signed(reg500) >> reg715) ?
                      {((8'haf) ? reg856 : reg569)} : (reg605 <<< reg568))))
                    begin
                      reg1022 <= $signed($signed($unsigned(reg928)));
                    end
                  else
                    begin
                      reg1022 <= $signed(reg1016);
                    end
                  if ((-reg758))
                    begin
                      reg1023 <= (($unsigned((reg171 == reg222)) ?
                              ((reg40 ? (8'ha1) : reg218) ?
                                  {reg222} : $unsigned(reg616)) : ((^~(8'ha6)) ?
                                  $signed(reg872) : reg512)) ?
                          {reg734[(3'h7):(1'h1)]} : reg1003[(4'h9):(1'h1)]);
                    end
                  else
                    begin
                      reg1023 <= ($unsigned(($unsigned((8'hb0)) || (reg1023 <<< reg729))) != reg719);
                      reg1024 <= $unsigned($signed(((reg686 ?
                              (8'hac) : reg731) ?
                          (8'ha5) : (reg114 < reg680))));
                      reg1025 <= (^((~^(reg592 ~^ reg121)) ?
                          (^~$unsigned((8'h9c))) : $unsigned($unsigned(reg970))));
                    end
                end
              else
                begin
                  reg1022 <= {forvar978};
                  reg1023 <= ($unsigned(((reg108 ? reg714 : reg929) > (reg22 ?
                          reg204 : reg873))) ?
                      $signed((reg103 <<< reg556)) : (~|reg497));
                  for (forvar1024 = (1'h0); (forvar1024 < (1'h1)); forvar1024 = (forvar1024 + (1'h1)))
                    begin
                      reg1025 <= (8'hb2);
                      reg1026 <= (~&($unsigned(reg673) ?
                          (|(+reg722)) : ($unsigned(reg209) <<< (reg193 + reg613))));
                      reg1027 <= (({reg599} ?
                          reg93[(2'h3):(1'h1)] : ({reg19} ?
                              {reg1018} : (^~reg905))) <= $signed(reg531[(4'ha):(3'h6)]));
                    end
                end
            end
          for (forvar1028 = (1'h0); (forvar1028 < (2'h3)); forvar1028 = (forvar1028 + (1'h1)))
            begin
              if (((^~reg680) == reg68[(2'h2):(2'h2)]))
                begin
                  reg1029 <= $unsigned((~|($signed((8'hae)) ?
                      reg592 : {reg796})));
                end
              else
                begin
                  if ({$signed(($signed((8'h9c)) ?
                          reg962 : (reg193 ? (8'ha4) : reg668)))})
                    begin
                      reg1029 <= (-$unsigned(reg692[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1029 <= $unsigned($signed((+(wire9 > reg506))));
                      reg1030 <= ((|reg984[(2'h3):(2'h3)]) ?
                          (&(reg531[(3'h6):(3'h6)] >>> (reg731 * reg119))) : ({$signed(reg713)} ^ $unsigned(reg1012[(1'h0):(1'h0)])));
                      reg1031 <= ((reg723 ?
                          reg605 : ((reg208 ? reg185 : (8'hb9)) ?
                              (reg553 ?
                                  reg671 : reg921) : $signed(reg100))) < (&reg192[(2'h2):(2'h2)]));
                    end
                end
              for (forvar1032 = (1'h0); (forvar1032 < (2'h3)); forvar1032 = (forvar1032 + (1'h1)))
                begin
                  for (forvar1033 = (1'h0); (forvar1033 < (2'h3)); forvar1033 = (forvar1033 + (1'h1)))
                    begin
                      reg1034 <= reg923[(2'h2):(1'h0)];
                      reg1035 <= (+$signed((!$signed(reg110))));
                    end
                  if ((-reg17[(4'hd):(2'h3)]))
                    begin
                      reg1036 <= (~((~$unsigned(reg39)) ?
                          ({reg501} ?
                              reg688[(1'h0):(1'h0)] : (reg768 >> reg130)) : reg641));
                      reg1037 <= ($signed({reg209}) <= $signed((8'hae)));
                    end
                  else
                    begin
                      reg1036 <= {$signed({((8'hb7) ? reg93 : (8'ha8))})};
                      reg1037 <= $unsigned(reg77);
                    end
                end
            end
        end
      for (forvar1038 = (1'h0); (forvar1038 < (2'h3)); forvar1038 = (forvar1038 + (1'h1)))
        begin
          reg1039 <= (~^reg677);
        end
    end
  assign wire1040 = reg966;
  always
    @(posedge clk) begin
      reg1041 <= (($signed((reg855 ? reg667 : reg215)) - ((reg513 & reg767) ?
          reg959[(2'h2):(2'h2)] : $signed(reg702))) ^~ (reg800 ^~ {reg710[(2'h3):(1'h0)]}));
      if ($signed($signed(reg16[(2'h3):(2'h3)])))
        begin
          for (forvar1042 = (1'h0); (forvar1042 < (2'h2)); forvar1042 = (forvar1042 + (1'h1)))
            begin
              reg1043 <= (^((~&reg152) ?
                  (-(reg898 << reg1004)) : (~|(!reg644))));
            end
          reg1044 <= ({{$signed(reg18)}} > (reg121[(4'h9):(3'h6)] ?
              ((~&reg220) ?
                  (reg712 && reg787) : $unsigned(reg653)) : reg211[(4'h9):(3'h7)]));
          for (forvar1045 = (1'h0); (forvar1045 < (2'h3)); forvar1045 = (forvar1045 + (1'h1)))
            begin
              if (reg609[(3'h6):(1'h0)])
                begin
                  for (forvar1046 = (1'h0); (forvar1046 < (2'h2)); forvar1046 = (forvar1046 + (1'h1)))
                    begin
                      reg1047 <= reg772;
                      reg1048 <= reg85[(3'h5):(3'h5)];
                      reg1049 <= reg669;
                      reg1050 <= {$unsigned(reg114[(3'h5):(2'h3)])};
                    end
                end
              else
                begin
                  if ($signed(($signed((reg686 ? reg667 : forvar1042)) ?
                      $signed($unsigned(reg835)) : (reg1000 ?
                          (-reg908) : (reg523 ? reg689 : (8'ha5))))))
                    begin
                      reg1046 <= {(reg605 ?
                              reg554[(3'h4):(2'h2)] : ({reg512} + $unsigned(reg516)))};
                      reg1047 <= (~&$signed((8'hb6)));
                      reg1048 <= ($unsigned(((reg10 >= reg110) ?
                              (reg103 ? reg1008 : reg862) : {reg840})) ?
                          (^~(!$signed((8'h9c)))) : (reg147 ?
                              (^(|reg126)) : ((reg713 ^ reg599) - (reg698 != reg942))));
                      reg1049 <= reg74[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1046 <= (&((~|(~^(8'hb9))) ?
                          reg586[(1'h1):(1'h1)] : reg142));
                      reg1047 <= reg664;
                      reg1048 <= (^~(8'ha2));
                    end
                  for (forvar1050 = (1'h0); (forvar1050 < (1'h1)); forvar1050 = (forvar1050 + (1'h1)))
                    begin
                      reg1051 <= reg591;
                      reg1052 <= reg974;
                      reg1053 <= {(($signed(reg1010) <<< {reg693}) ?
                              $signed($unsigned((8'hae))) : (8'ha4))};
                    end
                  for (forvar1054 = (1'h0); (forvar1054 < (1'h1)); forvar1054 = (forvar1054 + (1'h1)))
                    begin
                      reg1055 <= {$signed(((!reg634) > $signed(reg943)))};
                      reg1056 <= (&$signed((8'hba)));
                      reg1057 <= reg547;
                      reg1058 <= reg647[(2'h2):(1'h0)];
                    end
                  reg1059 <= ({((8'hae) ? (|reg177) : (-reg793))} ?
                      {reg671[(1'h1):(1'h1)]} : ((reg795[(2'h3):(1'h1)] ?
                              (reg1018 ? reg664 : reg203) : (reg1051 ?
                                  reg959 : reg501)) ?
                          {{reg106}} : ($signed(reg509) <= reg756)));
                end
              if (reg978[(3'h5):(1'h0)])
                begin
                  reg1060 <= (!((-$unsigned(reg706)) ?
                      ((reg935 + (8'ha6)) ?
                          ((8'haf) ?
                              wire1040 : reg124) : (reg866 | (8'hb1))) : reg157[(2'h2):(1'h0)]));
                end
              else
                begin
                  for (forvar1060 = (1'h0); (forvar1060 < (1'h0)); forvar1060 = (forvar1060 + (1'h1)))
                    begin
                      reg1061 <= reg743;
                      reg1062 <= $signed($signed(reg821));
                    end
                end
            end
        end
      else
        begin
          reg1042 <= $unsigned($signed($unsigned(reg720[(1'h1):(1'h0)])));
          for (forvar1043 = (1'h0); (forvar1043 < (2'h2)); forvar1043 = (forvar1043 + (1'h1)))
            begin
              if (((reg111[(1'h0):(1'h0)] ?
                  $signed((reg968 << reg599)) : ((reg722 ?
                      reg517 : (8'ha1)) ^~ reg167)) <= $unsigned(reg796)))
                begin
                  for (forvar1044 = (1'h0); (forvar1044 < (1'h1)); forvar1044 = (forvar1044 + (1'h1)))
                    begin
                      reg1045 <= (reg560 ?
                          reg513 : ({(reg157 ? reg958 : reg803)} ?
                              reg749 : (~|$unsigned(reg795))));
                      reg1046 <= reg1019;
                      reg1047 <= ((^reg865[(4'h8):(1'h1)]) ?
                          ($signed($signed((8'hab))) >>> (reg207[(4'hc):(3'h7)] ?
                              $unsigned(wire492) : reg714[(4'h8):(3'h4)])) : reg147[(1'h1):(1'h1)]);
                    end
                  reg1048 <= reg192;
                  if ((8'ha7))
                    begin
                      reg1049 <= reg34;
                      reg1050 <= ((-({reg1030} && $signed(reg109))) != (&reg220[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1049 <= $unsigned((+(~|reg556)));
                      reg1050 <= (reg820[(1'h1):(1'h0)] ?
                          (reg176 || (reg592[(2'h2):(2'h2)] != (!reg749))) : reg589);
                      reg1051 <= $unsigned(reg786);
                      reg1052 <= (~&reg1009[(3'h5):(1'h1)]);
                    end
                  reg1053 <= {(-($unsigned(reg901) ? {reg109} : (~&reg799)))};
                end
              else
                begin
                  for (forvar1044 = (1'h0); (forvar1044 < (2'h3)); forvar1044 = (forvar1044 + (1'h1)))
                    begin
                      reg1045 <= ($unsigned($unsigned((reg1043 ?
                          reg991 : reg194))) << reg767);
                    end
                  for (forvar1046 = (1'h0); (forvar1046 < (1'h0)); forvar1046 = (forvar1046 + (1'h1)))
                    begin
                      reg1047 <= ($signed((reg121 ?
                          $signed((8'h9d)) : $unsigned((8'ha5)))) << reg537);
                      reg1048 <= reg934[(3'h5):(3'h5)];
                      reg1049 <= $signed((^~reg1048));
                    end
                  if (reg148)
                    begin
                      reg1050 <= (-reg206[(1'h1):(1'h0)]);
                      reg1051 <= {($signed(reg560) ?
                              (-(reg42 ? (8'hb4) : reg737)) : ($signed(reg149) ?
                                  $signed(reg864) : $unsigned(reg36)))};
                      reg1052 <= reg975;
                      reg1053 <= (reg624[(2'h2):(2'h2)] && $signed(reg831));
                    end
                  else
                    begin
                      reg1050 <= reg799;
                      reg1051 <= reg516;
                      reg1052 <= (8'hb3);
                      reg1053 <= {(reg836 ?
                              $signed(reg774) : reg729[(1'h0):(1'h0)])};
                    end
                end
              for (forvar1054 = (1'h0); (forvar1054 < (2'h3)); forvar1054 = (forvar1054 + (1'h1)))
                begin
                  reg1055 <= reg184;
                end
              if (($signed(({reg723} * (reg858 ?
                  forvar1045 : reg70))) <= $unsigned($unsigned($unsigned((8'ha7))))))
                begin
                  for (forvar1056 = (1'h0); (forvar1056 < (2'h3)); forvar1056 = (forvar1056 + (1'h1)))
                    begin
                      reg1057 <= {reg847[(2'h2):(1'h1)]};
                    end
                  for (forvar1058 = (1'h0); (forvar1058 < (1'h1)); forvar1058 = (forvar1058 + (1'h1)))
                    begin
                      reg1059 <= ((($signed(reg987) * (reg88 | reg551)) >>> reg576[(3'h4):(1'h0)]) ?
                          $signed(((^~reg673) && {reg847})) : $signed($unsigned((8'ha4))));
                      reg1060 <= (8'ha3);
                      reg1061 <= (^$signed($unsigned((reg836 ?
                          reg580 : reg740))));
                    end
                end
              else
                begin
                  for (forvar1056 = (1'h0); (forvar1056 < (1'h0)); forvar1056 = (forvar1056 + (1'h1)))
                    begin
                      reg1057 <= $unsigned(($unsigned($unsigned(reg95)) ?
                          (~|reg547[(1'h1):(1'h0)]) : (~&(reg638 * reg684))));
                      reg1058 <= (^reg109);
                    end
                  reg1059 <= $signed(reg622);
                  for (forvar1060 = (1'h0); (forvar1060 < (1'h0)); forvar1060 = (forvar1060 + (1'h1)))
                    begin
                      reg1061 <= $unsigned(reg896);
                    end
                end
              reg1062 <= reg508[(3'h5):(3'h5)];
            end
          for (forvar1063 = (1'h0); (forvar1063 < (1'h0)); forvar1063 = (forvar1063 + (1'h1)))
            begin
              reg1064 <= reg183[(4'hd):(4'h8)];
            end
          reg1065 <= $signed((^(reg715 > (~&reg923))));
        end
      for (forvar1066 = (1'h0); (forvar1066 < (2'h2)); forvar1066 = (forvar1066 + (1'h1)))
        begin
          for (forvar1067 = (1'h0); (forvar1067 < (1'h0)); forvar1067 = (forvar1067 + (1'h1)))
            begin
              for (forvar1068 = (1'h0); (forvar1068 < (1'h0)); forvar1068 = (forvar1068 + (1'h1)))
                begin
                  if (reg216)
                    begin
                      reg1069 <= (~^reg95[(2'h2):(2'h2)]);
                      reg1070 <= ((reg16 * reg590) | $unsigned(reg788[(3'h4):(3'h4)]));
                      reg1071 <= wire9;
                    end
                  else
                    begin
                      reg1069 <= reg972[(4'hc):(2'h3)];
                      reg1070 <= $unsigned($signed((reg499[(2'h3):(1'h0)] ?
                          (reg968 >>> reg969) : reg992[(2'h2):(1'h1)])));
                      reg1071 <= reg946[(1'h1):(1'h0)];
                      reg1072 <= $unsigned(reg794);
                    end
                  reg1073 <= (^~(($unsigned(reg906) ?
                      $signed(reg174) : (reg905 >>> (8'h9f))) ^ reg30));
                  for (forvar1074 = (1'h0); (forvar1074 < (1'h0)); forvar1074 = (forvar1074 + (1'h1)))
                    begin
                      reg1075 <= (+$unsigned(((reg855 ?
                          reg171 : reg774) * reg41[(3'h6):(1'h0)])));
                      reg1076 <= reg678[(2'h2):(2'h2)];
                    end
                end
              for (forvar1077 = (1'h0); (forvar1077 < (2'h2)); forvar1077 = (forvar1077 + (1'h1)))
                begin
                  for (forvar1078 = (1'h0); (forvar1078 < (2'h3)); forvar1078 = (forvar1078 + (1'h1)))
                    begin
                      reg1079 <= (reg958 ?
                          (|($signed(reg45) ?
                              reg547[(2'h2):(1'h0)] : reg618[(1'h0):(1'h0)])) : {($signed(reg720) << $signed((8'ha0)))});
                      reg1080 <= $unsigned(reg921);
                      reg1081 <= ((&({reg946} <<< reg646[(3'h6):(3'h5)])) ?
                          $signed(reg745[(2'h2):(1'h0)]) : (~^reg146));
                      reg1082 <= $unsigned($unsigned((-(8'hb8))));
                    end
                  for (forvar1083 = (1'h0); (forvar1083 < (2'h2)); forvar1083 = (forvar1083 + (1'h1)))
                    begin
                      reg1084 <= ((((~|reg793) | (-reg624)) ?
                          reg956 : ($signed(reg751) ?
                              (&(8'hae)) : $signed((8'hb2)))) == {{(-reg562)}});
                      reg1085 <= ($signed((-reg918)) ? reg921 : reg126);
                    end
                  if ($signed(reg881[(1'h0):(1'h0)]))
                    begin
                      reg1086 <= reg792;
                      reg1087 <= $signed(reg1009);
                    end
                  else
                    begin
                      reg1086 <= ((forvar1043 || reg641[(4'hb):(3'h6)]) * {$signed($signed(reg949))});
                      reg1087 <= reg589[(4'hc):(3'h5)];
                      reg1088 <= reg880[(4'hc):(3'h7)];
                      reg1089 <= {(^((8'ha2) ?
                              (reg704 ? reg100 : reg149) : {(8'ha8)}))};
                    end
                end
              if (reg746)
                begin
                  for (forvar1090 = (1'h0); (forvar1090 < (1'h0)); forvar1090 = (forvar1090 + (1'h1)))
                    begin
                      reg1091 <= (^(wire492[(3'h6):(2'h3)] * $signed($unsigned(reg779))));
                      reg1092 <= (8'ha8);
                      reg1093 <= (!$unsigned($unsigned((reg804 ?
                          reg764 : reg1024))));
                      reg1094 <= (^{reg145});
                    end
                  if (reg829[(3'h5):(1'h1)])
                    begin
                      reg1095 <= ((~reg221[(2'h3):(2'h3)]) ?
                          ($unsigned($unsigned(reg660)) ?
                              reg100 : ((reg1025 ?
                                  reg13 : reg974) ^~ reg952[(2'h2):(1'h0)])) : $signed({(8'hae)}));
                    end
                  else
                    begin
                      reg1095 <= $unsigned(reg10);
                      reg1096 <= reg897;
                      reg1097 <= (-$unsigned(reg723));
                    end
                  for (forvar1098 = (1'h0); (forvar1098 < (2'h3)); forvar1098 = (forvar1098 + (1'h1)))
                    begin
                      reg1099 <= (reg548[(1'h1):(1'h1)] ?
                          $signed((|(reg881 & reg64))) : reg1044);
                    end
                end
              else
                begin
                  if ((!{reg1088[(4'hb):(4'hb)]}))
                    begin
                      reg1090 <= $signed(reg531);
                      reg1091 <= (8'ha6);
                      reg1092 <= (reg887[(2'h3):(2'h3)] ?
                          {(8'ha8)} : reg946[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1090 <= reg496[(3'h6):(1'h1)];
                      reg1091 <= $signed(reg511[(3'h6):(1'h0)]);
                      reg1092 <= ($unsigned($unsigned(((8'h9d) ?
                          reg889 : (8'ha3)))) & reg688);
                    end
                end
            end
          for (forvar1100 = (1'h0); (forvar1100 < (1'h1)); forvar1100 = (forvar1100 + (1'h1)))
            begin
              if ((~^((reg1011 ?
                  (reg33 ?
                      reg657 : reg132) : (reg796 >> reg779)) > $unsigned((|reg192)))))
                begin
                  if ($signed((^{(reg528 ? reg111 : reg784)})))
                    begin
                      reg1101 <= $unsigned({reg529});
                      reg1102 <= (({{reg595}} ?
                          (~|(8'ha5)) : {$unsigned((8'hb6))}) && $signed($signed((reg922 >>> (8'ha9)))));
                    end
                  else
                    begin
                      reg1101 <= $signed({$signed({reg75})});
                      reg1102 <= reg927;
                    end
                  if (($unsigned(reg741) >> reg548[(1'h1):(1'h1)]))
                    begin
                      reg1103 <= $unsigned(((&$signed(reg887)) ^ (+(+reg701))));
                      reg1104 <= reg111[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1103 <= {$unsigned({reg176})};
                      reg1104 <= reg1024;
                      reg1105 <= ((~^({reg32} ?
                              (reg921 > (8'hb3)) : (reg1036 ?
                                  (8'hab) : reg856))) ?
                          {(^~$unsigned(reg16))} : (reg609 && (&$unsigned(reg840))));
                      reg1106 <= reg105;
                    end
                  if (reg513)
                    begin
                      reg1107 <= reg103;
                      reg1108 <= reg26;
                    end
                  else
                    begin
                      reg1107 <= reg79[(3'h6):(3'h5)];
                      reg1108 <= reg696[(3'h5):(2'h2)];
                      reg1109 <= reg716;
                      reg1110 <= {{$unsigned($unsigned(reg1047))}};
                    end
                end
              else
                begin
                  if (reg1037)
                    begin
                      reg1101 <= $unsigned(reg729[(1'h0):(1'h0)]);
                      reg1102 <= (((&$unsigned(reg586)) != $signed(reg38[(1'h1):(1'h1)])) ?
                          ($unsigned((~|reg569)) ?
                              $unsigned(reg22) : ((!(8'had)) ?
                                  (~reg793) : (~reg927))) : reg48);
                    end
                  else
                    begin
                      reg1101 <= $signed({(~&(-reg902))});
                      reg1102 <= {reg651[(4'ha):(4'ha)]};
                    end
                  for (forvar1103 = (1'h0); (forvar1103 < (2'h2)); forvar1103 = (forvar1103 + (1'h1)))
                    begin
                      reg1104 <= (~(reg1089[(1'h1):(1'h1)] ?
                          ($unsigned((8'had)) <= reg654) : reg922));
                      reg1105 <= ($signed({reg17}) ?
                          reg163[(1'h1):(1'h0)] : ((^(reg1012 ?
                              reg513 : (8'haa))) ~^ ($unsigned(reg674) ?
                              $unsigned(reg670) : $signed(reg661))));
                      reg1106 <= $signed((reg862 ?
                          reg732[(1'h1):(1'h1)] : $signed($signed((8'ha2)))));
                    end
                  if ((8'hb7))
                    begin
                      reg1107 <= {(^~reg1106[(3'h5):(1'h0)])};
                    end
                  else
                    begin
                      reg1107 <= ((~|reg773) ?
                          {(^~(forvar1056 >= reg770))} : (reg637[(2'h3):(1'h0)] ?
                              (~^reg834[(2'h3):(1'h0)]) : ((~&reg643) ?
                                  (reg806 ?
                                      reg100 : reg622) : reg789[(2'h2):(1'h0)])));
                      reg1108 <= (reg930[(4'hd):(4'h8)] ?
                          reg588[(4'h8):(1'h1)] : (~&$unsigned($unsigned((8'ha6)))));
                      reg1109 <= (~$unsigned((^$unsigned(reg155))));
                    end
                  for (forvar1110 = (1'h0); (forvar1110 < (1'h1)); forvar1110 = (forvar1110 + (1'h1)))
                    begin
                      reg1111 <= reg76;
                      reg1112 <= reg704[(2'h2):(1'h0)];
                    end
                end
              if (reg599)
                begin
                  for (forvar1113 = (1'h0); (forvar1113 < (2'h2)); forvar1113 = (forvar1113 + (1'h1)))
                    begin
                      reg1114 <= ((reg684 | $signed(reg539)) | reg1087[(4'ha):(3'h5)]);
                      reg1115 <= ((~|{(reg816 ? (8'hb5) : reg940)}) ?
                          (&$signed($unsigned(reg967))) : (~$unsigned((^~(8'hac)))));
                    end
                end
              else
                begin
                  if (reg204[(3'h6):(3'h5)])
                    begin
                      reg1113 <= (reg592[(3'h5):(2'h2)] ?
                          (+reg156) : (~^{(reg523 | reg806)}));
                      reg1114 <= ((~^(reg1079[(3'h4):(1'h0)] + (~reg754))) || ((~&((8'hba) - reg783)) + ((~|reg785) <= (reg190 != reg952))));
                      reg1115 <= reg835[(2'h2):(1'h0)];
                      reg1116 <= $unsigned(reg781);
                    end
                  else
                    begin
                      reg1113 <= reg987;
                      reg1114 <= ($unsigned({(reg728 ^ reg857)}) == $unsigned($unsigned($signed(reg580))));
                      reg1115 <= ($signed(reg689[(3'h5):(1'h0)]) - reg925[(2'h2):(1'h1)]);
                    end
                  for (forvar1117 = (1'h0); (forvar1117 < (1'h0)); forvar1117 = (forvar1117 + (1'h1)))
                    begin
                      reg1118 <= reg1099[(2'h3):(2'h2)];
                      reg1119 <= $signed($signed((~|$unsigned(reg834))));
                      reg1120 <= ($unsigned((~reg767[(2'h3):(1'h1)])) ?
                          ({{(8'hb2)}} > reg509[(3'h4):(1'h0)]) : (&(((8'ha2) || reg665) && ((8'h9e) != reg743))));
                    end
                end
              if (reg1064)
                begin
                  for (forvar1121 = (1'h0); (forvar1121 < (1'h1)); forvar1121 = (forvar1121 + (1'h1)))
                    begin
                      reg1122 <= ($unsigned(((&reg650) ?
                              $signed(reg205) : $signed(reg938))) ?
                          (reg681 ?
                              $signed(reg1019[(1'h0):(1'h0)]) : (|$unsigned(reg117))) : reg546[(3'h6):(1'h1)]);
                      reg1123 <= ($unsigned(((~|reg544) ^ (~reg973))) == (^~{reg763[(4'hb):(4'h8)]}));
                      reg1124 <= reg553[(1'h0):(1'h0)];
                    end
                  for (forvar1125 = (1'h0); (forvar1125 < (1'h0)); forvar1125 = (forvar1125 + (1'h1)))
                    begin
                      reg1126 <= (reg701[(4'hd):(3'h7)] || (^~$signed((8'ha4))));
                      reg1127 <= reg652;
                    end
                  if ($unsigned(reg843[(2'h3):(1'h0)]))
                    begin
                      reg1128 <= ({{{reg518}}} == reg586[(2'h3):(2'h2)]);
                      reg1129 <= reg66;
                      reg1130 <= $signed(reg593);
                      reg1131 <= (&(reg22[(4'hc):(4'h8)] ?
                          $signed(reg221[(1'h0):(1'h0)]) : $unsigned({reg1091})));
                    end
                  else
                    begin
                      reg1128 <= reg76;
                      reg1129 <= ((reg506[(1'h1):(1'h1)] ?
                              $signed(reg905) : ($unsigned((8'h9c)) ?
                                  (reg973 <<< reg979) : reg962[(2'h2):(1'h1)])) ?
                          (~^((reg133 >>> reg1097) < reg1045)) : (reg855[(3'h5):(3'h4)] * reg511));
                    end
                end
              else
                begin
                  for (forvar1121 = (1'h0); (forvar1121 < (1'h0)); forvar1121 = (forvar1121 + (1'h1)))
                    begin
                      reg1122 <= reg698[(1'h1):(1'h0)];
                      reg1123 <= {reg192};
                      reg1124 <= reg1089;
                      reg1125 <= reg644[(2'h2):(2'h2)];
                    end
                end
              if ((reg497 ?
                  (reg982[(1'h1):(1'h1)] == {(reg555 ?
                          reg687 : reg930)}) : $unsigned($unsigned((+reg795)))))
                begin
                  reg1132 <= $signed(((8'haa) ?
                      $unsigned(reg978[(2'h3):(2'h2)]) : (reg834 ?
                          (~^reg563) : reg1120[(3'h7):(1'h0)])));
                  for (forvar1133 = (1'h0); (forvar1133 < (2'h2)); forvar1133 = (forvar1133 + (1'h1)))
                    begin
                      reg1134 <= reg561;
                      reg1135 <= {$signed({(reg555 ? reg207 : reg981)})};
                      reg1136 <= (({reg796} + reg1011) <<< reg194[(4'hc):(3'h7)]);
                    end
                  if (((^~(|(reg1049 == reg1132))) * reg554[(2'h3):(1'h0)]))
                    begin
                      reg1137 <= $signed({reg828[(3'h6):(2'h2)]});
                    end
                  else
                    begin
                      reg1137 <= reg960[(3'h6):(3'h5)];
                      reg1138 <= (-(8'hb3));
                    end
                  for (forvar1139 = (1'h0); (forvar1139 < (1'h1)); forvar1139 = (forvar1139 + (1'h1)))
                    begin
                      reg1140 <= forvar1074[(2'h3):(2'h3)];
                      reg1141 <= reg142[(2'h2):(1'h1)];
                      reg1142 <= ((~&((reg609 >= reg117) | (~&(8'h9e)))) && (8'ha8));
                      reg1143 <= $unsigned((&{(reg873 >> (8'h9e))}));
                    end
                end
              else
                begin
                  if ((^reg188))
                    begin
                      reg1132 <= reg1143[(3'h4):(2'h2)];
                      reg1133 <= (-({((8'h9e) ? reg939 : reg145)} ?
                          $signed(reg1134[(2'h3):(1'h1)]) : $signed((8'ha7))));
                      reg1134 <= $unsigned($unsigned($unsigned(reg616)));
                    end
                  else
                    begin
                      reg1132 <= $unsigned($unsigned(forvar1063));
                      reg1133 <= reg653;
                    end
                  if ((~^reg742))
                    begin
                      reg1135 <= (reg770 <= (($unsigned(reg526) ?
                          (reg803 ?
                              reg207 : wire8) : $unsigned(reg795)) - (&reg1076[(2'h3):(2'h2)])));
                      reg1136 <= reg198;
                      reg1137 <= (!$unsigned((^~(reg124 < reg639))));
                      reg1138 <= {(+{{reg883}})};
                    end
                  else
                    begin
                      reg1135 <= ($signed(reg50) ?
                          {{reg195}} : {reg687[(3'h5):(3'h4)]});
                      reg1136 <= (($unsigned($signed(reg578)) != (~(8'ha6))) <= ((reg940[(3'h7):(1'h1)] + ((8'hab) | reg1055)) - ((reg535 ?
                              reg42 : reg893) ?
                          (+reg129) : $unsigned(reg530))));
                      reg1137 <= ($unsigned(reg939[(2'h2):(2'h2)]) & ($unsigned({(8'ha7)}) < reg731[(2'h3):(1'h1)]));
                    end
                end
            end
          if ((((reg76[(2'h3):(1'h0)] != {(8'hba)}) ?
                  $unsigned(reg797[(4'hc):(2'h2)]) : ((reg638 >= reg860) << (~&reg779))) ?
              reg534[(3'h6):(3'h6)] : {$signed(reg139[(3'h6):(2'h3)])}))
            begin
              for (forvar1144 = (1'h0); (forvar1144 < (1'h0)); forvar1144 = (forvar1144 + (1'h1)))
                begin
                  for (forvar1145 = (1'h0); (forvar1145 < (2'h2)); forvar1145 = (forvar1145 + (1'h1)))
                    begin
                      reg1146 <= $unsigned(reg877);
                      reg1147 <= ((&$unsigned((!reg535))) + $unsigned(((reg1020 <= reg952) | $unsigned(forvar1125))));
                      reg1148 <= (($unsigned($unsigned((8'hba))) || reg720[(1'h1):(1'h1)]) >> (reg987 != reg820));
                      reg1149 <= $unsigned(reg917[(1'h0):(1'h0)]);
                    end
                  if ($signed($unsigned($signed((8'hb4)))))
                    begin
                      reg1150 <= (reg579 ?
                          ((8'hab) ?
                              $signed((reg883 ~^ (8'h9f))) : reg1136[(1'h1):(1'h0)]) : $signed(reg650[(2'h3):(1'h0)]));
                      reg1151 <= $unsigned($unsigned(reg501[(3'h6):(2'h2)]));
                      reg1152 <= $signed(reg696);
                      reg1153 <= $unsigned(reg729);
                    end
                  else
                    begin
                      reg1150 <= (!$unsigned((~&$unsigned((8'ha6)))));
                      reg1151 <= (((reg670 ~^ {reg745}) <= ((~^forvar1100) >> reg976)) && (reg1034[(4'h8):(3'h6)] >= reg36));
                      reg1152 <= (^~{{$unsigned(reg702)}});
                    end
                  if (reg1080)
                    begin
                      reg1154 <= forvar1103[(1'h1):(1'h1)];
                      reg1155 <= $signed({forvar1144[(3'h5):(1'h0)]});
                      reg1156 <= {$unsigned({reg1093})};
                      reg1157 <= reg741[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg1154 <= reg579;
                      reg1155 <= (~|(^{$signed(reg734)}));
                    end
                end
              if (((^~$signed((forvar1098 ?
                  reg1133 : reg216))) == reg790[(5'h10):(1'h1)]))
                begin
                  if (($signed(reg590) <= (|reg686[(3'h7):(2'h3)])))
                    begin
                      reg1158 <= $unsigned($signed({(+reg1116)}));
                      reg1159 <= reg877[(2'h2):(2'h2)];
                      reg1160 <= $signed(reg1110);
                      reg1161 <= (reg523 >>> $unsigned($signed(reg496)));
                    end
                  else
                    begin
                      reg1158 <= $signed(($unsigned(forvar1078[(1'h1):(1'h0)]) ?
                          ($unsigned(reg47) && (reg582 ?
                              reg214 : reg534)) : $signed((^~reg807))));
                      reg1159 <= reg968[(3'h6):(2'h3)];
                      reg1160 <= (~&$signed((~&reg967[(2'h2):(1'h0)])));
                      reg1161 <= (!$unsigned((reg200[(3'h5):(2'h3)] >= {reg1069})));
                    end
                  for (forvar1162 = (1'h0); (forvar1162 < (2'h2)); forvar1162 = (forvar1162 + (1'h1)))
                    begin
                      reg1163 <= (reg511 - $signed($unsigned((reg558 >>> (8'ha7)))));
                      reg1164 <= ((~^$signed(reg635)) + ((forvar1133[(3'h5):(3'h4)] || (reg627 & reg116)) <= $signed(reg33)));
                      reg1165 <= {(&reg958)};
                    end
                end
              else
                begin
                  if ($signed(($unsigned(reg814[(4'h9):(2'h3)]) ?
                      (8'ha1) : ((reg1136 - reg582) ? reg840 : reg981))))
                    begin
                      reg1158 <= (reg167[(2'h2):(2'h2)] ?
                          reg872[(1'h1):(1'h0)] : $signed((8'hb0)));
                      reg1159 <= reg1058;
                    end
                  else
                    begin
                      reg1158 <= reg193;
                      reg1159 <= ({reg790[(4'ha):(3'h5)]} ?
                          $unsigned($unsigned(((8'ha6) ?
                              reg838 : reg988))) : ($unsigned((reg115 + reg1125)) ?
                              ((8'ha7) ?
                                  $signed(reg503) : $signed(reg872)) : ((-reg717) < {reg187})));
                      reg1160 <= (~^($unsigned((reg98 ?
                          reg931 : (8'ha8))) * reg1095));
                      reg1161 <= reg1116[(3'h6):(3'h6)];
                    end
                end
            end
          else
            begin
              for (forvar1144 = (1'h0); (forvar1144 < (1'h1)); forvar1144 = (forvar1144 + (1'h1)))
                begin
                  reg1145 <= (^(((-reg698) >= (reg1153 << reg717)) ?
                      {(8'haf)} : (reg903 ?
                          {reg811} : (reg150 ? (8'ha4) : (8'ha9)))));
                end
              for (forvar1146 = (1'h0); (forvar1146 < (1'h1)); forvar1146 = (forvar1146 + (1'h1)))
                begin
                  if (reg593)
                    begin
                      reg1147 <= $unsigned(reg608);
                      reg1148 <= reg1021[(3'h7):(3'h6)];
                      reg1149 <= $signed((reg722 ?
                          $unsigned((8'ha9)) : reg896));
                    end
                  else
                    begin
                      reg1147 <= reg47;
                      reg1148 <= $unsigned(((~|(~&reg983)) ?
                          $unsigned($signed(reg533)) : $unsigned(reg1137)));
                      reg1149 <= {reg1021};
                      reg1150 <= ({((reg992 ?
                              reg801 : reg95) != $unsigned(reg140))} && $unsigned($signed($signed((8'ha7)))));
                    end
                  for (forvar1151 = (1'h0); (forvar1151 < (1'h1)); forvar1151 = (forvar1151 + (1'h1)))
                    begin
                      reg1152 <= ((|reg629[(3'h7):(1'h0)]) - ($signed(reg95) ?
                          reg922[(2'h3):(1'h0)] : ($unsigned(forvar1144) ?
                              (reg1101 ? reg17 : reg612) : $signed(reg610))));
                      reg1153 <= reg867;
                      reg1154 <= $signed(($signed($unsigned(reg762)) ?
                          $signed((reg1037 ?
                              (8'h9d) : reg151)) : ((reg905 > (8'hb6)) && (~^reg678))));
                      reg1155 <= reg111[(2'h2):(1'h0)];
                    end
                  reg1156 <= ({{reg517[(1'h0):(1'h0)]}} ?
                      (^reg1051[(1'h0):(1'h0)]) : $signed({reg980}));
                end
            end
          for (forvar1166 = (1'h0); (forvar1166 < (2'h2)); forvar1166 = (forvar1166 + (1'h1)))
            begin
              if ($unsigned({((~|reg947) ?
                      (reg627 ? reg545 : reg150) : (~reg494))}))
                begin
                  for (forvar1167 = (1'h0); (forvar1167 < (1'h1)); forvar1167 = (forvar1167 + (1'h1)))
                    begin
                      reg1168 <= reg815[(5'h10):(4'hc)];
                      reg1169 <= (!(reg604[(4'ha):(4'h8)] ?
                          ((reg984 >> (8'ha5)) >= (reg507 || reg1057)) : (8'hb4)));
                      reg1170 <= ($unsigned(((~^reg920) ?
                              $unsigned(reg1111) : reg145[(1'h0):(1'h0)])) ?
                          (-($signed(reg546) << $unsigned((8'ha2)))) : (~{$signed(forvar1083)}));
                    end
                  for (forvar1171 = (1'h0); (forvar1171 < (1'h0)); forvar1171 = (forvar1171 + (1'h1)))
                    begin
                      reg1172 <= (^{((^~reg1130) || (reg792 ?
                              reg967 : reg502))});
                      reg1173 <= {($signed((~^reg1149)) ?
                              reg1151[(1'h0):(1'h0)] : ($signed(forvar1151) ?
                                  $signed(reg893) : reg757))};
                      reg1174 <= reg193[(1'h0):(1'h0)];
                      reg1175 <= ($signed({$unsigned(reg1143)}) << (((~^(8'hb3)) ?
                              $signed(reg650) : $unsigned(reg516)) ?
                          ((!forvar1042) ?
                              (|(8'had)) : $unsigned(reg984)) : (8'hba)));
                    end
                  for (forvar1176 = (1'h0); (forvar1176 < (1'h1)); forvar1176 = (forvar1176 + (1'h1)))
                    begin
                      reg1177 <= $unsigned(reg690);
                      reg1178 <= (8'hb4);
                    end
                end
              else
                begin
                  if ((^(reg767 >>> reg1052)))
                    begin
                      reg1167 <= $unsigned({reg173});
                      reg1168 <= (8'ha3);
                      reg1169 <= $unsigned(($unsigned((8'hac)) >> reg508[(1'h1):(1'h1)]));
                      reg1170 <= $unsigned($signed((-reg891[(4'hf):(4'h8)])));
                    end
                  else
                    begin
                      reg1167 <= (reg510 ?
                          $unsigned((reg688 << {reg1157})) : $unsigned($unsigned((~(8'hb5)))));
                      reg1168 <= reg650;
                      reg1169 <= (reg1065[(2'h2):(2'h2)] << {$unsigned((reg1073 ?
                              reg989 : reg967))});
                      reg1170 <= reg1058[(4'h8):(3'h4)];
                    end
                  for (forvar1171 = (1'h0); (forvar1171 < (1'h1)); forvar1171 = (forvar1171 + (1'h1)))
                    begin
                      reg1172 <= (~^($unsigned($unsigned(reg975)) <= ($signed(reg937) * $unsigned(reg117))));
                      reg1173 <= ({(8'ha2)} ?
                          reg1167[(3'h6):(2'h2)] : $unsigned((!reg1128[(4'ha):(2'h3)])));
                      reg1174 <= ((^forvar1078) && reg73[(3'h6):(2'h2)]);
                    end
                  reg1175 <= $unsigned((8'hba));
                  if (((reg41[(3'h4):(3'h4)] ?
                          forvar1145[(3'h5):(1'h1)] : {reg581}) ?
                      (-($unsigned(reg34) ?
                          (^reg112) : (&reg168))) : $unsigned(reg524)))
                    begin
                      reg1176 <= ({$unsigned(reg127[(2'h2):(1'h1)])} ?
                          (8'hab) : (^($signed(reg1052) ?
                              (|reg879) : $unsigned((8'ha0)))));
                    end
                  else
                    begin
                      reg1176 <= ($signed($unsigned(((8'hac) & (8'hae)))) | ($unsigned(reg143) ?
                          (~&(~^(8'hb6))) : reg1042));
                    end
                end
            end
        end
    end
  assign wire1179 = (~($unsigned($unsigned((8'hb0))) || {(^~reg820)}));
  module1180 #() modinst3403 (.wire1181(reg1076), .wire1183(reg508), .y(wire3402), .wire1182(reg1099), .wire1184(reg901), .clk(clk));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1180  (y, clk, wire1181, wire1182, wire1183, wire1184);
  output wire [(32'h655):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire1181;
  input wire signed [(4'hd):(1'h0)] wire1182;
  input wire [(4'hf):(1'h0)] wire1183;
  input wire signed [(3'h4):(1'h0)] wire1184;
  wire [(3'h6):(1'h0)] wire3401;
  wire [(4'he):(1'h0)] wire3400;
  wire [(4'he):(1'h0)] wire3399;
  wire [(3'h4):(1'h0)] wire3227;
  wire [(3'h7):(1'h0)] wire3226;
  wire [(4'hd):(1'h0)] wire1185;
  wire signed [(4'h8):(1'h0)] wire3224;
  reg [(3'h5):(1'h0)] reg3398 = (1'h0);
  reg [(4'ha):(1'h0)] reg3397 = (1'h0);
  reg [(4'h9):(1'h0)] reg3395 = (1'h0);
  reg [(4'hb):(1'h0)] reg3394 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3393 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3392 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3391 = (1'h0);
  reg [(2'h2):(1'h0)] reg3390 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3388 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3380 = (1'h0);
  reg [(3'h6):(1'h0)] reg3373 = (1'h0);
  reg [(4'hd):(1'h0)] reg3387 = (1'h0);
  reg [(4'hf):(1'h0)] reg3386 = (1'h0);
  reg [(2'h2):(1'h0)] reg3385 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3384 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3383 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3382 = (1'h0);
  reg [(2'h2):(1'h0)] reg3381 = (1'h0);
  reg [(3'h6):(1'h0)] reg3379 = (1'h0);
  reg [(5'h10):(1'h0)] reg3378 = (1'h0);
  reg [(4'hf):(1'h0)] reg3377 = (1'h0);
  reg [(4'hc):(1'h0)] reg3376 = (1'h0);
  reg [(3'h5):(1'h0)] reg3375 = (1'h0);
  reg [(4'hd):(1'h0)] reg3374 = (1'h0);
  reg [(3'h7):(1'h0)] reg3371 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3370 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3369 = (1'h0);
  reg [(2'h2):(1'h0)] reg3368 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3367 = (1'h0);
  reg [(3'h5):(1'h0)] reg3366 = (1'h0);
  reg [(3'h4):(1'h0)] reg3365 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3364 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3363 = (1'h0);
  reg [(3'h7):(1'h0)] reg3360 = (1'h0);
  reg [(3'h5):(1'h0)] reg3359 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3358 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3357 = (1'h0);
  reg [(3'h5):(1'h0)] reg3355 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3353 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3352 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3351 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3350 = (1'h0);
  reg [(3'h7):(1'h0)] reg3349 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3348 = (1'h0);
  reg [(4'he):(1'h0)] reg3347 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3344 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3340 = (1'h0);
  reg [(4'hf):(1'h0)] reg3339 = (1'h0);
  reg [(4'hf):(1'h0)] reg3337 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3335 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3334 = (1'h0);
  reg [(3'h6):(1'h0)] reg3333 = (1'h0);
  reg [(4'hc):(1'h0)] reg3332 = (1'h0);
  reg [(2'h3):(1'h0)] reg3329 = (1'h0);
  reg [(4'hb):(1'h0)] reg3331 = (1'h0);
  reg [(4'hd):(1'h0)] reg3330 = (1'h0);
  reg [(4'hb):(1'h0)] reg3328 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3327 = (1'h0);
  reg [(3'h5):(1'h0)] reg3326 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3325 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3323 = (1'h0);
  reg [(2'h3):(1'h0)] reg3322 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3320 = (1'h0);
  reg [(4'hc):(1'h0)] reg3319 = (1'h0);
  reg [(3'h7):(1'h0)] reg3318 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3317 = (1'h0);
  reg [(2'h2):(1'h0)] reg3315 = (1'h0);
  reg [(5'h10):(1'h0)] reg3314 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3311 = (1'h0);
  reg [(4'hb):(1'h0)] reg3306 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3313 = (1'h0);
  reg [(3'h4):(1'h0)] reg3312 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3310 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3309 = (1'h0);
  reg [(4'hc):(1'h0)] reg3308 = (1'h0);
  reg [(2'h3):(1'h0)] reg3307 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3305 = (1'h0);
  reg [(5'h10):(1'h0)] reg3303 = (1'h0);
  reg [(4'h9):(1'h0)] reg3302 = (1'h0);
  reg [(4'ha):(1'h0)] reg3301 = (1'h0);
  reg [(4'h8):(1'h0)] reg3300 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3298 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3297 = (1'h0);
  reg [(4'hd):(1'h0)] reg3294 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3293 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3292 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3291 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3288 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3282 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3280 = (1'h0);
  reg [(3'h6):(1'h0)] reg3287 = (1'h0);
  reg [(4'he):(1'h0)] reg3286 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3285 = (1'h0);
  reg [(2'h2):(1'h0)] reg3284 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3283 = (1'h0);
  reg [(3'h6):(1'h0)] reg3281 = (1'h0);
  reg [(4'h8):(1'h0)] reg3279 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3277 = (1'h0);
  reg [(4'he):(1'h0)] reg3276 = (1'h0);
  reg [(4'ha):(1'h0)] reg3274 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3273 = (1'h0);
  reg [(5'h10):(1'h0)] reg3272 = (1'h0);
  reg [(2'h2):(1'h0)] reg3270 = (1'h0);
  reg [(2'h3):(1'h0)] reg3269 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3268 = (1'h0);
  reg [(4'hf):(1'h0)] reg3267 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3266 = (1'h0);
  reg [(2'h2):(1'h0)] reg3265 = (1'h0);
  reg [(5'h10):(1'h0)] reg3264 = (1'h0);
  reg [(2'h3):(1'h0)] reg3261 = (1'h0);
  reg [(3'h4):(1'h0)] reg3260 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3259 = (1'h0);
  reg [(2'h3):(1'h0)] reg3258 = (1'h0);
  reg [(4'hb):(1'h0)] reg3257 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3256 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3255 = (1'h0);
  reg [(2'h3):(1'h0)] reg3254 = (1'h0);
  reg [(5'h10):(1'h0)] reg3253 = (1'h0);
  reg [(3'h4):(1'h0)] reg3251 = (1'h0);
  reg [(2'h2):(1'h0)] reg3250 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3249 = (1'h0);
  reg [(4'hc):(1'h0)] reg3248 = (1'h0);
  reg [(4'ha):(1'h0)] reg3246 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3245 = (1'h0);
  reg [(4'ha):(1'h0)] reg3244 = (1'h0);
  reg [(5'h10):(1'h0)] reg3243 = (1'h0);
  reg [(3'h4):(1'h0)] reg3242 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3241 = (1'h0);
  reg [(4'hd):(1'h0)] reg3239 = (1'h0);
  reg [(3'h5):(1'h0)] reg3238 = (1'h0);
  reg [(4'h9):(1'h0)] reg3237 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3236 = (1'h0);
  reg [(2'h3):(1'h0)] reg3235 = (1'h0);
  reg [(4'hd):(1'h0)] reg3234 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3233 = (1'h0);
  reg [(2'h2):(1'h0)] reg3229 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3396 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3389 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3380 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3373 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3372 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3362 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3361 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3356 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3354 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3346 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3345 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3343 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3342 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3341 = (1'h0);
  reg [(4'he):(1'h0)] forvar3338 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3336 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3329 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3324 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3321 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3316 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3313 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3305 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3311 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3306 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3304 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3299 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3296 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3295 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3290 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3289 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3282 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3280 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3278 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3275 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3271 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3263 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3262 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3252 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3247 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3240 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3232 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3231 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3230 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3228 = (1'h0);
  assign y = {wire3401,
                 wire3400,
                 wire3399,
                 wire3227,
                 wire3226,
                 wire1185,
                 wire3224,
                 reg3398,
                 reg3397,
                 reg3395,
                 reg3394,
                 reg3393,
                 reg3392,
                 reg3391,
                 reg3390,
                 reg3388,
                 reg3380,
                 reg3373,
                 reg3387,
                 reg3386,
                 reg3385,
                 reg3384,
                 reg3383,
                 reg3382,
                 reg3381,
                 reg3379,
                 reg3378,
                 reg3377,
                 reg3376,
                 reg3375,
                 reg3374,
                 reg3371,
                 reg3370,
                 reg3369,
                 reg3368,
                 reg3367,
                 reg3366,
                 reg3365,
                 reg3364,
                 reg3363,
                 reg3360,
                 reg3359,
                 reg3358,
                 reg3357,
                 reg3355,
                 reg3353,
                 reg3352,
                 reg3351,
                 reg3350,
                 reg3349,
                 reg3348,
                 reg3347,
                 reg3344,
                 reg3340,
                 reg3339,
                 reg3337,
                 reg3335,
                 reg3334,
                 reg3333,
                 reg3332,
                 reg3329,
                 reg3331,
                 reg3330,
                 reg3328,
                 reg3327,
                 reg3326,
                 reg3325,
                 reg3323,
                 reg3322,
                 reg3320,
                 reg3319,
                 reg3318,
                 reg3317,
                 reg3315,
                 reg3314,
                 reg3311,
                 reg3306,
                 reg3313,
                 reg3312,
                 reg3310,
                 reg3309,
                 reg3308,
                 reg3307,
                 reg3305,
                 reg3303,
                 reg3302,
                 reg3301,
                 reg3300,
                 reg3298,
                 reg3297,
                 reg3294,
                 reg3293,
                 reg3292,
                 reg3291,
                 reg3288,
                 reg3282,
                 reg3280,
                 reg3287,
                 reg3286,
                 reg3285,
                 reg3284,
                 reg3283,
                 reg3281,
                 reg3279,
                 reg3277,
                 reg3276,
                 reg3274,
                 reg3273,
                 reg3272,
                 reg3270,
                 reg3269,
                 reg3268,
                 reg3267,
                 reg3266,
                 reg3265,
                 reg3264,
                 reg3261,
                 reg3260,
                 reg3259,
                 reg3258,
                 reg3257,
                 reg3256,
                 reg3255,
                 reg3254,
                 reg3253,
                 reg3251,
                 reg3250,
                 reg3249,
                 reg3248,
                 reg3246,
                 reg3245,
                 reg3244,
                 reg3243,
                 reg3242,
                 reg3241,
                 reg3239,
                 reg3238,
                 reg3237,
                 reg3236,
                 reg3235,
                 reg3234,
                 reg3233,
                 reg3229,
                 forvar3396,
                 forvar3389,
                 forvar3380,
                 forvar3373,
                 forvar3372,
                 forvar3362,
                 forvar3361,
                 forvar3356,
                 forvar3354,
                 forvar3346,
                 forvar3345,
                 forvar3343,
                 forvar3342,
                 forvar3341,
                 forvar3338,
                 forvar3336,
                 forvar3329,
                 forvar3324,
                 forvar3321,
                 forvar3316,
                 forvar3313,
                 forvar3305,
                 forvar3311,
                 forvar3306,
                 forvar3304,
                 forvar3299,
                 forvar3296,
                 forvar3295,
                 forvar3290,
                 forvar3289,
                 forvar3282,
                 forvar3280,
                 forvar3278,
                 forvar3275,
                 forvar3271,
                 forvar3263,
                 forvar3262,
                 forvar3252,
                 forvar3247,
                 forvar3240,
                 forvar3232,
                 forvar3231,
                 forvar3230,
                 forvar3228,
                 (1'h0)};
  assign wire1185 = wire1184[(3'h4):(2'h3)];
  module1186 #() modinst3225 (.wire1189(wire1183), .wire1188(wire1181), .wire1187(wire1184), .y(wire3224), .clk(clk), .wire1190(wire1185), .wire1191(wire1182));
  assign wire3226 = (($unsigned(wire1185) ?
                        $unsigned(wire1185[(4'h8):(3'h4)]) : ($unsigned((8'hab)) ?
                            $signed(wire1183) : {(8'hb9)})) & (+(!$unsigned((8'hb7)))));
  assign wire3227 = (({wire1183} ? $unsigned((-(8'hb8))) : wire3226) ?
                        (($signed(wire3224) ?
                                $signed(wire1182) : (wire1184 < wire1184)) ?
                            wire1184 : (+(wire1181 ?
                                wire3224 : (8'hb3)))) : wire1183);
  always
    @(posedge clk) begin
      for (forvar3228 = (1'h0); (forvar3228 < (2'h3)); forvar3228 = (forvar3228 + (1'h1)))
        begin
          reg3229 <= $signed((wire3227[(3'h4):(2'h3)] >= $unsigned(wire3224[(4'h8):(4'h8)])));
          for (forvar3230 = (1'h0); (forvar3230 < (2'h3)); forvar3230 = (forvar3230 + (1'h1)))
            begin
              for (forvar3231 = (1'h0); (forvar3231 < (1'h0)); forvar3231 = (forvar3231 + (1'h1)))
                begin
                  for (forvar3232 = (1'h0); (forvar3232 < (2'h3)); forvar3232 = (forvar3232 + (1'h1)))
                    begin
                      reg3233 <= $unsigned((wire1181 ?
                          wire3227[(2'h2):(1'h1)] : ($unsigned(reg3229) ?
                              $unsigned((8'h9f)) : $signed(wire3226))));
                      reg3234 <= ({(wire1184 ?
                              (forvar3232 ?
                                  wire3227 : forvar3232) : $unsigned(wire1185))} ~^ (($unsigned(wire1181) * forvar3230) && $signed($signed(wire3226))));
                    end
                  reg3235 <= ($signed({(8'had)}) <<< wire1183[(4'ha):(4'ha)]);
                  if (reg3235)
                    begin
                      reg3236 <= (wire1181 ?
                          reg3233[(1'h0):(1'h0)] : (forvar3231 ?
                              ((8'ha2) ?
                                  (forvar3228 <= wire1185) : $unsigned(wire1181)) : $unsigned($signed(reg3229))));
                      reg3237 <= ((wire1181 ?
                              $signed(wire1181[(4'ha):(2'h3)]) : reg3234) ?
                          forvar3230[(4'h8):(2'h2)] : (&wire1184[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg3236 <= (-({(8'h9f)} <= forvar3228[(3'h4):(2'h2)]));
                      reg3237 <= $unsigned(reg3234);
                      reg3238 <= ((&(forvar3228 ^ $signed((8'ha1)))) ?
                          $signed({(wire1185 ?
                                  forvar3230 : wire1181)}) : $unsigned($signed(reg3229)));
                      reg3239 <= (forvar3228 >>> (~|reg3236[(3'h7):(3'h5)]));
                    end
                  for (forvar3240 = (1'h0); (forvar3240 < (2'h3)); forvar3240 = (forvar3240 + (1'h1)))
                    begin
                      reg3241 <= $signed((^wire1183));
                      reg3242 <= ({wire1183} ?
                          forvar3230[(4'hb):(3'h6)] : forvar3230[(2'h2):(1'h0)]);
                    end
                end
              if ((|$unsigned(forvar3230[(4'h8):(1'h0)])))
                begin
                  if ($signed({(reg3241[(1'h0):(1'h0)] ?
                          (+wire1183) : (reg3236 ? (8'ha6) : reg3233))}))
                    begin
                      reg3243 <= (~&(~&reg3238[(2'h3):(1'h1)]));
                      reg3244 <= reg3236[(3'h7):(2'h3)];
                      reg3245 <= (wire3227[(1'h0):(1'h0)] < forvar3231);
                    end
                  else
                    begin
                      reg3243 <= wire3227[(1'h0):(1'h0)];
                      reg3244 <= forvar3231;
                      reg3245 <= $unsigned($unsigned(reg3241));
                    end
                end
              else
                begin
                  if (reg3244[(2'h2):(1'h1)])
                    begin
                      reg3243 <= reg3233;
                      reg3244 <= ($unsigned((8'h9d)) + ($unsigned((wire3227 ?
                          wire1184 : reg3243)) || ((reg3245 || wire3227) ?
                          $signed(forvar3232) : (forvar3230 ?
                              wire1183 : reg3239))));
                    end
                  else
                    begin
                      reg3243 <= (($signed(reg3236) & reg3237[(3'h7):(2'h3)]) ?
                          wire3224 : $unsigned((reg3238[(3'h4):(2'h2)] || forvar3232[(1'h1):(1'h0)])));
                    end
                  reg3245 <= $signed((({reg3238} ?
                      {(8'h9c)} : reg3238) << (~|(reg3245 << reg3235))));
                  reg3246 <= (8'ha5);
                end
              for (forvar3247 = (1'h0); (forvar3247 < (2'h3)); forvar3247 = (forvar3247 + (1'h1)))
                begin
                  if ((^~wire1183))
                    begin
                      reg3248 <= reg3245;
                      reg3249 <= (-$signed({reg3237[(3'h7):(1'h1)]}));
                      reg3250 <= (reg3239[(4'ha):(2'h2)] - $signed((^(^~forvar3228))));
                      reg3251 <= (8'ha5);
                    end
                  else
                    begin
                      reg3248 <= $unsigned(($unsigned($signed(forvar3240)) >>> reg3250));
                    end
                  for (forvar3252 = (1'h0); (forvar3252 < (1'h1)); forvar3252 = (forvar3252 + (1'h1)))
                    begin
                      reg3253 <= (8'hb8);
                      reg3254 <= $signed((~^((^reg3238) * $signed(forvar3228))));
                    end
                  if (wire3227)
                    begin
                      reg3255 <= wire3224[(3'h6):(2'h2)];
                      reg3256 <= $unsigned(($unsigned(forvar3240[(1'h1):(1'h0)]) ?
                          {(reg3254 ?
                                  reg3239 : (8'hb5))} : {(reg3248 << (8'hb4))}));
                      reg3257 <= forvar3247;
                      reg3258 <= forvar3252[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3255 <= (reg3243[(4'ha):(2'h2)] ?
                          $signed(reg3244) : reg3234);
                      reg3256 <= $unsigned({reg3242});
                      reg3257 <= ((|{$signed(wire1185)}) ?
                          $unsigned((^reg3233)) : (8'ha1));
                    end
                  if ($unsigned(wire1183[(4'hd):(4'h8)]))
                    begin
                      reg3259 <= (~^($signed($signed((8'ha0))) * (8'ha0)));
                      reg3260 <= wire1185;
                      reg3261 <= $unsigned($signed(($unsigned(reg3257) ?
                          ((8'hb4) ? wire1184 : reg3246) : (wire1183 ?
                              wire1184 : (8'ha9)))));
                    end
                  else
                    begin
                      reg3259 <= reg3229[(1'h1):(1'h0)];
                      reg3260 <= reg3251[(1'h1):(1'h0)];
                    end
                end
            end
          for (forvar3262 = (1'h0); (forvar3262 < (1'h0)); forvar3262 = (forvar3262 + (1'h1)))
            begin
              for (forvar3263 = (1'h0); (forvar3263 < (1'h1)); forvar3263 = (forvar3263 + (1'h1)))
                begin
                  if (forvar3230[(3'h5):(1'h0)])
                    begin
                      reg3264 <= $unsigned(({(forvar3240 ? reg3251 : reg3238)} ?
                          ((~forvar3252) ?
                              forvar3252 : wire3227[(1'h0):(1'h0)]) : {{wire1182}}));
                      reg3265 <= $signed((&$unsigned((forvar3232 ?
                          (8'hb6) : reg3261))));
                      reg3266 <= (8'hb8);
                      reg3267 <= $signed(((~|reg3259) ?
                          (!forvar3247) : reg3256));
                    end
                  else
                    begin
                      reg3264 <= wire1182;
                      reg3265 <= (|(+{reg3249}));
                      reg3266 <= $unsigned((($unsigned(forvar3232) ?
                              (-forvar3232) : reg3241) ?
                          $signed($unsigned(reg3259)) : $signed(reg3249[(3'h4):(1'h0)])));
                      reg3267 <= forvar3240;
                    end
                  if ((($signed((|reg3238)) >>> (|(reg3264 <= forvar3230))) - (~$unsigned(((8'hb8) >>> reg3251)))))
                    begin
                      reg3268 <= ($unsigned(reg3245) && $signed((reg3258 ?
                          (8'hb4) : $unsigned(reg3235))));
                      reg3269 <= wire3226[(1'h0):(1'h0)];
                      reg3270 <= $unsigned($unsigned(({forvar3232} ?
                          $signed((8'ha9)) : (|reg3236))));
                    end
                  else
                    begin
                      reg3268 <= (+reg3250[(2'h2):(1'h0)]);
                      reg3269 <= reg3267;
                      reg3270 <= $unsigned($signed($unsigned((reg3257 ~^ wire3224))));
                    end
                  for (forvar3271 = (1'h0); (forvar3271 < (1'h1)); forvar3271 = (forvar3271 + (1'h1)))
                    begin
                      reg3272 <= {(-(&(forvar3271 ? (8'ha4) : reg3261)))};
                      reg3273 <= ((((forvar3263 | reg3264) > (^~reg3254)) ?
                          ($unsigned((8'ha1)) ?
                              (reg3238 == forvar3263) : reg3261) : reg3242[(1'h0):(1'h0)]) << $unsigned($signed($unsigned(reg3233))));
                      reg3274 <= ((8'ha4) ?
                          ($unsigned($unsigned(reg3255)) || (reg3236[(4'hb):(3'h7)] * {wire1184})) : $unsigned((|reg3257)));
                    end
                  for (forvar3275 = (1'h0); (forvar3275 < (1'h0)); forvar3275 = (forvar3275 + (1'h1)))
                    begin
                      reg3276 <= (((~&{wire3227}) ? forvar3271 : reg3260) ?
                          reg3238[(2'h2):(1'h0)] : (^~reg3248[(1'h0):(1'h0)]));
                      reg3277 <= $unsigned((~^((-reg3257) | (8'ha7))));
                    end
                end
            end
        end
      for (forvar3278 = (1'h0); (forvar3278 < (2'h3)); forvar3278 = (forvar3278 + (1'h1)))
        begin
          reg3279 <= reg3242[(1'h0):(1'h0)];
          if (reg3257[(4'h9):(2'h2)])
            begin
              for (forvar3280 = (1'h0); (forvar3280 < (1'h1)); forvar3280 = (forvar3280 + (1'h1)))
                begin
                  reg3281 <= reg3257;
                  for (forvar3282 = (1'h0); (forvar3282 < (2'h3)); forvar3282 = (forvar3282 + (1'h1)))
                    begin
                      reg3283 <= $unsigned($signed($unsigned(reg3274)));
                      reg3284 <= (((~(forvar3228 >>> reg3258)) ?
                          wire1182[(3'h5):(2'h3)] : reg3283[(1'h0):(1'h0)]) <= $unsigned($signed((^forvar3231))));
                      reg3285 <= reg3277;
                      reg3286 <= $unsigned((|$unsigned(((8'ha6) ^~ (8'hb3)))));
                    end
                  reg3287 <= ($unsigned($signed((reg3283 - reg3250))) + $unsigned($unsigned({forvar3230})));
                end
            end
          else
            begin
              if (forvar3228[(3'h6):(3'h4)])
                begin
                  if ($unsigned({(8'haa)}))
                    begin
                      reg3280 <= $unsigned($unsigned($unsigned(reg3274[(3'h7):(3'h7)])));
                      reg3281 <= (&reg3268[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg3280 <= {$signed((8'h9e))};
                      reg3281 <= (~reg3238[(2'h3):(1'h0)]);
                      reg3282 <= (reg3283[(3'h4):(1'h1)] ?
                          {{reg3260[(3'h4):(2'h2)]}} : $signed((reg3260[(1'h1):(1'h0)] ?
                              $unsigned(reg3244) : (reg3274 ?
                                  (8'hb1) : reg3248))));
                    end
                  if ((&(((~&reg3234) ?
                      forvar3232 : (reg3254 >>> (8'ha2))) ^~ reg3254[(1'h1):(1'h1)])))
                    begin
                      reg3283 <= (~^(+$signed((+reg3235))));
                      reg3284 <= $signed((-(reg3279 > $signed(reg3244))));
                      reg3285 <= ($unsigned(((reg3261 < wire1183) ?
                              reg3253 : $unsigned(reg3283))) ?
                          (&((reg3257 ? reg3268 : (8'ha2)) ?
                              wire3227 : (8'hac))) : $unsigned(((reg3273 ?
                                  forvar3240 : wire3227) ?
                              $unsigned(wire1183) : $signed(forvar3247))));
                    end
                  else
                    begin
                      reg3283 <= reg3277;
                      reg3284 <= (((&reg3284) == {$unsigned(wire3226)}) ?
                          (~|wire3224) : (reg3273[(1'h0):(1'h0)] & $unsigned((!reg3248))));
                      reg3285 <= ((((reg3279 ? forvar3275 : (8'h9d)) ?
                          (&reg3265) : $signed(reg3237)) & (8'ha7)) >= (^$unsigned((8'ha9))));
                      reg3286 <= reg3242;
                    end
                  reg3287 <= ((&$signed((^reg3276))) ?
                      (!(-reg3266)) : wire3227);
                  reg3288 <= (8'hae);
                end
              else
                begin
                  reg3280 <= $signed((8'hb4));
                end
              for (forvar3289 = (1'h0); (forvar3289 < (1'h0)); forvar3289 = (forvar3289 + (1'h1)))
                begin
                  for (forvar3290 = (1'h0); (forvar3290 < (2'h2)); forvar3290 = (forvar3290 + (1'h1)))
                    begin
                      reg3291 <= $unsigned((reg3279 << $unsigned(reg3256)));
                    end
                  if ($signed(((reg3272[(3'h6):(1'h0)] >> {(8'hac)}) ?
                      (^wire1185) : wire1181)))
                    begin
                      reg3292 <= (reg3279 ^ forvar3280);
                      reg3293 <= (reg3244[(4'h8):(3'h4)] ?
                          reg3239[(1'h0):(1'h0)] : (reg3259[(3'h4):(2'h3)] - {forvar3275[(3'h4):(3'h4)]}));
                    end
                  else
                    begin
                      reg3292 <= $unsigned($signed(((reg3276 != reg3288) ?
                          $unsigned((8'hb3)) : $unsigned(reg3280))));
                      reg3293 <= $unsigned((!reg3287));
                      reg3294 <= ($signed(((reg3244 ?
                          forvar3282 : forvar3271) >= (|reg3244))) >= (|(^(^~(8'hb5)))));
                    end
                end
              for (forvar3295 = (1'h0); (forvar3295 < (2'h2)); forvar3295 = (forvar3295 + (1'h1)))
                begin
                  for (forvar3296 = (1'h0); (forvar3296 < (2'h2)); forvar3296 = (forvar3296 + (1'h1)))
                    begin
                      reg3297 <= forvar3252;
                      reg3298 <= (~|($signed((reg3235 * reg3291)) ?
                          ((+reg3277) ?
                              reg3276 : forvar3282[(4'ha):(2'h2)]) : ((+reg3248) >> reg3276)));
                    end
                  for (forvar3299 = (1'h0); (forvar3299 < (1'h1)); forvar3299 = (forvar3299 + (1'h1)))
                    begin
                      reg3300 <= (&(8'hb4));
                      reg3301 <= $unsigned(reg3284[(2'h2):(1'h0)]);
                      reg3302 <= (&reg3229);
                    end
                end
            end
          reg3303 <= reg3254[(2'h2):(1'h0)];
        end
      for (forvar3304 = (1'h0); (forvar3304 < (1'h1)); forvar3304 = (forvar3304 + (1'h1)))
        begin
          if (reg3248[(1'h1):(1'h1)])
            begin
              reg3305 <= $unsigned(reg3292);
              for (forvar3306 = (1'h0); (forvar3306 < (1'h0)); forvar3306 = (forvar3306 + (1'h1)))
                begin
                  if ($unsigned((!reg3285)))
                    begin
                      reg3307 <= $signed(reg3294[(4'h8):(4'h8)]);
                      reg3308 <= $signed(reg3249);
                      reg3309 <= (((reg3239 + (reg3274 << wire3227)) >>> $signed((reg3283 ^~ reg3260))) >>> $signed({forvar3306[(4'ha):(2'h3)]}));
                      reg3310 <= (!reg3276[(4'hc):(3'h7)]);
                    end
                  else
                    begin
                      reg3307 <= forvar3271[(1'h1):(1'h1)];
                      reg3308 <= reg3264[(3'h7):(1'h1)];
                      reg3309 <= forvar3306[(3'h7):(2'h2)];
                    end
                  for (forvar3311 = (1'h0); (forvar3311 < (2'h2)); forvar3311 = (forvar3311 + (1'h1)))
                    begin
                      reg3312 <= (((&reg3305[(3'h5):(2'h3)]) + reg3229[(1'h0):(1'h0)]) ?
                          $signed(reg3235) : (((reg3241 - reg3243) ?
                                  (8'ha8) : (wire1184 == reg3286)) ?
                              {$signed(forvar3232)} : ($unsigned(forvar3299) >> (!reg3242))));
                      reg3313 <= reg3251[(2'h3):(1'h1)];
                    end
                end
            end
          else
            begin
              if ($signed((~^forvar3282)))
                begin
                  reg3305 <= reg3286[(3'h6):(1'h0)];
                  for (forvar3306 = (1'h0); (forvar3306 < (1'h0)); forvar3306 = (forvar3306 + (1'h1)))
                    begin
                      reg3307 <= forvar3282;
                    end
                end
              else
                begin
                  for (forvar3305 = (1'h0); (forvar3305 < (2'h2)); forvar3305 = (forvar3305 + (1'h1)))
                    begin
                      reg3306 <= (~$unsigned(((!(8'hab)) ?
                          (8'ha0) : reg3260[(1'h0):(1'h0)])));
                      reg3307 <= wire1181[(3'h6):(3'h4)];
                      reg3308 <= $unsigned(reg3251[(2'h3):(2'h3)]);
                    end
                  if ((^~(($signed(forvar3290) ?
                      reg3312[(2'h2):(1'h1)] : (-reg3305)) == ($unsigned(reg3233) <<< $signed(reg3282)))))
                    begin
                      reg3309 <= reg3308;
                      reg3310 <= reg3313[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3309 <= forvar3262[(2'h2):(2'h2)];
                      reg3310 <= $signed({(&(+reg3300))});
                      reg3311 <= reg3259[(3'h4):(3'h4)];
                      reg3312 <= (^~$signed($unsigned(forvar3282[(4'hc):(4'hc)])));
                    end
                  for (forvar3313 = (1'h0); (forvar3313 < (2'h2)); forvar3313 = (forvar3313 + (1'h1)))
                    begin
                      reg3314 <= (8'ha1);
                      reg3315 <= forvar3247[(3'h6):(1'h0)];
                    end
                end
              for (forvar3316 = (1'h0); (forvar3316 < (1'h0)); forvar3316 = (forvar3316 + (1'h1)))
                begin
                  if ($unsigned((!((~reg3287) ?
                      (8'hb0) : $unsigned(forvar3232)))))
                    begin
                      reg3317 <= reg3235[(2'h3):(2'h2)];
                      reg3318 <= $signed(reg3264);
                    end
                  else
                    begin
                      reg3317 <= reg3257[(3'h4):(1'h0)];
                      reg3318 <= ((-((reg3236 >= reg3301) <<< (&wire1183))) < $signed(wire3226[(1'h0):(1'h0)]));
                      reg3319 <= (((|reg3249[(4'ha):(2'h2)]) >= $unsigned((&reg3246))) ?
                          (~forvar3299) : (~reg3266[(1'h0):(1'h0)]));
                      reg3320 <= reg3305;
                    end
                  for (forvar3321 = (1'h0); (forvar3321 < (1'h1)); forvar3321 = (forvar3321 + (1'h1)))
                    begin
                      reg3322 <= $unsigned(($signed($signed(forvar3296)) ?
                          (^(reg3293 && reg3253)) : reg3294));
                      reg3323 <= (forvar3231 ?
                          (reg3267[(2'h3):(1'h0)] & $unsigned(reg3283[(3'h4):(2'h2)])) : (forvar3316 ?
                              $signed(reg3317) : (^reg3302)));
                    end
                  for (forvar3324 = (1'h0); (forvar3324 < (2'h3)); forvar3324 = (forvar3324 + (1'h1)))
                    begin
                      reg3325 <= $unsigned(({$unsigned(forvar3316)} <= (^$signed(reg3229))));
                      reg3326 <= (|(((+reg3310) ?
                              (reg3260 ?
                                  wire1184 : forvar3240) : reg3300[(2'h3):(1'h0)]) ?
                          $signed((&reg3270)) : ((reg3264 ?
                              reg3281 : reg3245) <= reg3319[(3'h7):(2'h2)])));
                      reg3327 <= $signed(reg3280[(1'h0):(1'h0)]);
                      reg3328 <= wire1184;
                    end
                end
              if ($unsigned((((forvar3305 ^ reg3251) ?
                      $unsigned(reg3284) : (&wire1181)) ?
                  $unsigned((&forvar3247)) : $signed((~reg3284)))))
                begin
                  for (forvar3329 = (1'h0); (forvar3329 < (2'h2)); forvar3329 = (forvar3329 + (1'h1)))
                    begin
                      reg3330 <= (+(~|wire3226));
                      reg3331 <= {($signed($unsigned(reg3257)) <<< $unsigned(forvar3280[(1'h0):(1'h0)]))};
                    end
                end
              else
                begin
                  if ($signed((|reg3260)))
                    begin
                      reg3329 <= $signed(($signed(reg3237[(3'h4):(3'h4)]) >>> reg3288[(3'h5):(2'h2)]));
                      reg3330 <= (!(reg3234 * {{reg3256}}));
                      reg3331 <= {$unsigned($signed(reg3293[(2'h3):(2'h3)]))};
                      reg3332 <= $unsigned(((reg3291 ?
                          (^~reg3255) : wire1185[(4'hd):(1'h1)]) ^~ (~&forvar3295[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg3329 <= (8'haf);
                      reg3330 <= (~&(&((reg3331 ? reg3298 : reg3238) ?
                          reg3318[(1'h1):(1'h0)] : {(8'hba)})));
                      reg3331 <= (~&(&reg3286));
                      reg3332 <= {(reg3288[(2'h2):(1'h1)] + reg3229)};
                    end
                  if ((reg3285[(1'h0):(1'h0)] ^~ reg3325))
                    begin
                      reg3333 <= $unsigned(((~(forvar3280 & forvar3316)) ?
                          $signed((reg3314 << forvar3313)) : $unsigned((wire1181 != reg3264))));
                    end
                  else
                    begin
                      reg3333 <= (reg3268[(3'h5):(3'h5)] ?
                          (-(reg3300[(2'h3):(2'h2)] ?
                              {reg3258} : reg3332[(1'h0):(1'h0)])) : (~&({reg3274} ?
                              (forvar3324 ? reg3283 : reg3307) : (&(8'h9e)))));
                      reg3334 <= (-(reg3256[(3'h4):(2'h2)] ?
                          ((forvar3271 - reg3254) && forvar3289) : reg3285[(3'h6):(2'h2)]));
                      reg3335 <= (((&(+reg3257)) ? (8'hae) : reg3276) ?
                          $signed(($signed(reg3244) << $signed(reg3245))) : $unsigned(reg3300));
                    end
                end
            end
          for (forvar3336 = (1'h0); (forvar3336 < (1'h1)); forvar3336 = (forvar3336 + (1'h1)))
            begin
              if ((^(wire3226 & (~|$unsigned((8'ha3))))))
                begin
                  if ($unsigned(reg3326))
                    begin
                      reg3337 <= (|reg3267);
                    end
                  else
                    begin
                      reg3337 <= (reg3320[(3'h5):(3'h5)] ?
                          forvar3231[(2'h3):(2'h2)] : (^~reg3334[(1'h1):(1'h0)]));
                    end
                end
              else
                begin
                  reg3337 <= ($unsigned((forvar3247 ?
                          (!reg3235) : $signed(reg3309))) ?
                      ($signed((~|forvar3316)) ^ reg3320) : {($signed(reg3254) ?
                              (~|(8'ha3)) : (~|wire1182))});
                  for (forvar3338 = (1'h0); (forvar3338 < (2'h2)); forvar3338 = (forvar3338 + (1'h1)))
                    begin
                      reg3339 <= forvar3231;
                      reg3340 <= reg3245[(2'h3):(2'h3)];
                    end
                end
            end
        end
      for (forvar3341 = (1'h0); (forvar3341 < (2'h3)); forvar3341 = (forvar3341 + (1'h1)))
        begin
          for (forvar3342 = (1'h0); (forvar3342 < (2'h2)); forvar3342 = (forvar3342 + (1'h1)))
            begin
              for (forvar3343 = (1'h0); (forvar3343 < (2'h3)); forvar3343 = (forvar3343 + (1'h1)))
                begin
                  reg3344 <= ($unsigned(forvar3305[(3'h4):(2'h2)]) ^~ reg3308[(2'h2):(2'h2)]);
                end
              for (forvar3345 = (1'h0); (forvar3345 < (2'h3)); forvar3345 = (forvar3345 + (1'h1)))
                begin
                  for (forvar3346 = (1'h0); (forvar3346 < (2'h3)); forvar3346 = (forvar3346 + (1'h1)))
                    begin
                      reg3347 <= $unsigned($unsigned(reg3332));
                      reg3348 <= (~(((&forvar3336) ^ reg3298[(2'h2):(1'h0)]) == ($unsigned(reg3333) >= $unsigned(reg3242))));
                    end
                  reg3349 <= (reg3329 || $unsigned($signed((wire1182 ?
                      reg3258 : reg3229))));
                  if (forvar3316[(3'h7):(1'h1)])
                    begin
                      reg3350 <= {((~|$unsigned(reg3315)) ^~ (8'ha1))};
                      reg3351 <= reg3333;
                      reg3352 <= $signed(((-$unsigned(reg3237)) ?
                          {$signed(reg3250)} : $unsigned($signed(reg3317))));
                      reg3353 <= reg3268;
                    end
                  else
                    begin
                      reg3350 <= $signed((((reg3255 <= (8'ha8)) ?
                          $unsigned((8'haa)) : ((8'hb2) >>> forvar3336)) ^~ $signed((-reg3352))));
                      reg3351 <= reg3319;
                      reg3352 <= ((!$signed((^forvar3278))) && (8'h9f));
                      reg3353 <= (((~|reg3277) <= ((8'ha0) ^ $unsigned((8'hb9)))) ^~ $signed($signed(reg3308[(4'h9):(3'h7)])));
                    end
                end
              for (forvar3354 = (1'h0); (forvar3354 < (1'h1)); forvar3354 = (forvar3354 + (1'h1)))
                begin
                  reg3355 <= reg3279[(3'h5):(1'h1)];
                  for (forvar3356 = (1'h0); (forvar3356 < (1'h0)); forvar3356 = (forvar3356 + (1'h1)))
                    begin
                      reg3357 <= {reg3320[(2'h3):(2'h2)]};
                      reg3358 <= $signed($signed((|wire1182)));
                      reg3359 <= {$unsigned($signed($unsigned(forvar3232)))};
                      reg3360 <= reg3300[(1'h0):(1'h0)];
                    end
                end
              for (forvar3361 = (1'h0); (forvar3361 < (2'h3)); forvar3361 = (forvar3361 + (1'h1)))
                begin
                  for (forvar3362 = (1'h0); (forvar3362 < (1'h1)); forvar3362 = (forvar3362 + (1'h1)))
                    begin
                      reg3363 <= (8'ha5);
                      reg3364 <= $signed(reg3273);
                      reg3365 <= (8'ha6);
                      reg3366 <= ($signed(((wire1182 == reg3285) ?
                              ((8'ha8) + reg3258) : (reg3334 ~^ reg3337))) ?
                          (~|reg3239) : (((reg3359 && reg3301) >> reg3298) ?
                              (8'ha2) : $unsigned($signed(forvar3305))));
                    end
                  if ((!reg3317))
                    begin
                      reg3367 <= $unsigned(reg3323[(3'h4):(2'h3)]);
                      reg3368 <= reg3367[(4'h8):(3'h4)];
                      reg3369 <= (8'h9e);
                      reg3370 <= (((8'hb4) ?
                          forvar3231[(3'h4):(2'h3)] : (^~(reg3334 ?
                              forvar3313 : reg3332))) <<< forvar3228);
                    end
                  else
                    begin
                      reg3367 <= ($unsigned(({(8'ha1)} ?
                          reg3301 : {reg3329})) | {$unsigned((wire1183 ?
                              forvar3230 : (8'ha1)))});
                      reg3368 <= reg3318;
                      reg3369 <= (~|(~^reg3256));
                    end
                end
            end
          reg3371 <= (~|$signed((reg3311 ?
              $unsigned(wire1185) : {forvar3299})));
          for (forvar3372 = (1'h0); (forvar3372 < (2'h2)); forvar3372 = (forvar3372 + (1'h1)))
            begin
              if (wire1182)
                begin
                  for (forvar3373 = (1'h0); (forvar3373 < (2'h2)); forvar3373 = (forvar3373 + (1'h1)))
                    begin
                      reg3374 <= (|{{(!forvar3313)}});
                      reg3375 <= ($signed($signed((reg3285 >= reg3319))) & ({(reg3249 ?
                                  reg3366 : forvar3345)} ?
                          (^~reg3355[(2'h3):(1'h0)]) : reg3229));
                      reg3376 <= {forvar3361[(3'h5):(3'h5)]};
                    end
                  if ({$unsigned($signed((&reg3363)))})
                    begin
                      reg3377 <= (8'hb9);
                    end
                  else
                    begin
                      reg3377 <= ($unsigned((-(reg3374 ~^ reg3237))) ?
                          {$signed({reg3323})} : reg3364[(3'h6):(3'h4)]);
                      reg3378 <= $unsigned((!$unsigned(reg3320)));
                      reg3379 <= (+(((forvar3305 >> forvar3338) ?
                              ((8'hb0) >= (8'hab)) : (reg3357 || (8'h9d))) ?
                          {reg3238} : ((reg3337 ?
                              reg3337 : wire3226) < $unsigned(reg3317))));
                    end
                  for (forvar3380 = (1'h0); (forvar3380 < (2'h3)); forvar3380 = (forvar3380 + (1'h1)))
                    begin
                      reg3381 <= ($unsigned(forvar3343[(3'h7):(3'h4)]) >> (8'h9e));
                      reg3382 <= $unsigned((($signed(reg3234) ?
                              ((8'ha1) ?
                                  forvar3247 : forvar3341) : $unsigned((8'hb4))) ?
                          reg3315 : forvar3329[(1'h0):(1'h0)]));
                      reg3383 <= ((^((^~forvar3280) ?
                              reg3288 : reg3352[(3'h6):(2'h3)])) ?
                          $signed($signed($signed(reg3246))) : {$unsigned({reg3381})});
                      reg3384 <= ((~|$unsigned((reg3378 - forvar3361))) <<< $unsigned(reg3284[(1'h0):(1'h0)]));
                    end
                  if ($signed((~|$signed((reg3307 & reg3238)))))
                    begin
                      reg3385 <= $signed(wire3227);
                      reg3386 <= ((reg3308[(3'h4):(2'h2)] == forvar3232) ?
                          $signed((reg3267 ?
                              reg3310[(2'h3):(2'h3)] : {(8'h9d)})) : reg3347[(3'h6):(2'h2)]);
                      reg3387 <= (~|{({forvar3282} ^ (reg3348 ?
                              reg3254 : (8'hb7)))});
                    end
                  else
                    begin
                      reg3385 <= reg3310;
                      reg3386 <= reg3297;
                    end
                end
              else
                begin
                  if (reg3303)
                    begin
                      reg3373 <= ($signed(({(8'hba)} ?
                              (^~forvar3271) : (forvar3296 ?
                                  reg3351 : (8'hae)))) ?
                          reg3358 : reg3292);
                      reg3374 <= $unsigned($unsigned((reg3292[(3'h6):(3'h6)] >>> (reg3382 == reg3318))));
                      reg3375 <= $unsigned(((reg3277 ?
                          (reg3366 >> reg3382) : $signed(forvar3290)) >>> ((~reg3307) ?
                          $signed(reg3260) : {reg3292})));
                      reg3376 <= $unsigned($signed((^(forvar3313 ?
                          reg3243 : wire1181))));
                    end
                  else
                    begin
                      reg3373 <= reg3259[(1'h0):(1'h0)];
                    end
                  if ($signed({forvar3289[(4'h9):(2'h3)]}))
                    begin
                      reg3377 <= {$signed($unsigned(reg3258[(1'h1):(1'h0)]))};
                      reg3378 <= {$signed(reg3266)};
                      reg3379 <= $unsigned($signed(reg3308[(1'h1):(1'h0)]));
                      reg3380 <= (8'ha1);
                    end
                  else
                    begin
                      reg3377 <= (8'h9e);
                    end
                end
              reg3388 <= {$signed(($signed(reg3309) > (forvar3362 ?
                      (8'hb7) : reg3292)))};
              if ({$unsigned(reg3293[(3'h4):(1'h1)])})
                begin
                  for (forvar3389 = (1'h0); (forvar3389 < (2'h2)); forvar3389 = (forvar3389 + (1'h1)))
                    begin
                      reg3390 <= (reg3267 + reg3305[(2'h3):(1'h1)]);
                    end
                  if ({reg3333[(3'h4):(3'h4)]})
                    begin
                      reg3391 <= reg3352;
                    end
                  else
                    begin
                      reg3391 <= $signed($unsigned($signed(forvar3329[(1'h0):(1'h0)])));
                      reg3392 <= forvar3343[(3'h7):(3'h6)];
                      reg3393 <= ($signed(forvar3380) ^ reg3234);
                    end
                end
              else
                begin
                  for (forvar3389 = (1'h0); (forvar3389 < (2'h2)); forvar3389 = (forvar3389 + (1'h1)))
                    begin
                      reg3390 <= ($signed(forvar3231) ?
                          {((~forvar3342) ?
                                  (&(8'hb2)) : reg3379)} : (~(^{reg3352})));
                    end
                  reg3391 <= $unsigned(reg3272);
                  reg3392 <= (wire3226 <= forvar3341);
                  if ($signed(reg3380[(4'hb):(1'h0)]))
                    begin
                      reg3393 <= (^({(8'ha9)} ?
                          forvar3324[(1'h1):(1'h0)] : (forvar3231[(3'h6):(3'h4)] ?
                              {(8'had)} : $unsigned(forvar3311))));
                      reg3394 <= $signed($unsigned((reg3326 ?
                          {reg3298} : reg3329[(1'h1):(1'h0)])));
                      reg3395 <= reg3333;
                    end
                  else
                    begin
                      reg3393 <= (|(8'haf));
                      reg3394 <= ({reg3237} ?
                          {((forvar3341 ? (8'hb8) : forvar3321) - (reg3301 ?
                                  reg3258 : forvar3336))} : reg3238);
                    end
                end
              for (forvar3396 = (1'h0); (forvar3396 < (2'h3)); forvar3396 = (forvar3396 + (1'h1)))
                begin
                  if (($signed({(reg3331 ?
                          reg3344 : forvar3263)}) | reg3233[(3'h5):(2'h2)]))
                    begin
                      reg3397 <= reg3239;
                    end
                  else
                    begin
                      reg3397 <= ({$unsigned((reg3353 == reg3391))} || reg3385[(2'h2):(2'h2)]);
                      reg3398 <= (reg3291[(3'h5):(1'h0)] >> reg3374[(2'h2):(2'h2)]);
                    end
                end
            end
        end
    end
  assign wire3399 = $unsigned(reg3363[(2'h3):(2'h3)]);
  assign wire3400 = ((8'ha1) != wire3224[(2'h3):(2'h3)]);
  assign wire3401 = reg3390[(2'h2):(1'h1)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module226
#(parameter param491 = (^~((^{(8'hb2)}) ? ({(8'hb5)} ? ((8'hb3) << (8'hb9)) : ((8'hac) ? (8'ha4) : (8'hba))) : ((^(8'h9e)) << ((8'ha1) - (8'ha0))))))
(y, clk, wire231, wire230, wire229, wire228, wire227);
  output wire [(32'hbbb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire231;
  input wire signed [(3'h7):(1'h0)] wire230;
  input wire [(4'hb):(1'h0)] wire229;
  input wire [(2'h2):(1'h0)] wire228;
  input wire signed [(4'h8):(1'h0)] wire227;
  wire signed [(3'h5):(1'h0)] wire490;
  wire signed [(4'hb):(1'h0)] wire489;
  wire [(4'hd):(1'h0)] wire488;
  wire signed [(3'h5):(1'h0)] wire349;
  wire [(4'he):(1'h0)] wire348;
  wire [(3'h5):(1'h0)] wire347;
  wire [(2'h3):(1'h0)] wire346;
  wire signed [(4'hf):(1'h0)] wire234;
  wire [(4'hb):(1'h0)] wire233;
  wire [(5'h10):(1'h0)] wire232;
  reg signed [(4'he):(1'h0)] reg471 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg483 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg478 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg487 = (1'h0);
  reg [(4'h9):(1'h0)] reg486 = (1'h0);
  reg [(5'h10):(1'h0)] reg485 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg484 = (1'h0);
  reg [(3'h7):(1'h0)] reg482 = (1'h0);
  reg signed [(4'he):(1'h0)] reg481 = (1'h0);
  reg [(4'hc):(1'h0)] reg480 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg479 = (1'h0);
  reg [(3'h6):(1'h0)] reg470 = (1'h0);
  reg [(3'h4):(1'h0)] reg477 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg476 = (1'h0);
  reg [(4'hc):(1'h0)] reg475 = (1'h0);
  reg [(4'hc):(1'h0)] reg473 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg472 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg457 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg445 = (1'h0);
  reg [(4'h8):(1'h0)] reg442 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg469 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg468 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg467 = (1'h0);
  reg [(3'h7):(1'h0)] reg466 = (1'h0);
  reg [(4'h9):(1'h0)] reg465 = (1'h0);
  reg [(4'hd):(1'h0)] reg464 = (1'h0);
  reg [(3'h4):(1'h0)] reg463 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg462 = (1'h0);
  reg [(5'h10):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg460 = (1'h0);
  reg [(5'h10):(1'h0)] reg459 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg458 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg455 = (1'h0);
  reg [(4'hd):(1'h0)] reg454 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg453 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg452 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg451 = (1'h0);
  reg [(3'h7):(1'h0)] reg450 = (1'h0);
  reg [(3'h7):(1'h0)] reg449 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg448 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg447 = (1'h0);
  reg [(4'hf):(1'h0)] reg446 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg444 = (1'h0);
  reg [(3'h7):(1'h0)] reg443 = (1'h0);
  reg [(4'ha):(1'h0)] reg441 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg440 = (1'h0);
  reg signed [(4'he):(1'h0)] reg439 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg438 = (1'h0);
  reg [(4'hc):(1'h0)] reg437 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg436 = (1'h0);
  reg [(4'hc):(1'h0)] reg435 = (1'h0);
  reg [(4'h8):(1'h0)] reg434 = (1'h0);
  reg [(3'h5):(1'h0)] reg433 = (1'h0);
  reg [(2'h3):(1'h0)] reg432 = (1'h0);
  reg [(4'he):(1'h0)] reg431 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg428 = (1'h0);
  reg [(4'ha):(1'h0)] reg427 = (1'h0);
  reg [(4'hd):(1'h0)] reg426 = (1'h0);
  reg [(4'he):(1'h0)] reg424 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg423 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg422 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg420 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg419 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg418 = (1'h0);
  reg [(4'h9):(1'h0)] reg417 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg416 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg415 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg414 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg413 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg412 = (1'h0);
  reg [(5'h10):(1'h0)] reg411 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg410 = (1'h0);
  reg [(4'hf):(1'h0)] reg409 = (1'h0);
  reg [(3'h5):(1'h0)] reg408 = (1'h0);
  reg [(4'hf):(1'h0)] reg406 = (1'h0);
  reg [(4'hd):(1'h0)] reg403 = (1'h0);
  reg [(2'h3):(1'h0)] reg388 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg376 = (1'h0);
  reg [(3'h6):(1'h0)] reg373 = (1'h0);
  reg [(4'he):(1'h0)] reg370 = (1'h0);
  reg [(3'h5):(1'h0)] reg366 = (1'h0);
  reg [(4'he):(1'h0)] reg365 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg360 = (1'h0);
  reg [(3'h7):(1'h0)] reg350 = (1'h0);
  reg [(2'h3):(1'h0)] reg402 = (1'h0);
  reg [(4'hd):(1'h0)] reg401 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg400 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg399 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg397 = (1'h0);
  reg [(4'hd):(1'h0)] reg396 = (1'h0);
  reg [(4'he):(1'h0)] reg395 = (1'h0);
  reg signed [(4'he):(1'h0)] reg394 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg392 = (1'h0);
  reg [(4'ha):(1'h0)] reg391 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg390 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg389 = (1'h0);
  reg [(5'h10):(1'h0)] reg381 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg387 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg386 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg385 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg384 = (1'h0);
  reg [(5'h10):(1'h0)] reg383 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg382 = (1'h0);
  reg [(4'he):(1'h0)] reg380 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg378 = (1'h0);
  reg [(4'hc):(1'h0)] reg377 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg375 = (1'h0);
  reg [(4'hf):(1'h0)] reg374 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg372 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg371 = (1'h0);
  reg [(4'hb):(1'h0)] reg369 = (1'h0);
  reg [(4'hc):(1'h0)] reg368 = (1'h0);
  reg [(4'hd):(1'h0)] reg367 = (1'h0);
  reg [(4'h8):(1'h0)] reg364 = (1'h0);
  reg [(3'h7):(1'h0)] reg363 = (1'h0);
  reg [(4'hf):(1'h0)] reg362 = (1'h0);
  reg [(2'h3):(1'h0)] reg361 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg359 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg358 = (1'h0);
  reg signed [(4'he):(1'h0)] reg357 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg356 = (1'h0);
  reg [(4'hf):(1'h0)] reg355 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg354 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg353 = (1'h0);
  reg [(4'hc):(1'h0)] reg352 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg345 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg344 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg343 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg342 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg340 = (1'h0);
  reg [(4'hb):(1'h0)] reg339 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg338 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg337 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg336 = (1'h0);
  reg [(4'h9):(1'h0)] reg335 = (1'h0);
  reg [(4'hd):(1'h0)] reg334 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg333 = (1'h0);
  reg [(2'h2):(1'h0)] reg332 = (1'h0);
  reg [(4'he):(1'h0)] reg330 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg329 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg328 = (1'h0);
  reg [(4'he):(1'h0)] reg327 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg326 = (1'h0);
  reg signed [(4'he):(1'h0)] reg325 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg317 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg323 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg322 = (1'h0);
  reg [(4'he):(1'h0)] reg321 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg320 = (1'h0);
  reg [(2'h3):(1'h0)] reg319 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg318 = (1'h0);
  reg signed [(4'he):(1'h0)] reg262 = (1'h0);
  reg [(3'h5):(1'h0)] reg311 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg307 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg304 = (1'h0);
  reg [(4'he):(1'h0)] reg315 = (1'h0);
  reg [(4'hf):(1'h0)] reg314 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg313 = (1'h0);
  reg [(4'h9):(1'h0)] reg312 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg310 = (1'h0);
  reg [(2'h3):(1'h0)] reg309 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg308 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg306 = (1'h0);
  reg [(3'h6):(1'h0)] reg303 = (1'h0);
  reg [(3'h5):(1'h0)] reg302 = (1'h0);
  reg [(2'h2):(1'h0)] reg301 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg300 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg299 = (1'h0);
  reg [(4'ha):(1'h0)] reg298 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg297 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg294 = (1'h0);
  reg [(4'h8):(1'h0)] reg293 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg291 = (1'h0);
  reg [(4'hd):(1'h0)] reg290 = (1'h0);
  reg [(4'h9):(1'h0)] reg289 = (1'h0);
  reg [(3'h4):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg285 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg283 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg282 = (1'h0);
  reg [(2'h2):(1'h0)] reg281 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg280 = (1'h0);
  reg signed [(4'he):(1'h0)] reg278 = (1'h0);
  reg [(2'h2):(1'h0)] reg277 = (1'h0);
  reg [(3'h7):(1'h0)] reg276 = (1'h0);
  reg [(4'he):(1'h0)] reg275 = (1'h0);
  reg [(2'h3):(1'h0)] reg274 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg273 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg272 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg271 = (1'h0);
  reg [(2'h3):(1'h0)] reg270 = (1'h0);
  reg [(2'h3):(1'h0)] reg269 = (1'h0);
  reg [(3'h5):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg267 = (1'h0);
  reg [(3'h6):(1'h0)] reg235 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg247 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg236 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg265 = (1'h0);
  reg [(4'hc):(1'h0)] reg264 = (1'h0);
  reg [(4'h8):(1'h0)] reg263 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg261 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg260 = (1'h0);
  reg [(4'he):(1'h0)] reg259 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg258 = (1'h0);
  reg [(3'h7):(1'h0)] reg257 = (1'h0);
  reg [(4'hc):(1'h0)] reg256 = (1'h0);
  reg [(4'h8):(1'h0)] reg255 = (1'h0);
  reg [(4'he):(1'h0)] reg254 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg253 = (1'h0);
  reg [(3'h4):(1'h0)] reg252 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg250 = (1'h0);
  reg [(4'hf):(1'h0)] reg249 = (1'h0);
  reg [(5'h10):(1'h0)] reg248 = (1'h0);
  reg [(3'h6):(1'h0)] reg246 = (1'h0);
  reg [(3'h5):(1'h0)] reg245 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg244 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg243 = (1'h0);
  reg [(5'h10):(1'h0)] reg242 = (1'h0);
  reg [(4'ha):(1'h0)] reg241 = (1'h0);
  reg [(4'hf):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg239 = (1'h0);
  reg [(4'hf):(1'h0)] reg238 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg237 = (1'h0);
  reg [(2'h2):(1'h0)] forvar452 = (1'h0);
  reg [(5'h10):(1'h0)] forvar448 = (1'h0);
  reg [(4'ha):(1'h0)] forvar444 = (1'h0);
  reg [(3'h5):(1'h0)] forvar481 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar484 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar482 = (1'h0);
  reg [(4'ha):(1'h0)] forvar483 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar478 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar474 = (1'h0);
  reg [(4'hb):(1'h0)] forvar471 = (1'h0);
  reg [(4'h8):(1'h0)] forvar470 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar466 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar465 = (1'h0);
  reg [(2'h2):(1'h0)] forvar463 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar459 = (1'h0);
  reg [(5'h10):(1'h0)] forvar455 = (1'h0);
  reg [(3'h5):(1'h0)] forvar443 = (1'h0);
  reg [(4'hd):(1'h0)] forvar447 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar450 = (1'h0);
  reg [(5'h10):(1'h0)] forvar457 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar445 = (1'h0);
  reg [(4'hc):(1'h0)] forvar442 = (1'h0);
  reg [(4'hd):(1'h0)] forvar430 = (1'h0);
  reg [(4'hf):(1'h0)] forvar429 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar425 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar421 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar407 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar405 = (1'h0);
  reg [(4'h8):(1'h0)] forvar404 = (1'h0);
  reg [(2'h2):(1'h0)] forvar384 = (1'h0);
  reg [(4'h9):(1'h0)] forvar374 = (1'h0);
  reg [(4'hb):(1'h0)] forvar368 = (1'h0);
  reg [(4'hb):(1'h0)] forvar367 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar359 = (1'h0);
  reg [(3'h7):(1'h0)] forvar358 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar353 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar352 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar398 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar393 = (1'h0);
  reg [(2'h3):(1'h0)] forvar388 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar385 = (1'h0);
  reg [(2'h2):(1'h0)] forvar382 = (1'h0);
  reg [(4'hb):(1'h0)] forvar381 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar379 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar376 = (1'h0);
  reg [(2'h3):(1'h0)] forvar373 = (1'h0);
  reg [(4'hb):(1'h0)] forvar370 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar366 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar365 = (1'h0);
  reg [(4'h9):(1'h0)] forvar360 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar351 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar350 = (1'h0);
  reg [(4'hd):(1'h0)] forvar341 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar331 = (1'h0);
  reg [(4'h8):(1'h0)] forvar324 = (1'h0);
  reg [(3'h5):(1'h0)] forvar321 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar317 = (1'h0);
  reg [(4'h8):(1'h0)] forvar316 = (1'h0);
  reg [(4'hc):(1'h0)] forvar258 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar252 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar248 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar237 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar238 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar308 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar306 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar311 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar307 = (1'h0);
  reg [(5'h10):(1'h0)] forvar305 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar304 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar296 = (1'h0);
  reg [(4'hf):(1'h0)] forvar295 = (1'h0);
  reg [(4'hf):(1'h0)] forvar292 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar288 = (1'h0);
  reg [(3'h4):(1'h0)] forvar286 = (1'h0);
  reg [(3'h4):(1'h0)] forvar279 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar271 = (1'h0);
  reg [(4'h9):(1'h0)] forvar267 = (1'h0);
  reg [(4'ha):(1'h0)] forvar266 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar244 = (1'h0);
  reg [(5'h10):(1'h0)] forvar262 = (1'h0);
  reg [(3'h7):(1'h0)] forvar251 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar247 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar236 = (1'h0);
  reg [(3'h5):(1'h0)] forvar235 = (1'h0);
  assign y = {wire490,
                 wire489,
                 wire488,
                 wire349,
                 wire348,
                 wire347,
                 wire346,
                 wire234,
                 wire233,
                 wire232,
                 reg471,
                 reg483,
                 reg478,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg482,
                 reg481,
                 reg480,
                 reg479,
                 reg470,
                 reg477,
                 reg476,
                 reg475,
                 reg473,
                 reg472,
                 reg457,
                 reg445,
                 reg442,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 reg447,
                 reg446,
                 reg444,
                 reg443,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 reg428,
                 reg427,
                 reg426,
                 reg424,
                 reg423,
                 reg422,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg406,
                 reg403,
                 reg388,
                 reg376,
                 reg373,
                 reg370,
                 reg366,
                 reg365,
                 reg360,
                 reg350,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg381,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg380,
                 reg378,
                 reg377,
                 reg375,
                 reg374,
                 reg372,
                 reg371,
                 reg369,
                 reg368,
                 reg367,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg317,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg262,
                 reg311,
                 reg307,
                 reg304,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg310,
                 reg309,
                 reg308,
                 reg306,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg294,
                 reg293,
                 reg291,
                 reg290,
                 reg289,
                 reg287,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg235,
                 reg247,
                 reg236,
                 reg265,
                 reg264,
                 reg263,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg250,
                 reg249,
                 reg248,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 forvar452,
                 forvar448,
                 forvar444,
                 forvar481,
                 forvar484,
                 forvar482,
                 forvar483,
                 forvar478,
                 forvar474,
                 forvar471,
                 forvar470,
                 forvar466,
                 forvar465,
                 forvar463,
                 forvar459,
                 forvar455,
                 forvar443,
                 forvar447,
                 forvar450,
                 forvar457,
                 forvar445,
                 forvar442,
                 forvar430,
                 forvar429,
                 forvar425,
                 forvar421,
                 forvar407,
                 forvar405,
                 forvar404,
                 forvar384,
                 forvar374,
                 forvar368,
                 forvar367,
                 forvar359,
                 forvar358,
                 forvar353,
                 forvar352,
                 forvar398,
                 forvar393,
                 forvar388,
                 forvar385,
                 forvar382,
                 forvar381,
                 forvar379,
                 forvar376,
                 forvar373,
                 forvar370,
                 forvar366,
                 forvar365,
                 forvar360,
                 forvar351,
                 forvar350,
                 forvar341,
                 forvar331,
                 forvar324,
                 forvar321,
                 forvar317,
                 forvar316,
                 forvar258,
                 forvar252,
                 forvar248,
                 forvar237,
                 forvar238,
                 forvar308,
                 forvar306,
                 forvar311,
                 forvar307,
                 forvar305,
                 forvar304,
                 forvar296,
                 forvar295,
                 forvar292,
                 forvar288,
                 forvar286,
                 forvar279,
                 forvar271,
                 forvar267,
                 forvar266,
                 forvar244,
                 forvar262,
                 forvar251,
                 forvar247,
                 forvar236,
                 forvar235,
                 (1'h0)};
  assign wire232 = wire227;
  assign wire233 = {wire227[(2'h2):(2'h2)]};
  assign wire234 = ({(~^wire229)} ?
                       (({wire232} & wire229) >= ((^~wire227) ^ wire229[(4'hb):(2'h2)])) : wire227);
  always
    @(posedge clk) begin
      if ($signed(wire230[(2'h3):(1'h1)]))
        begin
          if (wire232)
            begin
              for (forvar235 = (1'h0); (forvar235 < (1'h1)); forvar235 = (forvar235 + (1'h1)))
                begin
                  for (forvar236 = (1'h0); (forvar236 < (2'h3)); forvar236 = (forvar236 + (1'h1)))
                    begin
                      reg237 <= wire232;
                      reg238 <= $signed(wire228[(1'h0):(1'h0)]);
                    end
                  if (reg237)
                    begin
                      reg239 <= (($unsigned($signed(wire227)) ?
                              (~&reg237) : $signed(forvar235[(1'h1):(1'h1)])) ?
                          ($signed($unsigned(wire232)) < wire227) : {$signed($unsigned(reg237))});
                      reg240 <= (~&forvar236);
                      reg241 <= ($unsigned({wire227[(4'h8):(3'h6)]}) ?
                          $signed($signed($unsigned(wire228))) : $signed({(^wire228)}));
                    end
                  else
                    begin
                      reg239 <= forvar236;
                      reg240 <= $signed($unsigned((8'ha8)));
                      reg241 <= (~|($unsigned(reg241[(2'h2):(1'h1)]) & $unsigned(((8'ha3) - reg239))));
                      reg242 <= $unsigned($unsigned(($unsigned(wire234) >>> wire227)));
                    end
                  if (forvar236[(3'h6):(3'h6)])
                    begin
                      reg243 <= $signed(reg238[(3'h6):(2'h2)]);
                      reg244 <= $signed(forvar236[(4'h8):(3'h6)]);
                      reg245 <= (wire233[(3'h4):(2'h3)] == wire234[(3'h6):(1'h0)]);
                      reg246 <= (($unsigned({forvar235}) ?
                          $signed((^(8'hb5))) : reg240) & $unsigned($signed($unsigned(wire228))));
                    end
                  else
                    begin
                      reg243 <= reg245[(1'h1):(1'h0)];
                    end
                end
              for (forvar247 = (1'h0); (forvar247 < (2'h2)); forvar247 = (forvar247 + (1'h1)))
                begin
                  if ({(^~((wire231 && reg239) >= $signed(reg238)))})
                    begin
                      reg248 <= (~^reg240);
                      reg249 <= wire233;
                    end
                  else
                    begin
                      reg248 <= $unsigned((8'ha2));
                      reg249 <= ((~|reg245) >>> (8'hb7));
                      reg250 <= $unsigned($unsigned((~$unsigned(forvar247))));
                    end
                end
              for (forvar251 = (1'h0); (forvar251 < (2'h2)); forvar251 = (forvar251 + (1'h1)))
                begin
                  reg252 <= wire229[(4'ha):(3'h4)];
                  if ((wire228 < (~&reg245)))
                    begin
                      reg253 <= $unsigned((((~wire232) ?
                          (8'ha6) : {reg242}) - {$unsigned(forvar251)}));
                      reg254 <= ($unsigned(((wire231 ? (8'ha5) : reg249) ?
                              $signed(reg249) : (wire229 ? reg248 : reg239))) ?
                          {(-(|forvar236))} : (&$unsigned($unsigned(forvar247))));
                      reg255 <= ($signed({(reg246 ?
                              reg238 : reg249)}) * (-$unsigned(forvar251)));
                      reg256 <= reg250;
                    end
                  else
                    begin
                      reg253 <= reg243;
                    end
                end
              if ((&$signed($unsigned((wire234 >> reg246)))))
                begin
                  reg257 <= reg246[(1'h0):(1'h0)];
                end
              else
                begin
                  reg257 <= reg250[(4'h8):(3'h4)];
                  if ((!wire230[(3'h4):(1'h0)]))
                    begin
                      reg258 <= wire227;
                      reg259 <= (!reg243[(1'h1):(1'h0)]);
                      reg260 <= {reg255[(4'h8):(1'h1)]};
                      reg261 <= reg250[(4'h8):(2'h2)];
                    end
                  else
                    begin
                      reg258 <= $signed(reg239);
                      reg259 <= {reg260};
                      reg260 <= (({reg243[(1'h1):(1'h1)]} >= reg246[(2'h3):(2'h3)]) * $unsigned($signed($unsigned(wire228))));
                      reg261 <= wire230[(3'h6):(2'h3)];
                    end
                  for (forvar262 = (1'h0); (forvar262 < (2'h3)); forvar262 = (forvar262 + (1'h1)))
                    begin
                      reg263 <= (~($unsigned((forvar262 || reg244)) ?
                          (wire228[(1'h1):(1'h1)] ?
                              $signed(reg243) : $signed(reg243)) : $unsigned((~&wire227))));
                      reg264 <= ((!(reg260[(3'h4):(2'h3)] ?
                              wire227[(3'h5):(1'h1)] : (reg248 & forvar236))) ?
                          $signed(((reg249 ?
                              wire227 : reg241) - (^~wire228))) : wire230);
                      reg265 <= ($unsigned(reg239[(4'ha):(2'h3)]) + $unsigned($unsigned($unsigned(reg239))));
                    end
                end
            end
          else
            begin
              if ($unsigned((~^(reg243[(2'h3):(1'h1)] ?
                  (wire228 ? reg242 : reg260) : $unsigned((8'ha8))))))
                begin
                  for (forvar235 = (1'h0); (forvar235 < (1'h0)); forvar235 = (forvar235 + (1'h1)))
                    begin
                      reg236 <= $unsigned($unsigned((8'ha1)));
                      reg237 <= ($signed((8'hb8)) > {wire232[(5'h10):(1'h0)]});
                      reg238 <= $unsigned($unsigned(reg245));
                      reg239 <= (reg261 ^~ reg265);
                    end
                  if ((($signed(forvar236[(3'h6):(2'h3)]) > $signed((-(8'ha2)))) ?
                      ({(^~wire231)} ?
                          ((reg237 ? forvar247 : (8'hb0)) ?
                              $unsigned(wire230) : (reg259 != reg245)) : $signed(wire232)) : forvar236[(3'h7):(3'h6)]))
                    begin
                      reg240 <= {$signed($signed($signed((8'hab))))};
                      reg241 <= $signed($unsigned((8'ha2)));
                      reg242 <= reg263[(3'h5):(1'h0)];
                      reg243 <= (|wire227);
                    end
                  else
                    begin
                      reg240 <= ($unsigned((reg252 ?
                              $unsigned(reg259) : reg264[(1'h1):(1'h0)])) ?
                          forvar247[(4'h8):(3'h5)] : $unsigned(($unsigned(reg258) ?
                              (forvar235 ? wire232 : reg248) : (+wire229))));
                    end
                  for (forvar244 = (1'h0); (forvar244 < (1'h1)); forvar244 = (forvar244 + (1'h1)))
                    begin
                      reg245 <= reg265[(3'h7):(2'h2)];
                      reg246 <= $signed(({forvar244[(1'h0):(1'h0)]} ?
                          ($signed((8'ha3)) | reg236[(4'h8):(3'h6)]) : ($signed(reg252) & (reg264 <= reg248))));
                      reg247 <= $unsigned((~|((reg245 && reg265) == (wire231 ?
                          wire230 : reg264))));
                    end
                end
              else
                begin
                  if ($unsigned($signed({(reg248 ^ (8'h9e))})))
                    begin
                      reg235 <= $unsigned(wire233);
                      reg236 <= $signed(forvar244);
                      reg237 <= $unsigned((reg238 + {$signed(wire232)}));
                    end
                  else
                    begin
                      reg235 <= $unsigned(($unsigned((&wire233)) ?
                          $signed((wire228 ?
                              reg245 : reg245)) : (~^$unsigned(forvar247))));
                      reg236 <= (~^(^((|reg239) ^~ $unsigned(wire228))));
                      reg237 <= ((|$signed({(8'hba)})) >= (reg257[(1'h0):(1'h0)] ?
                          $unsigned($unsigned(reg258)) : $unsigned((wire233 < forvar244))));
                    end
                end
            end
          for (forvar266 = (1'h0); (forvar266 < (1'h0)); forvar266 = (forvar266 + (1'h1)))
            begin
              if (reg248)
                begin
                  if (reg253)
                    begin
                      reg267 <= (8'ha9);
                      reg268 <= {(($signed(reg242) && $unsigned(forvar247)) - {$unsigned(wire234)})};
                      reg269 <= wire228;
                      reg270 <= ((wire227[(3'h5):(1'h0)] <<< $signed(reg263[(2'h2):(2'h2)])) ?
                          reg240 : reg241[(3'h5):(2'h2)]);
                    end
                  else
                    begin
                      reg267 <= reg245;
                      reg268 <= wire227;
                    end
                  if (reg259[(4'h9):(3'h4)])
                    begin
                      reg271 <= $signed(reg270);
                      reg272 <= reg244[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg271 <= $signed((~(reg269 >> $unsigned(wire232))));
                      reg272 <= ($signed((~|reg255[(2'h2):(1'h1)])) ?
                          (&((forvar236 ? reg271 : reg259) ?
                              reg242 : $unsigned(reg242))) : $signed($signed((~|wire232))));
                      reg273 <= {reg252};
                      reg274 <= {{forvar266}};
                    end
                  if (((((~^reg263) ?
                          (reg235 ?
                              wire234 : reg246) : reg244[(4'h9):(4'h9)]) >> $signed(((8'hb3) ?
                          forvar235 : reg264))) ?
                      (&$unsigned((wire230 >> reg268))) : $unsigned(forvar247)))
                    begin
                      reg275 <= $unsigned(($signed($signed(reg254)) * ($signed(reg246) < {forvar247})));
                    end
                  else
                    begin
                      reg275 <= $signed($unsigned((&(reg255 ?
                          forvar236 : wire232))));
                    end
                  if ($unsigned((+{((8'hab) ? (8'ha1) : (8'hb6))})))
                    begin
                      reg276 <= reg275[(4'hd):(4'ha)];
                    end
                  else
                    begin
                      reg276 <= wire228[(1'h1):(1'h0)];
                      reg277 <= $unsigned($unsigned((~^{(8'h9e)})));
                      reg278 <= ((^~reg261[(4'hb):(4'hb)]) < (reg257[(1'h0):(1'h0)] ?
                          (-reg246[(2'h2):(2'h2)]) : forvar266[(3'h5):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar267 = (1'h0); (forvar267 < (1'h1)); forvar267 = (forvar267 + (1'h1)))
                    begin
                      reg268 <= $unsigned($signed((((8'hb1) < reg237) && {reg276})));
                      reg269 <= forvar247[(4'hb):(2'h3)];
                    end
                  reg270 <= reg273[(4'h8):(3'h5)];
                  for (forvar271 = (1'h0); (forvar271 < (1'h1)); forvar271 = (forvar271 + (1'h1)))
                    begin
                      reg272 <= $signed((^~(-reg263)));
                      reg273 <= $signed(reg241);
                      reg274 <= (-((^~reg246[(3'h6):(3'h5)]) ?
                          reg239 : ((reg276 | reg277) ^ wire228[(1'h0):(1'h0)])));
                      reg275 <= (|$unsigned(((^~reg239) ?
                          {(8'hb3)} : $signed(reg277))));
                    end
                  reg276 <= forvar235[(2'h3):(1'h0)];
                end
              for (forvar279 = (1'h0); (forvar279 < (2'h2)); forvar279 = (forvar279 + (1'h1)))
                begin
                  if ($signed((^((&(8'ha3)) ?
                      reg236[(3'h6):(3'h5)] : $signed((8'h9e))))))
                    begin
                      reg280 <= ((&$signed((~|reg264))) ?
                          forvar279 : $signed($signed((^reg238))));
                      reg281 <= (-(^~forvar271));
                    end
                  else
                    begin
                      reg280 <= (reg235[(3'h4):(2'h3)] ?
                          ((8'ha0) ?
                              forvar235[(3'h5):(3'h4)] : $signed($unsigned((8'ha3)))) : ((forvar266 ?
                                  (reg256 >= wire230) : {reg235}) ?
                              ((~reg273) != $signed(reg271)) : $unsigned(forvar236[(4'h9):(3'h6)])));
                    end
                  if ($unsigned((!reg280[(4'ha):(3'h4)])))
                    begin
                      reg282 <= (~^{{(reg273 ? reg275 : (8'ha4))}});
                      reg283 <= ((&{reg274[(1'h0):(1'h0)]}) ?
                          $signed((8'h9f)) : $unsigned(reg238[(4'h9):(2'h2)]));
                      reg284 <= ((^((8'hb5) ?
                              reg254[(3'h7):(2'h3)] : wire233[(4'hb):(2'h3)])) ?
                          $signed(forvar247) : (~|(reg264[(4'hc):(3'h6)] ?
                              $signed(reg246) : ((8'hba) ? reg276 : wire228))));
                      reg285 <= reg281[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg282 <= $unsigned(reg236[(4'hb):(4'h8)]);
                      reg283 <= reg242;
                    end
                  for (forvar286 = (1'h0); (forvar286 < (2'h2)); forvar286 = (forvar286 + (1'h1)))
                    begin
                      reg287 <= reg276[(2'h3):(2'h2)];
                    end
                end
              for (forvar288 = (1'h0); (forvar288 < (2'h3)); forvar288 = (forvar288 + (1'h1)))
                begin
                  if (reg241[(1'h0):(1'h0)])
                    begin
                      reg289 <= reg250;
                    end
                  else
                    begin
                      reg289 <= ($signed((8'hae)) ?
                          ($signed(reg250[(1'h0):(1'h0)]) ?
                              (~reg249[(4'hd):(1'h1)]) : $unsigned(forvar266[(4'h8):(4'h8)])) : reg246);
                      reg290 <= (|reg285[(3'h4):(2'h3)]);
                      reg291 <= ($unsigned({reg235[(1'h1):(1'h1)]}) ?
                          $unsigned($signed(reg247[(3'h5):(1'h0)])) : reg245);
                    end
                  for (forvar292 = (1'h0); (forvar292 < (2'h3)); forvar292 = (forvar292 + (1'h1)))
                    begin
                      reg293 <= $signed({$signed(reg247)});
                    end
                  reg294 <= (reg264[(2'h3):(1'h0)] ?
                      (^~forvar244) : ($signed(reg293) ?
                          ((^~reg275) && wire227[(2'h3):(2'h2)]) : (((8'haa) >>> reg287) ^ (~&reg264))));
                end
              for (forvar295 = (1'h0); (forvar295 < (2'h3)); forvar295 = (forvar295 + (1'h1)))
                begin
                  for (forvar296 = (1'h0); (forvar296 < (2'h3)); forvar296 = (forvar296 + (1'h1)))
                    begin
                      reg297 <= reg287;
                      reg298 <= $unsigned(reg297);
                      reg299 <= (&$signed(((reg252 ^~ reg298) ?
                          $unsigned((8'hb1)) : (wire231 && reg240))));
                    end
                  reg300 <= (-reg272);
                  if ((&reg294[(3'h4):(3'h4)]))
                    begin
                      reg301 <= (8'ha2);
                      reg302 <= $signed($unsigned(reg275[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg301 <= ({(&reg259[(4'hb):(4'h8)])} ?
                          $unsigned($unsigned({wire231})) : $signed({forvar279}));
                      reg302 <= (!(-{{reg301}}));
                      reg303 <= (((forvar292 ?
                                  wire230[(3'h5):(1'h0)] : (~&forvar279)) ?
                              (~&(reg258 <<< reg294)) : reg238[(3'h5):(2'h2)]) ?
                          $unsigned({$signed(reg284)}) : reg280[(4'h9):(3'h6)]);
                    end
                end
            end
          if ($signed($unsigned((reg259 ~^ $unsigned(reg269)))))
            begin
              for (forvar304 = (1'h0); (forvar304 < (1'h1)); forvar304 = (forvar304 + (1'h1)))
                begin
                  for (forvar305 = (1'h0); (forvar305 < (2'h2)); forvar305 = (forvar305 + (1'h1)))
                    begin
                      reg306 <= ({$unsigned((forvar236 ?
                              reg261 : forvar267))} + forvar251);
                    end
                  for (forvar307 = (1'h0); (forvar307 < (2'h3)); forvar307 = (forvar307 + (1'h1)))
                    begin
                      reg308 <= (8'hb1);
                    end
                  if ($signed($signed((~^(reg291 - reg287)))))
                    begin
                      reg309 <= reg253;
                    end
                  else
                    begin
                      reg309 <= {(^~(wire232 ^~ (reg267 ? reg273 : reg264)))};
                      reg310 <= forvar236;
                    end
                  for (forvar311 = (1'h0); (forvar311 < (1'h1)); forvar311 = (forvar311 + (1'h1)))
                    begin
                      reg312 <= forvar296[(3'h7):(2'h2)];
                      reg313 <= $signed({reg252[(1'h0):(1'h0)]});
                      reg314 <= (~^reg308);
                      reg315 <= $unsigned(reg310[(1'h1):(1'h0)]);
                    end
                end
            end
          else
            begin
              reg304 <= ((~|{$unsigned((8'hb1))}) < reg293[(4'h8):(3'h5)]);
              for (forvar305 = (1'h0); (forvar305 < (2'h3)); forvar305 = (forvar305 + (1'h1)))
                begin
                  for (forvar306 = (1'h0); (forvar306 < (1'h0)); forvar306 = (forvar306 + (1'h1)))
                    begin
                      reg307 <= ($unsigned(reg264[(3'h5):(1'h0)]) ?
                          $signed($unsigned((~|wire232))) : reg258);
                    end
                  for (forvar308 = (1'h0); (forvar308 < (1'h0)); forvar308 = (forvar308 + (1'h1)))
                    begin
                      reg309 <= reg267[(3'h5):(2'h3)];
                      reg310 <= $signed((&((reg310 ? reg276 : reg307) ?
                          $unsigned(reg299) : $unsigned(reg302))));
                      reg311 <= $signed(((wire230 != $signed(reg304)) ?
                          ((-reg304) ?
                              (reg268 * reg255) : wire230) : {$signed(reg270)}));
                      reg312 <= (($signed(forvar308) ^ {reg299[(1'h1):(1'h0)]}) ?
                          $unsigned(reg307) : reg280[(4'hf):(3'h7)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar235 = (1'h0); (forvar235 < (1'h1)); forvar235 = (forvar235 + (1'h1)))
            begin
              if ((^reg250[(2'h2):(2'h2)]))
                begin
                  if ((reg237[(1'h1):(1'h0)] <<< ($unsigned((reg300 >> reg253)) << ((~|(8'h9d)) ^ reg273[(3'h5):(1'h0)]))))
                    begin
                      reg236 <= $signed(reg264[(4'hc):(4'hb)]);
                      reg237 <= reg264[(4'hc):(1'h1)];
                    end
                  else
                    begin
                      reg236 <= ({$signed(reg270[(1'h1):(1'h1)])} ?
                          $unsigned(forvar244) : (8'haa));
                      reg237 <= ($unsigned((reg276 ?
                              (reg249 ? reg293 : reg248) : {forvar304})) ?
                          (-{(+reg272)}) : forvar308[(1'h1):(1'h0)]);
                    end
                  for (forvar238 = (1'h0); (forvar238 < (1'h0)); forvar238 = (forvar238 + (1'h1)))
                    begin
                      reg239 <= $unsigned((+(^reg237[(3'h4):(3'h4)])));
                      reg240 <= (({(reg303 != (8'hb3))} > reg267[(4'hc):(4'h9)]) ^ (($unsigned(forvar279) ?
                              (reg261 ? reg283 : reg267) : (~^reg302)) ?
                          $signed($signed(forvar244)) : {{reg249}}));
                    end
                end
              else
                begin
                  reg236 <= (~&reg272);
                  for (forvar237 = (1'h0); (forvar237 < (1'h1)); forvar237 = (forvar237 + (1'h1)))
                    begin
                      reg238 <= $signed($unsigned(($unsigned(reg297) + (|(8'hb4)))));
                      reg239 <= reg255[(3'h7):(3'h6)];
                      reg240 <= (-(-$unsigned($signed(reg293))));
                      reg241 <= (((+forvar235) ?
                          ({reg261} ?
                              (reg257 <<< reg275) : (reg272 ^~ forvar288)) : $signed(reg242)) == ((~&reg242[(1'h1):(1'h1)]) ?
                          $unsigned($signed(forvar247)) : {reg301[(1'h0):(1'h0)]}));
                    end
                  if (reg314[(3'h7):(2'h3)])
                    begin
                      reg242 <= ($unsigned((~forvar296)) >>> reg273[(2'h2):(1'h0)]);
                      reg243 <= ((($unsigned(wire227) ?
                          reg301[(2'h2):(2'h2)] : (~forvar238)) << forvar244[(1'h0):(1'h0)]) != (reg293[(3'h7):(3'h6)] <<< reg274));
                      reg244 <= {wire228[(1'h1):(1'h1)]};
                    end
                  else
                    begin
                      reg242 <= (((reg272[(1'h0):(1'h0)] ?
                          (~^reg250) : $signed(forvar311)) || $unsigned($unsigned(forvar292))) < $signed($unsigned({reg274})));
                      reg243 <= (((8'ha6) && wire230) ?
                          $unsigned($signed($signed(reg299))) : $signed(((reg242 ?
                              reg287 : forvar286) >> $signed(reg314))));
                    end
                  if (($unsigned($signed(reg258[(4'hb):(3'h6)])) ?
                      forvar267 : (((&reg255) ?
                              reg268 : (reg240 ? (8'h9c) : (8'hb9))) ?
                          reg280[(1'h0):(1'h0)] : {(8'haf)})))
                    begin
                      reg245 <= ($signed(reg263) ?
                          ($signed((forvar235 ? wire228 : reg255)) ?
                              (&forvar305[(4'hc):(4'h8)]) : (8'haf)) : $unsigned($unsigned((forvar307 ?
                              reg309 : reg289))));
                    end
                  else
                    begin
                      reg245 <= (8'hb0);
                      reg246 <= $unsigned(($unsigned(reg315) < reg265));
                      reg247 <= ((-(~(|forvar235))) || (((reg294 ?
                              (8'hb8) : reg236) ?
                          (reg248 ?
                              reg280 : wire229) : reg310[(3'h5):(1'h0)]) || reg236));
                    end
                end
            end
          if (((({wire233} ? (reg313 >> (8'hba)) : forvar295) ?
                  $unsigned($signed(reg246)) : ((^~reg274) > $signed(reg242))) ?
              $signed(($signed(reg268) ^~ reg293)) : $signed((((8'hb0) | reg269) < $unsigned(forvar236)))))
            begin
              for (forvar248 = (1'h0); (forvar248 < (1'h0)); forvar248 = (forvar248 + (1'h1)))
                begin
                  if ((8'hb7))
                    begin
                      reg249 <= reg255;
                    end
                  else
                    begin
                      reg249 <= reg284[(3'h5):(1'h0)];
                    end
                end
              reg250 <= ((($signed(reg241) ? reg274 : forvar307) ?
                      ($signed((8'hb3)) - $signed(forvar279)) : ((reg304 || (8'hba)) <<< $unsigned(reg274))) ?
                  $unsigned($unsigned((forvar244 * reg307))) : ({forvar236} < ((forvar251 ?
                      reg241 : reg294) <<< $signed(forvar237))));
              for (forvar251 = (1'h0); (forvar251 < (2'h2)); forvar251 = (forvar251 + (1'h1)))
                begin
                  for (forvar252 = (1'h0); (forvar252 < (1'h1)); forvar252 = (forvar252 + (1'h1)))
                    begin
                      reg253 <= (forvar304[(2'h2):(1'h0)] ?
                          $signed($unsigned({reg255})) : $unsigned($unsigned($signed(reg241))));
                      reg254 <= reg291;
                      reg255 <= ({(^reg264)} ?
                          (((&reg269) ? (|forvar267) : (wire231 == reg310)) ?
                              ($unsigned(forvar288) ?
                                  {reg310} : reg283[(4'ha):(3'h5)]) : reg247[(3'h5):(3'h5)]) : wire234);
                      reg256 <= $unsigned($signed({(^~reg244)}));
                    end
                  reg257 <= reg310;
                  for (forvar258 = (1'h0); (forvar258 < (2'h3)); forvar258 = (forvar258 + (1'h1)))
                    begin
                      reg259 <= (~|$signed($unsigned(forvar305)));
                      reg260 <= forvar266[(3'h4):(1'h0)];
                    end
                  if ((forvar236[(3'h4):(3'h4)] * $unsigned(reg282)))
                    begin
                      reg261 <= forvar237;
                      reg262 <= $unsigned(wire230[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg261 <= $signed(((|(&reg270)) >> $signed(reg307)));
                    end
                end
              reg263 <= (~(forvar258 <= forvar251));
            end
          else
            begin
              reg248 <= $unsigned(($signed(forvar296[(3'h6):(2'h3)]) ?
                  $signed((reg309 ?
                      forvar251 : reg287)) : $signed($unsigned((8'hac)))));
            end
        end
      for (forvar316 = (1'h0); (forvar316 < (1'h0)); forvar316 = (forvar316 + (1'h1)))
        begin
          if ($signed(((-$signed(reg298)) * (((8'hae) - reg275) >>> (forvar247 <<< wire230)))))
            begin
              for (forvar317 = (1'h0); (forvar317 < (1'h1)); forvar317 = (forvar317 + (1'h1)))
                begin
                  reg318 <= (($signed((reg313 < reg314)) ?
                      reg263 : $signed(reg302)) - (!forvar311));
                end
              reg319 <= (+reg247);
            end
          else
            begin
              if (reg304)
                begin
                  for (forvar317 = (1'h0); (forvar317 < (1'h0)); forvar317 = (forvar317 + (1'h1)))
                    begin
                      reg318 <= ($signed((~&((8'haa) + reg250))) >> ({reg263} <<< {reg298}));
                      reg319 <= ((^reg271[(4'h9):(3'h7)]) ?
                          $unsigned(((reg311 ?
                              forvar306 : reg249) >>> $signed(reg284))) : (~&({(8'hb5)} < (forvar271 ?
                              forvar308 : forvar235))));
                    end
                  if ({forvar279[(3'h4):(3'h4)]})
                    begin
                      reg320 <= (~|reg291);
                      reg321 <= ({$unsigned(reg243[(3'h4):(2'h2)])} ?
                          (+$signed((forvar236 & reg240))) : (^~($unsigned(reg244) ?
                              (reg249 ?
                                  reg257 : (8'ha7)) : $unsigned(reg258))));
                    end
                  else
                    begin
                      reg320 <= (~&{((wire234 ?
                              forvar266 : (8'haa)) <= (8'hb7))});
                      reg321 <= wire229[(3'h4):(2'h3)];
                    end
                  reg322 <= reg237;
                  reg323 <= $signed((~&($signed(forvar317) >> reg291[(4'hb):(3'h6)])));
                end
              else
                begin
                  if (reg280)
                    begin
                      reg317 <= (~^reg268);
                      reg318 <= $unsigned($signed(((&wire230) ?
                          $signed(forvar244) : $signed(reg241))));
                      reg319 <= reg256;
                      reg320 <= (-(((reg238 + wire228) <= $signed(reg235)) > (-$signed(reg277))));
                    end
                  else
                    begin
                      reg317 <= reg238;
                      reg318 <= $signed(reg297);
                      reg319 <= (((~|$unsigned(reg254)) ^~ reg293[(2'h2):(1'h0)]) ?
                          (^{(!reg307)}) : (((reg311 ^~ reg270) ?
                              (forvar295 ?
                                  reg310 : reg321) : reg235) * reg310));
                      reg320 <= (~|$signed(reg285));
                    end
                  for (forvar321 = (1'h0); (forvar321 < (1'h0)); forvar321 = (forvar321 + (1'h1)))
                    begin
                      reg322 <= (^$unsigned(((forvar311 ?
                          reg236 : forvar266) | $unsigned(forvar252))));
                      reg323 <= {(-$unsigned((+reg297)))};
                    end
                  for (forvar324 = (1'h0); (forvar324 < (1'h1)); forvar324 = (forvar324 + (1'h1)))
                    begin
                      reg325 <= $signed(((~(forvar238 ? (8'h9c) : reg237)) ?
                          {reg306} : (reg243 ~^ {reg278})));
                      reg326 <= ((|$signed(reg272[(2'h2):(1'h0)])) ?
                          reg291[(3'h4):(1'h0)] : (!reg307));
                      reg327 <= $unsigned($signed((reg249[(1'h0):(1'h0)] >= reg252)));
                    end
                  if (forvar244)
                    begin
                      reg328 <= $unsigned(forvar235);
                      reg329 <= (~&(8'hb7));
                      reg330 <= $unsigned($unsigned(forvar306));
                    end
                  else
                    begin
                      reg328 <= reg258[(3'h5):(2'h3)];
                    end
                end
              if ($signed(reg260[(2'h2):(1'h1)]))
                begin
                  for (forvar331 = (1'h0); (forvar331 < (2'h2)); forvar331 = (forvar331 + (1'h1)))
                    begin
                      reg332 <= forvar251;
                    end
                  if ($unsigned(reg299))
                    begin
                      reg333 <= $unsigned(($unsigned($signed(reg278)) << $signed($unsigned((8'hb8)))));
                      reg334 <= (((8'hb4) ?
                          (8'ha4) : {((8'haa) ^~ (8'hac))}) & ($signed({(8'hb0)}) ?
                          (~$signed(wire231)) : ((reg322 - reg238) ?
                              $signed(forvar286) : (^(8'hb0)))));
                    end
                  else
                    begin
                      reg333 <= (~|(~&reg297[(3'h4):(2'h3)]));
                      reg334 <= reg321;
                      reg335 <= ($unsigned(((8'hb9) == $unsigned(reg289))) ?
                          (forvar305 << {(~|reg328)}) : $signed($signed($signed(reg312))));
                      reg336 <= {forvar307};
                    end
                  if (reg334[(3'h5):(2'h2)])
                    begin
                      reg337 <= reg289;
                      reg338 <= {{$unsigned(((8'hb9) - forvar316))}};
                      reg339 <= $signed($unsigned((reg274 ^ (-forvar262))));
                      reg340 <= {reg311};
                    end
                  else
                    begin
                      reg337 <= (~|(&(reg306 & {reg311})));
                      reg338 <= (|{(|(reg249 ? reg254 : forvar295))});
                    end
                  for (forvar341 = (1'h0); (forvar341 < (2'h2)); forvar341 = (forvar341 + (1'h1)))
                    begin
                      reg342 <= $unsigned((+((reg336 ~^ forvar248) ?
                          forvar266 : {reg259})));
                      reg343 <= (&(^~((~^reg269) >> (reg283 ?
                          reg269 : reg281))));
                      reg344 <= (reg343 ?
                          (((!forvar258) ^ reg250[(2'h2):(1'h0)]) ?
                              $unsigned((~reg330)) : $unsigned(forvar266)) : $signed(((forvar288 ?
                                  forvar308 : forvar238) ?
                              (forvar306 - forvar316) : $signed((8'ha2)))));
                    end
                end
              else
                begin
                  for (forvar331 = (1'h0); (forvar331 < (2'h3)); forvar331 = (forvar331 + (1'h1)))
                    begin
                      reg332 <= $signed(reg241);
                      reg333 <= ((~&reg238) ?
                          $unsigned($unsigned((forvar262 ?
                              reg275 : wire230))) : reg330[(4'h8):(2'h3)]);
                      reg334 <= (!reg272[(1'h0):(1'h0)]);
                    end
                end
              reg345 <= (8'had);
            end
        end
    end
  assign wire346 = reg297[(3'h4):(1'h1)];
  assign wire347 = reg293[(1'h1):(1'h1)];
  assign wire348 = (reg312 <<< $signed(reg325));
  assign wire349 = $unsigned($unsigned($signed(reg276[(3'h4):(2'h3)])));
  always
    @(posedge clk) begin
      if ($unsigned((($signed(reg318) ?
          reg325 : {wire232}) * ($unsigned(reg330) ?
          ((8'h9d) || wire230) : (-reg237)))))
        begin
          for (forvar350 = (1'h0); (forvar350 < (1'h0)); forvar350 = (forvar350 + (1'h1)))
            begin
              for (forvar351 = (1'h0); (forvar351 < (1'h0)); forvar351 = (forvar351 + (1'h1)))
                begin
                  if (reg312[(4'h8):(3'h6)])
                    begin
                      reg352 <= (8'h9e);
                      reg353 <= (8'haa);
                    end
                  else
                    begin
                      reg352 <= $unsigned(reg311);
                      reg353 <= $signed((($unsigned(reg290) == $unsigned(reg342)) | $unsigned(reg237)));
                      reg354 <= ($signed((reg330[(4'ha):(3'h7)] ?
                          (reg285 ?
                              reg291 : reg329) : (-reg253))) > reg239[(3'h7):(3'h6)]);
                      reg355 <= (8'ha7);
                    end
                  if (((^~$signed((wire233 ? reg293 : reg311))) >> reg311))
                    begin
                      reg356 <= $signed(reg241[(3'h6):(3'h5)]);
                      reg357 <= {(reg235 ?
                              ($unsigned(reg237) ?
                                  reg321 : (^~wire234)) : $unsigned($unsigned(reg271)))};
                      reg358 <= $unsigned(($unsigned(reg260) <= $signed((reg294 ?
                          (8'haa) : reg240))));
                      reg359 <= ((reg285 ?
                              $unsigned($unsigned(reg301)) : reg245[(2'h3):(1'h0)]) ?
                          ($unsigned($unsigned(wire233)) & (reg353[(2'h2):(1'h1)] + reg258)) : (wire228[(2'h2):(1'h1)] ?
                              $unsigned((reg256 <= reg353)) : {reg241}));
                    end
                  else
                    begin
                      reg356 <= reg309;
                      reg357 <= $signed(reg244[(2'h3):(1'h1)]);
                    end
                  for (forvar360 = (1'h0); (forvar360 < (2'h2)); forvar360 = (forvar360 + (1'h1)))
                    begin
                      reg361 <= {($unsigned($unsigned(reg283)) ?
                              (~|(-wire232)) : $unsigned(((8'hba) <= reg306)))};
                      reg362 <= reg312[(3'h4):(1'h1)];
                      reg363 <= reg260[(4'h9):(2'h3)];
                      reg364 <= $unsigned((&(reg242 ?
                          reg262 : $signed(reg246))));
                    end
                end
              for (forvar365 = (1'h0); (forvar365 < (2'h2)); forvar365 = (forvar365 + (1'h1)))
                begin
                  for (forvar366 = (1'h0); (forvar366 < (2'h2)); forvar366 = (forvar366 + (1'h1)))
                    begin
                      reg367 <= reg245;
                      reg368 <= ({((wire228 ? reg235 : reg362) ?
                                  {reg355} : $signed(forvar365))} ?
                          (((!reg342) ~^ (reg301 + reg359)) ?
                              reg293 : ($unsigned(reg287) ?
                                  (reg364 << reg336) : $signed((8'ha9)))) : (!$signed(reg307)));
                      reg369 <= $unsigned($signed({$unsigned(reg275)}));
                    end
                  for (forvar370 = (1'h0); (forvar370 < (2'h2)); forvar370 = (forvar370 + (1'h1)))
                    begin
                      reg371 <= reg297;
                      reg372 <= forvar350[(3'h6):(2'h3)];
                    end
                  for (forvar373 = (1'h0); (forvar373 < (1'h1)); forvar373 = (forvar373 + (1'h1)))
                    begin
                      reg374 <= reg273[(1'h0):(1'h0)];
                      reg375 <= (~^$signed($unsigned(reg274[(1'h1):(1'h1)])));
                    end
                  for (forvar376 = (1'h0); (forvar376 < (1'h0)); forvar376 = (forvar376 + (1'h1)))
                    begin
                      reg377 <= (~$unsigned((-(~reg246))));
                      reg378 <= $unsigned((~&{{wire346}}));
                    end
                end
            end
          for (forvar379 = (1'h0); (forvar379 < (2'h2)); forvar379 = (forvar379 + (1'h1)))
            begin
              reg380 <= reg297;
              if ({(((+reg328) ?
                      reg369[(4'hb):(2'h3)] : reg335) ~^ (reg254[(4'h9):(4'h9)] ~^ reg306[(1'h0):(1'h0)]))})
                begin
                  for (forvar381 = (1'h0); (forvar381 < (1'h1)); forvar381 = (forvar381 + (1'h1)))
                    begin
                      reg382 <= (8'hb7);
                      reg383 <= $signed(reg238);
                    end
                  if (reg308[(1'h1):(1'h1)])
                    begin
                      reg384 <= (($unsigned((reg303 > wire346)) < reg368[(4'h9):(3'h6)]) ?
                          $signed(reg315[(4'hd):(2'h2)]) : $unsigned(((reg274 ?
                                  reg308 : (8'hb3)) ?
                              reg241[(3'h5):(2'h3)] : (reg243 && reg328))));
                    end
                  else
                    begin
                      reg384 <= (|(((forvar370 <<< reg323) ?
                          reg375 : $signed(reg282)) & {$unsigned(reg375)}));
                      reg385 <= ((8'h9c) || (~^reg281));
                      reg386 <= (forvar360[(4'h8):(2'h3)] >>> forvar379);
                    end
                  reg387 <= $signed((8'ha4));
                end
              else
                begin
                  reg381 <= $signed(forvar381);
                  for (forvar382 = (1'h0); (forvar382 < (2'h3)); forvar382 = (forvar382 + (1'h1)))
                    begin
                      reg383 <= (((^~$unsigned(reg318)) ?
                              (~|reg243) : reg333[(1'h0):(1'h0)]) ?
                          $signed((~|((8'hab) || (8'hb0)))) : wire231[(3'h5):(3'h4)]);
                      reg384 <= (reg326[(4'hc):(4'ha)] ?
                          ((!$signed(reg282)) ?
                              reg235 : (8'ha9)) : $signed((reg241 ?
                              reg330[(4'ha):(2'h2)] : (^reg368))));
                    end
                  for (forvar385 = (1'h0); (forvar385 < (2'h3)); forvar385 = (forvar385 + (1'h1)))
                    begin
                      reg386 <= reg387;
                    end
                end
              for (forvar388 = (1'h0); (forvar388 < (1'h1)); forvar388 = (forvar388 + (1'h1)))
                begin
                  reg389 <= {wire230[(3'h4):(1'h1)]};
                  if ((reg285[(3'h7):(3'h7)] == $unsigned((((8'ha9) < reg339) && (reg362 ?
                      forvar382 : wire232)))))
                    begin
                      reg390 <= reg283[(4'ha):(2'h2)];
                    end
                  else
                    begin
                      reg390 <= ((reg255 > $unsigned($signed((8'h9e)))) | $signed((~|$signed((8'ha9)))));
                      reg391 <= ((^~($unsigned(reg323) ?
                          reg273[(1'h0):(1'h0)] : (8'ha7))) && $signed({reg384[(4'he):(4'he)]}));
                      reg392 <= forvar350[(4'ha):(3'h4)];
                    end
                  for (forvar393 = (1'h0); (forvar393 < (1'h0)); forvar393 = (forvar393 + (1'h1)))
                    begin
                      reg394 <= $signed(reg356[(2'h3):(2'h2)]);
                      reg395 <= (reg369 ?
                          {$signed((~|reg374))} : $signed($unsigned($signed(forvar381))));
                      reg396 <= (8'ha8);
                      reg397 <= reg368;
                    end
                  for (forvar398 = (1'h0); (forvar398 < (2'h2)); forvar398 = (forvar398 + (1'h1)))
                    begin
                      reg399 <= reg317;
                      reg400 <= $unsigned(reg236);
                      reg401 <= {($unsigned({reg280}) & ((forvar398 ^~ reg375) + $unsigned((8'h9c))))};
                      reg402 <= reg241;
                    end
                end
            end
        end
      else
        begin
          reg350 <= ($unsigned($signed((8'hb5))) ?
              {reg299[(1'h1):(1'h1)]} : $unsigned($signed($unsigned(reg275))));
          for (forvar351 = (1'h0); (forvar351 < (1'h0)); forvar351 = (forvar351 + (1'h1)))
            begin
              for (forvar352 = (1'h0); (forvar352 < (2'h2)); forvar352 = (forvar352 + (1'h1)))
                begin
                  for (forvar353 = (1'h0); (forvar353 < (1'h1)); forvar353 = (forvar353 + (1'h1)))
                    begin
                      reg354 <= (^$unsigned({$signed((8'h9d))}));
                      reg355 <= {$unsigned(((^(8'ha2)) <<< $signed(reg378)))};
                      reg356 <= forvar381[(1'h0):(1'h0)];
                    end
                end
              reg357 <= (~&(8'hb2));
            end
          if ($signed((|reg343)))
            begin
              if ($signed({{(+(8'haa))}}))
                begin
                  for (forvar358 = (1'h0); (forvar358 < (1'h0)); forvar358 = (forvar358 + (1'h1)))
                    begin
                      reg359 <= reg371[(4'h9):(3'h6)];
                      reg360 <= (reg276 > $unsigned($signed($unsigned(reg255))));
                      reg361 <= (reg264 || $unsigned($unsigned((8'hb4))));
                    end
                end
              else
                begin
                  if ($signed(($signed((reg261 ^ reg329)) << ((reg313 ~^ reg317) ?
                      $unsigned(reg387) : ((8'h9f) != reg267)))))
                    begin
                      reg358 <= reg237[(1'h1):(1'h0)];
                      reg359 <= (~^({$unsigned(reg307)} <= {reg363[(3'h5):(2'h3)]}));
                    end
                  else
                    begin
                      reg358 <= ($unsigned($unsigned({reg315})) << ($unsigned(forvar376) ?
                          {(reg278 ?
                                  reg391 : reg386)} : $unsigned((forvar358 ^~ reg267))));
                      reg359 <= $signed(({reg236} ?
                          ($unsigned((8'ha9)) + forvar379) : (8'h9d)));
                      reg360 <= $unsigned(reg247[(2'h2):(1'h1)]);
                      reg361 <= $unsigned(reg278);
                    end
                  reg362 <= (($unsigned({(8'h9e)}) ^~ {(wire346 ?
                              forvar365 : reg335)}) ?
                      (reg350[(3'h4):(3'h4)] ?
                          (-{reg262}) : ($signed(reg277) ?
                              (reg237 <= reg254) : (reg308 ?
                                  reg362 : forvar398))) : reg241);
                  if (wire229[(1'h0):(1'h0)])
                    begin
                      reg363 <= $signed($unsigned(reg236[(3'h7):(1'h1)]));
                      reg364 <= ($unsigned(($signed(reg299) ?
                          ((8'h9e) ? reg278 : reg271) : reg361)) >>> reg239);
                      reg365 <= {(^(~|$unsigned(reg285)))};
                    end
                  else
                    begin
                      reg363 <= reg312[(4'h9):(1'h0)];
                      reg364 <= {(8'hba)};
                    end
                  for (forvar366 = (1'h0); (forvar366 < (2'h2)); forvar366 = (forvar366 + (1'h1)))
                    begin
                      reg367 <= $unsigned(reg236);
                      reg368 <= ($unsigned({((8'ha4) <<< reg264)}) ?
                          (((+forvar360) ?
                              $unsigned(reg241) : $signed(reg357)) != (forvar398[(1'h1):(1'h0)] ?
                              reg246[(2'h3):(2'h3)] : $signed(reg328))) : ((reg345 ?
                                  (reg319 ?
                                      (8'hba) : reg238) : $unsigned(reg328)) ?
                              reg368 : $unsigned((forvar352 && forvar376))));
                    end
                end
            end
          else
            begin
              reg358 <= $unsigned(((reg323[(3'h6):(1'h1)] <= (reg278 ?
                  reg371 : reg328)) * reg273[(3'h4):(2'h3)]));
              for (forvar359 = (1'h0); (forvar359 < (2'h2)); forvar359 = (forvar359 + (1'h1)))
                begin
                  if (forvar385)
                    begin
                      reg360 <= (~^(&{$signed(forvar365)}));
                      reg361 <= (reg386 * reg267);
                      reg362 <= reg330[(3'h7):(1'h1)];
                      reg363 <= forvar360;
                    end
                  else
                    begin
                      reg360 <= reg395;
                      reg361 <= $signed(reg253[(1'h0):(1'h0)]);
                      reg362 <= reg387[(1'h1):(1'h0)];
                      reg363 <= reg299[(2'h3):(2'h2)];
                    end
                  if ({((8'ha4) && ((reg290 && forvar388) ?
                          (forvar359 ?
                              reg255 : reg257) : reg306[(3'h5):(2'h3)]))})
                    begin
                      reg364 <= reg321;
                      reg365 <= $signed((((reg241 ?
                              reg320 : reg263) ^ $signed((8'hb5))) ?
                          (~&reg320[(4'h9):(3'h4)]) : (~$signed(forvar350))));
                    end
                  else
                    begin
                      reg364 <= (~^$signed($signed((8'ha0))));
                      reg365 <= (reg386 ?
                          reg262[(4'hc):(2'h3)] : (~^((reg263 ?
                                  (8'hb2) : (8'h9c)) ?
                              $unsigned(forvar350) : (reg342 - forvar373))));
                      reg366 <= $unsigned((($unsigned(reg335) - (~&reg319)) > ((reg282 ?
                              reg262 : (8'h9e)) ?
                          reg263 : {reg333})));
                    end
                end
              for (forvar367 = (1'h0); (forvar367 < (2'h3)); forvar367 = (forvar367 + (1'h1)))
                begin
                  for (forvar368 = (1'h0); (forvar368 < (2'h2)); forvar368 = (forvar368 + (1'h1)))
                    begin
                      reg369 <= ({(^~forvar373[(1'h1):(1'h0)])} >>> (~{((8'hab) <<< reg336)}));
                    end
                  if ((~|reg247))
                    begin
                      reg370 <= $signed(reg367[(1'h1):(1'h1)]);
                      reg371 <= ((((reg395 ? reg344 : forvar351) ?
                          (reg238 ? reg396 : reg259) : {reg396}) ^~ ((reg238 ?
                              reg364 : (8'ha2)) ?
                          (reg322 >>> (8'hb2)) : $unsigned((8'h9e)))) >> reg402);
                    end
                  else
                    begin
                      reg370 <= reg301[(2'h2):(2'h2)];
                      reg371 <= ((((reg321 ~^ reg261) < $signed(reg383)) * $signed({reg285})) * $unsigned($unsigned((8'ha8))));
                      reg372 <= wire346[(1'h1):(1'h0)];
                      reg373 <= {{reg253}};
                    end
                end
              for (forvar374 = (1'h0); (forvar374 < (2'h3)); forvar374 = (forvar374 + (1'h1)))
                begin
                  if ((~|$unsigned($signed(reg256))))
                    begin
                      reg375 <= $signed($signed({(reg382 ? reg385 : reg242)}));
                      reg376 <= $unsigned($signed($unsigned($unsigned((8'hb8)))));
                      reg377 <= {$unsigned((-reg344))};
                      reg378 <= reg339[(4'ha):(1'h1)];
                    end
                  else
                    begin
                      reg375 <= reg271[(4'ha):(4'ha)];
                      reg376 <= reg310[(4'h8):(3'h6)];
                      reg377 <= (&(reg262 - (-(~&wire346))));
                    end
                  for (forvar379 = (1'h0); (forvar379 < (2'h2)); forvar379 = (forvar379 + (1'h1)))
                    begin
                      reg380 <= reg365;
                      reg381 <= ((!forvar351[(2'h2):(1'h0)]) ?
                          $signed(($unsigned(forvar388) ?
                              (forvar374 < reg376) : wire346)) : ($unsigned((reg332 ?
                              reg270 : (8'hab))) << $unsigned({forvar376})));
                      reg382 <= (^$signed($unsigned({forvar353})));
                      reg383 <= forvar368[(1'h0):(1'h0)];
                    end
                end
            end
          if (((((+reg311) & $signed(reg280)) ^~ ((reg238 ?
                  (8'h9c) : reg303) <= (-reg358))) ?
              $signed(($signed(reg258) & (reg343 >> (8'hab)))) : reg360[(3'h5):(1'h0)]))
            begin
              if ((($unsigned((~^reg338)) ?
                  reg303 : ((reg258 <<< reg317) <= $signed(reg255))) ^ (reg271[(4'ha):(3'h5)] - $unsigned(reg281))))
                begin
                  for (forvar384 = (1'h0); (forvar384 < (1'h0)); forvar384 = (forvar384 + (1'h1)))
                    begin
                      reg385 <= $unsigned((((8'ha7) != forvar351) ?
                          ($unsigned(reg366) ?
                              forvar359[(3'h5):(2'h2)] : reg334) : (-$signed((8'ha4)))));
                      reg386 <= reg274;
                    end
                  reg387 <= (reg380 ?
                      ($unsigned((8'h9f)) ?
                          {(-wire233)} : reg283[(3'h4):(1'h1)]) : forvar351[(1'h0):(1'h0)]);
                  reg388 <= ({$unsigned((forvar385 ?
                          (8'h9f) : reg280))} && $signed(reg274[(1'h0):(1'h0)]));
                  reg389 <= $signed(reg303);
                end
              else
                begin
                  for (forvar384 = (1'h0); (forvar384 < (2'h3)); forvar384 = (forvar384 + (1'h1)))
                    begin
                      reg385 <= $unsigned(reg397);
                      reg386 <= $signed(($unsigned(reg272[(1'h1):(1'h1)]) ?
                          reg402 : {forvar352[(3'h6):(2'h2)]}));
                      reg387 <= $signed((~|{reg373}));
                    end
                end
            end
          else
            begin
              for (forvar384 = (1'h0); (forvar384 < (1'h0)); forvar384 = (forvar384 + (1'h1)))
                begin
                  if ($unsigned(reg313))
                    begin
                      reg385 <= reg399;
                      reg386 <= reg274[(1'h1):(1'h0)];
                      reg387 <= reg371;
                      reg388 <= reg303;
                    end
                  else
                    begin
                      reg385 <= ($signed(reg284) ?
                          (8'hac) : $signed((-(reg243 <= reg253))));
                      reg386 <= (8'hb4);
                      reg387 <= $unsigned(((wire233[(1'h1):(1'h1)] && $signed((8'ha7))) ?
                          reg345[(4'h9):(3'h7)] : (~|(reg260 != reg242))));
                      reg388 <= $unsigned(({((8'haf) ^ forvar370)} & (reg372 - (8'hb3))));
                    end
                end
            end
        end
      if ((&{{reg366[(2'h2):(1'h0)]}}))
        begin
          reg403 <= reg321;
          for (forvar404 = (1'h0); (forvar404 < (1'h1)); forvar404 = (forvar404 + (1'h1)))
            begin
              for (forvar405 = (1'h0); (forvar405 < (2'h3)); forvar405 = (forvar405 + (1'h1)))
                begin
                  if ({reg363[(3'h4):(1'h0)]})
                    begin
                      reg406 <= $unsigned(forvar370);
                    end
                  else
                    begin
                      reg406 <= wire348;
                    end
                  for (forvar407 = (1'h0); (forvar407 < (2'h3)); forvar407 = (forvar407 + (1'h1)))
                    begin
                      reg408 <= ($unsigned(($signed(reg388) ?
                              (~^reg332) : $unsigned(reg317))) ?
                          (($unsigned(reg302) ?
                              $signed(wire349) : (reg342 ?
                                  reg339 : reg271)) == reg293) : (&((&reg268) ?
                              $signed(reg352) : reg236[(4'ha):(3'h6)])));
                      reg409 <= ($unsigned($signed($signed((8'hb3)))) ?
                          $unsigned(($unsigned(reg370) ?
                              $signed(reg355) : $signed((8'ha0)))) : $signed((reg254 <<< $unsigned(reg290))));
                      reg410 <= (forvar359[(2'h2):(2'h2)] >= forvar350);
                      reg411 <= reg390;
                    end
                end
              if (reg303)
                begin
                  reg412 <= reg370;
                  if (reg399)
                    begin
                      reg413 <= $unsigned(reg275[(3'h6):(2'h2)]);
                      reg414 <= $unsigned((((|reg250) < (reg352 ?
                              reg403 : reg397)) ?
                          ($signed(reg342) ?
                              (^~reg277) : (reg394 ^ (8'hb0))) : $signed($signed(reg317))));
                    end
                  else
                    begin
                      reg413 <= forvar398[(1'h1):(1'h1)];
                      reg414 <= ($unsigned(reg320[(2'h3):(2'h2)]) ?
                          (8'hab) : (reg257[(3'h4):(2'h3)] != $signed($signed(reg358))));
                      reg415 <= ((((~&reg285) ?
                              (reg327 ? reg281 : reg376) : (^(8'ha7))) ?
                          $unsigned(reg317) : (^{reg343})) >= $signed(reg344[(4'hd):(3'h5)]));
                      reg416 <= reg282[(3'h5):(3'h4)];
                    end
                  if (reg332)
                    begin
                      reg417 <= {reg329};
                      reg418 <= (8'hb4);
                      reg419 <= reg257[(3'h7):(3'h5)];
                      reg420 <= ({$signed((^~reg272))} | $unsigned(reg340));
                    end
                  else
                    begin
                      reg417 <= (($signed((wire349 ?
                              reg242 : (8'hb0))) << $signed($unsigned(reg392))) ?
                          $signed((+$signed(forvar385))) : (reg326 ?
                              {(~forvar367)} : reg290[(1'h0):(1'h0)]));
                      reg418 <= forvar360;
                    end
                end
              else
                begin
                  if ($unsigned((reg352[(3'h6):(3'h5)] ?
                      $unsigned(((8'hac) | reg284)) : reg388[(1'h1):(1'h1)])))
                    begin
                      reg412 <= $unsigned(reg371[(4'h9):(3'h4)]);
                      reg413 <= (reg382 || reg245);
                      reg414 <= {$signed($signed($unsigned(reg371)))};
                    end
                  else
                    begin
                      reg412 <= reg364;
                      reg413 <= (^~reg267[(3'h6):(3'h6)]);
                    end
                end
            end
          for (forvar421 = (1'h0); (forvar421 < (2'h3)); forvar421 = (forvar421 + (1'h1)))
            begin
              reg422 <= reg401;
              reg423 <= $unsigned(($signed((!wire233)) != $signed((reg419 ?
                  reg338 : reg363))));
              reg424 <= (reg237 ? reg258 : $unsigned((~^forvar393)));
            end
          for (forvar425 = (1'h0); (forvar425 < (1'h1)); forvar425 = (forvar425 + (1'h1)))
            begin
              reg426 <= (~&(~&((wire346 ^~ forvar365) ?
                  (forvar367 ? forvar388 : (8'haf)) : (reg373 ?
                      reg381 : (8'haa)))));
              reg427 <= ($signed(reg371) && {($unsigned(reg309) ?
                      reg370 : reg388)});
              reg428 <= $signed(forvar421);
              for (forvar429 = (1'h0); (forvar429 < (2'h3)); forvar429 = (forvar429 + (1'h1)))
                begin
                  for (forvar430 = (1'h0); (forvar430 < (1'h0)); forvar430 = (forvar430 + (1'h1)))
                    begin
                      reg431 <= (^~$signed(reg375));
                      reg432 <= (reg314[(3'h4):(2'h2)] ?
                          {$signed((reg323 ^ reg388))} : {(reg258 ^~ (reg380 && forvar407))});
                      reg433 <= reg315[(2'h2):(1'h0)];
                    end
                  if ($signed(reg245[(3'h5):(2'h3)]))
                    begin
                      reg434 <= (8'had);
                      reg435 <= (8'hb8);
                      reg436 <= reg265[(4'he):(4'ha)];
                    end
                  else
                    begin
                      reg434 <= reg422[(2'h3):(2'h2)];
                      reg435 <= reg391;
                      reg436 <= (reg406[(4'he):(4'hd)] && wire347[(3'h4):(1'h0)]);
                    end
                  if (reg406)
                    begin
                      reg437 <= (^~$unsigned(reg402[(1'h0):(1'h0)]));
                      reg438 <= ({({reg307} ?
                                  reg343[(2'h3):(1'h0)] : $signed((8'ha1)))} ?
                          $signed(reg418) : reg383);
                      reg439 <= (8'hb6);
                    end
                  else
                    begin
                      reg437 <= (((^~reg302) ?
                          reg434[(3'h7):(2'h3)] : ((~&reg322) ?
                              (^~reg252) : reg386[(2'h2):(2'h2)])) || (($unsigned(reg373) ?
                          $unsigned(reg261) : (forvar352 ?
                              reg270 : reg386)) >= ($signed(reg400) ?
                          ((8'hb7) ?
                              reg244 : reg312) : reg265[(4'hb):(1'h1)])));
                      reg438 <= {(~^(^~((8'haf) ? reg371 : reg354)))};
                      reg439 <= $unsigned($signed(reg358[(1'h0):(1'h0)]));
                      reg440 <= ($signed(reg338) > $signed(((reg431 ?
                              reg265 : reg285) ?
                          $signed((8'hb4)) : (reg327 <= reg368))));
                    end
                end
            end
        end
      else
        begin
          reg403 <= $unsigned($signed(forvar421));
        end
      reg441 <= {forvar367[(1'h0):(1'h0)]};
      if (forvar398)
        begin
          if ($unsigned(reg377))
            begin
              for (forvar442 = (1'h0); (forvar442 < (2'h3)); forvar442 = (forvar442 + (1'h1)))
                begin
                  if ($signed($signed((reg291 <= reg417[(3'h5):(1'h0)]))))
                    begin
                      reg443 <= reg374[(4'ha):(3'h4)];
                      reg444 <= ((((reg320 && reg276) + forvar393) ~^ (!(8'hb3))) ?
                          (^reg247) : $signed($signed($unsigned(forvar374))));
                    end
                  else
                    begin
                      reg443 <= reg255[(1'h1):(1'h0)];
                      reg444 <= (~(^~$unsigned(forvar398[(1'h1):(1'h1)])));
                    end
                  for (forvar445 = (1'h0); (forvar445 < (1'h1)); forvar445 = (forvar445 + (1'h1)))
                    begin
                      reg446 <= $unsigned((reg414[(2'h2):(1'h1)] * $unsigned((reg358 ?
                          reg291 : reg327))));
                      reg447 <= reg446[(2'h2):(1'h0)];
                      reg448 <= ((({reg272} > reg281[(2'h2):(1'h0)]) ?
                              reg239 : ($unsigned(forvar388) >= reg293[(3'h7):(3'h6)])) ?
                          ($signed((^reg284)) > ($unsigned(forvar407) == reg440)) : $unsigned(reg432));
                    end
                end
              reg449 <= (forvar445 >> (8'hb1));
              if ({$unsigned($unsigned((8'hb4)))})
                begin
                  if ((~|$signed(((reg297 ? reg326 : reg257) ?
                      reg447 : {reg313}))))
                    begin
                      reg450 <= $signed((((reg384 | reg440) <<< reg441) ?
                          (^~(reg388 << forvar393)) : forvar351[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg450 <= $unsigned({reg373[(1'h1):(1'h1)]});
                      reg451 <= {((reg415[(1'h0):(1'h0)] + reg321[(4'ha):(3'h4)]) == ((reg409 == forvar393) && $signed((8'h9d))))};
                      reg452 <= (reg258 & ($unsigned((8'ha9)) != (+$signed(forvar374))));
                    end
                  if (((~^($unsigned(reg452) ?
                      $unsigned(reg389) : (reg420 | forvar367))) >>> reg321[(1'h0):(1'h0)]))
                    begin
                      reg453 <= reg397[(2'h3):(1'h1)];
                      reg454 <= reg453;
                      reg455 <= (&reg252);
                      reg456 <= reg356;
                    end
                  else
                    begin
                      reg453 <= (wire349 && ((~^reg343) ?
                          ($signed(reg427) <<< reg257) : $signed((reg309 ?
                              forvar404 : reg270))));
                      reg454 <= reg242;
                      reg455 <= ((&$signed(reg318[(1'h0):(1'h0)])) ?
                          ((reg297[(1'h1):(1'h0)] ?
                                  (reg309 > reg449) : (reg374 ?
                                      reg387 : reg415)) ?
                              reg328[(3'h5):(2'h3)] : ((forvar382 ?
                                      reg259 : reg253) ?
                                  (^~(8'hb2)) : reg334)) : reg276);
                      reg456 <= (-reg263[(2'h3):(2'h2)]);
                    end
                  for (forvar457 = (1'h0); (forvar457 < (1'h0)); forvar457 = (forvar457 + (1'h1)))
                    begin
                      reg458 <= {reg250};
                    end
                end
              else
                begin
                  for (forvar450 = (1'h0); (forvar450 < (2'h2)); forvar450 = (forvar450 + (1'h1)))
                    begin
                      reg451 <= ((~^((wire233 >= reg334) >= (reg310 != forvar388))) & (-((reg322 ?
                              reg367 : forvar382) ?
                          (reg300 & reg261) : forvar384)));
                      reg452 <= $signed((reg275 && $unsigned(wire348)));
                    end
                  reg453 <= reg418;
                end
              if ($signed($unsigned($signed(reg426[(3'h5):(3'h4)]))))
                begin
                  if (reg317[(3'h5):(1'h0)])
                    begin
                      reg459 <= forvar429;
                      reg460 <= reg326;
                      reg461 <= (forvar398 ?
                          $signed(reg417[(1'h1):(1'h1)]) : $signed(reg298));
                      reg462 <= reg370[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg459 <= {reg459[(4'hb):(4'ha)]};
                      reg460 <= $signed($signed(((reg355 ~^ forvar398) <<< reg350[(3'h4):(2'h3)])));
                      reg461 <= $unsigned(reg391[(3'h5):(3'h5)]);
                    end
                  if ({$unsigned((reg454[(2'h2):(2'h2)] ?
                          {(8'h9d)} : $signed(reg283)))})
                    begin
                      reg463 <= reg253[(3'h7):(2'h2)];
                    end
                  else
                    begin
                      reg463 <= reg313[(1'h0):(1'h0)];
                      reg464 <= ($unsigned($unsigned(forvar351[(1'h0):(1'h0)])) << reg289[(3'h7):(3'h4)]);
                    end
                  if ((&(((reg350 ? forvar359 : reg350) ?
                      (^~reg383) : (reg329 ? forvar384 : (8'ha8))) >> wire349)))
                    begin
                      reg465 <= (($unsigned($unsigned((8'ha7))) * reg272[(1'h0):(1'h0)]) ?
                          reg256 : reg360[(3'h5):(1'h1)]);
                      reg466 <= $signed((~^reg437[(3'h5):(3'h4)]));
                      reg467 <= forvar352[(3'h5):(1'h1)];
                      reg468 <= ((((reg383 ? reg459 : reg396) >>> (~^reg455)) ?
                              forvar351[(2'h2):(1'h0)] : reg463[(3'h4):(1'h1)]) ?
                          (-reg373) : ($signed((reg432 > (8'hb3))) ?
                              ((|reg293) || (reg314 ?
                                  reg380 : forvar382)) : ((+reg383) ?
                                  reg256 : (&reg298))));
                    end
                  else
                    begin
                      reg465 <= reg322[(4'h8):(3'h5)];
                      reg466 <= $signed(({(~^reg310)} ^ reg390[(2'h3):(1'h1)]));
                      reg467 <= reg381[(4'h9):(4'h8)];
                    end
                  reg469 <= (-($unsigned((+reg310)) - $signed(reg359)));
                end
              else
                begin
                  reg459 <= (($unsigned(reg350[(3'h5):(2'h3)]) ?
                      $signed(((8'h9f) ?
                          (8'hb9) : reg412)) : reg370[(1'h0):(1'h0)]) >>> {(&reg339[(4'h8):(3'h4)])});
                end
            end
          else
            begin
              if (reg343)
                begin
                  if (reg334[(4'ha):(4'h8)])
                    begin
                      reg442 <= reg363;
                      reg443 <= $signed(reg360[(1'h1):(1'h0)]);
                      reg444 <= (+(^~$unsigned({reg414})));
                      reg445 <= reg402;
                    end
                  else
                    begin
                      reg442 <= {(($signed(reg363) ?
                              ((8'h9e) - reg258) : $signed(forvar373)) != ($signed(reg270) << reg289))};
                    end
                  reg446 <= {(8'hac)};
                  for (forvar447 = (1'h0); (forvar447 < (2'h3)); forvar447 = (forvar447 + (1'h1)))
                    begin
                      reg448 <= (^(&(&(forvar388 && forvar359))));
                      reg449 <= $signed($signed((^(reg317 <= (8'ha7)))));
                    end
                  for (forvar450 = (1'h0); (forvar450 < (1'h1)); forvar450 = (forvar450 + (1'h1)))
                    begin
                      reg451 <= $signed(reg440[(2'h2):(1'h1)]);
                      reg452 <= (!$unsigned(reg394));
                      reg453 <= ((|(~^$signed(reg411))) ?
                          ($unsigned(reg419[(3'h7):(3'h7)]) ?
                              ((reg253 ?
                                  reg261 : (8'hb3)) >> (reg434 <= reg386)) : (~|forvar368)) : reg417);
                      reg454 <= {$unsigned({reg301[(2'h2):(1'h1)]})};
                    end
                end
              else
                begin
                  reg442 <= ($unsigned($signed((^forvar447))) >> (!((reg370 ?
                      (8'hb3) : reg301) != reg322)));
                  for (forvar443 = (1'h0); (forvar443 < (2'h2)); forvar443 = (forvar443 + (1'h1)))
                    begin
                      reg444 <= reg375[(1'h0):(1'h0)];
                    end
                  for (forvar445 = (1'h0); (forvar445 < (1'h1)); forvar445 = (forvar445 + (1'h1)))
                    begin
                      reg446 <= ($signed((~|$unsigned(reg406))) ?
                          forvar404 : {reg419[(3'h6):(2'h2)]});
                      reg447 <= $signed((~^$signed((reg374 != reg356))));
                    end
                  reg448 <= reg468;
                end
              if ($unsigned(((~((8'hac) ?
                  reg443 : reg320)) + ($signed((8'ha6)) & (reg249 ?
                  reg307 : reg444)))))
                begin
                  for (forvar455 = (1'h0); (forvar455 < (1'h0)); forvar455 = (forvar455 + (1'h1)))
                    begin
                      reg456 <= (forvar358[(2'h3):(1'h0)] & reg260);
                    end
                  if ($unsigned($signed(((reg418 < (8'had)) ?
                      (reg369 ? (8'hae) : reg317) : forvar450[(1'h1):(1'h1)]))))
                    begin
                      reg457 <= $unsigned((((reg325 ? reg345 : reg444) ?
                          (+(8'haf)) : $signed((8'haa))) >= reg388[(1'h0):(1'h0)]));
                      reg458 <= (^($signed(((8'h9f) ^ forvar360)) ?
                          {{forvar382}} : ((reg457 ? reg327 : reg314) ?
                              reg258[(2'h2):(1'h0)] : $signed(forvar457))));
                    end
                  else
                    begin
                      reg457 <= reg376[(1'h1):(1'h0)];
                      reg458 <= $unsigned(reg256);
                    end
                end
              else
                begin
                  for (forvar455 = (1'h0); (forvar455 < (2'h3)); forvar455 = (forvar455 + (1'h1)))
                    begin
                      reg456 <= reg278;
                      reg457 <= ($signed(reg387[(2'h2):(2'h2)]) ?
                          forvar425[(4'h8):(1'h1)] : reg287[(2'h2):(1'h0)]);
                      reg458 <= reg431;
                    end
                end
              if ($signed(forvar447[(3'h6):(1'h1)]))
                begin
                  if (($signed(($signed((8'h9f)) << {(8'ha0)})) & reg408[(3'h4):(1'h0)]))
                    begin
                      reg459 <= wire233;
                      reg460 <= {(reg243 < $signed((8'ha7)))};
                      reg461 <= (reg257 <= reg385);
                      reg462 <= (~|$signed((-(!reg361))));
                    end
                  else
                    begin
                      reg459 <= ((~(forvar376[(2'h3):(1'h0)] ?
                          (reg261 ^ reg359) : (reg297 > reg318))) ~^ (forvar455 ?
                          reg451 : ((reg394 - reg328) ^ forvar382)));
                      reg460 <= (~&($unsigned($signed(forvar367)) ?
                          $signed($signed(reg283)) : reg322));
                    end
                end
              else
                begin
                  for (forvar459 = (1'h0); (forvar459 < (1'h0)); forvar459 = (forvar459 + (1'h1)))
                    begin
                      reg460 <= {$signed(forvar450)};
                      reg461 <= $signed($signed((&(^~(8'h9c)))));
                    end
                  reg462 <= $unsigned((~|{(-forvar388)}));
                  for (forvar463 = (1'h0); (forvar463 < (1'h0)); forvar463 = (forvar463 + (1'h1)))
                    begin
                      reg464 <= (8'hb5);
                    end
                end
              for (forvar465 = (1'h0); (forvar465 < (1'h0)); forvar465 = (forvar465 + (1'h1)))
                begin
                  for (forvar466 = (1'h0); (forvar466 < (2'h2)); forvar466 = (forvar466 + (1'h1)))
                    begin
                      reg467 <= {$unsigned((+forvar447[(1'h0):(1'h0)]))};
                      reg468 <= ($signed((reg340 && (-(8'hab)))) >= reg364[(3'h4):(3'h4)]);
                      reg469 <= $unsigned((^~$signed({reg368})));
                    end
                end
            end
          if ((reg247 ? (&reg283[(4'hb):(4'h8)]) : reg411[(3'h6):(1'h0)]))
            begin
              for (forvar470 = (1'h0); (forvar470 < (2'h3)); forvar470 = (forvar470 + (1'h1)))
                begin
                  for (forvar471 = (1'h0); (forvar471 < (1'h0)); forvar471 = (forvar471 + (1'h1)))
                    begin
                      reg472 <= (~|$signed(reg318[(1'h1):(1'h0)]));
                      reg473 <= (-reg249[(4'hb):(4'h8)]);
                    end
                  for (forvar474 = (1'h0); (forvar474 < (2'h2)); forvar474 = (forvar474 + (1'h1)))
                    begin
                      reg475 <= reg370;
                      reg476 <= (|$unsigned(reg382[(3'h7):(1'h0)]));
                      reg477 <= reg435[(3'h6):(3'h4)];
                    end
                end
            end
          else
            begin
              reg470 <= $unsigned($unsigned((8'ha3)));
            end
          if ($unsigned($signed(((8'ha6) && {reg360}))))
            begin
              if (((~$signed($unsigned(wire232))) >>> reg423))
                begin
                  for (forvar478 = (1'h0); (forvar478 < (2'h3)); forvar478 = (forvar478 + (1'h1)))
                    begin
                      reg479 <= reg374[(2'h3):(1'h1)];
                      reg480 <= (((^~(forvar404 ?
                          forvar443 : reg323)) ^~ reg438[(1'h1):(1'h0)]) && reg475);
                      reg481 <= $unsigned(reg336[(4'hc):(1'h1)]);
                      reg482 <= (reg306 ^ $unsigned(reg355));
                    end
                  for (forvar483 = (1'h0); (forvar483 < (1'h1)); forvar483 = (forvar483 + (1'h1)))
                    begin
                      reg484 <= $signed(reg355[(4'hc):(4'h8)]);
                      reg485 <= (8'hb5);
                      reg486 <= (((reg366[(3'h5):(3'h5)] << $signed(forvar374)) || $unsigned($signed(reg481))) ?
                          $unsigned($unsigned(reg409[(1'h1):(1'h1)])) : (-(reg361[(1'h0):(1'h0)] <= ((8'h9c) ?
                              reg414 : reg482))));
                      reg487 <= ((~(~|reg399)) && $signed(reg342[(3'h5):(3'h5)]));
                    end
                end
              else
                begin
                  if (((forvar353[(2'h2):(2'h2)] ?
                          $signed((+forvar430)) : ((-forvar359) ~^ reg402)) ?
                      (~$signed(reg298[(4'ha):(1'h1)])) : ((reg385[(2'h2):(1'h1)] ?
                          (~&(8'haf)) : (+forvar425)) && ((reg462 & reg247) ?
                          (+reg273) : reg357[(2'h2):(1'h0)]))))
                    begin
                      reg478 <= wire234[(3'h4):(2'h3)];
                      reg479 <= {(~^($signed(reg259) ?
                              (forvar351 ? forvar360 : reg410) : ((8'hb4) ?
                                  reg243 : (8'ha1))))};
                      reg480 <= reg260[(3'h6):(3'h5)];
                      reg481 <= $signed($unsigned((^~reg365)));
                    end
                  else
                    begin
                      reg478 <= $signed(reg432);
                      reg479 <= ($unsigned(($unsigned(reg482) >> ((8'h9d) ?
                              reg436 : reg306))) ?
                          reg442[(3'h5):(2'h2)] : reg383[(4'ha):(2'h2)]);
                    end
                  for (forvar482 = (1'h0); (forvar482 < (1'h1)); forvar482 = (forvar482 + (1'h1)))
                    begin
                      reg483 <= $signed((((reg311 > reg440) >>> $signed(reg323)) & reg285[(1'h0):(1'h0)]));
                    end
                  for (forvar484 = (1'h0); (forvar484 < (1'h1)); forvar484 = (forvar484 + (1'h1)))
                    begin
                      reg485 <= (forvar360 ?
                          ((~^(reg447 & reg431)) ?
                              $unsigned((+wire346)) : reg461[(3'h5):(3'h5)]) : ($unsigned($unsigned(reg448)) << (reg338 ?
                              $signed(reg370) : (reg289 & reg343))));
                      reg486 <= $signed($signed((reg356[(2'h2):(1'h1)] ?
                          $signed(reg291) : reg406)));
                    end
                end
            end
          else
            begin
              if ({$signed({(forvar381 ^ (8'ha5))})})
                begin
                  for (forvar478 = (1'h0); (forvar478 < (2'h3)); forvar478 = (forvar478 + (1'h1)))
                    begin
                      reg479 <= $signed(reg475);
                      reg480 <= (((~&(^~reg477)) - (reg415 != (reg273 ?
                          reg369 : reg241))) || (~reg417[(3'h4):(2'h2)]));
                    end
                  if (((((reg248 ? reg264 : forvar429) ?
                          $signed(reg449) : $signed(reg261)) < $signed($signed((8'ha8)))) ?
                      forvar455[(2'h3):(2'h3)] : $signed((forvar457 ?
                          reg280[(3'h4):(2'h2)] : $unsigned(reg306)))))
                    begin
                      reg481 <= reg411;
                      reg482 <= {reg339[(3'h6):(3'h4)]};
                      reg483 <= reg484[(4'hc):(3'h7)];
                    end
                  else
                    begin
                      reg481 <= $signed((($signed(reg391) << {reg240}) - (^~(reg326 >> reg306))));
                      reg482 <= ($unsigned(reg478[(1'h1):(1'h1)]) >= $signed(((reg314 ?
                              reg239 : reg381) ?
                          reg261[(3'h4):(1'h1)] : wire228[(1'h1):(1'h0)])));
                    end
                  for (forvar484 = (1'h0); (forvar484 < (2'h3)); forvar484 = (forvar484 + (1'h1)))
                    begin
                      reg485 <= {$unsigned(reg389)};
                      reg486 <= reg448;
                      reg487 <= (reg463 + ({{reg329}} ~^ {(8'hb8)}));
                    end
                end
              else
                begin
                  for (forvar478 = (1'h0); (forvar478 < (1'h0)); forvar478 = (forvar478 + (1'h1)))
                    begin
                      reg479 <= $unsigned(forvar470[(4'h8):(3'h4)]);
                      reg480 <= (reg371 ?
                          reg319 : ((~^$unsigned(reg242)) ?
                              (~$signed((8'haa))) : (!$unsigned(forvar445))));
                    end
                  for (forvar481 = (1'h0); (forvar481 < (1'h1)); forvar481 = (forvar481 + (1'h1)))
                    begin
                      reg482 <= {(((reg330 >> reg273) <<< $unsigned((8'hb2))) * reg373[(1'h0):(1'h0)])};
                      reg483 <= reg371;
                      reg484 <= (reg388 ?
                          (reg469[(2'h2):(1'h0)] ?
                              reg241 : (~|(reg313 ?
                                  reg333 : reg417))) : {(^(~reg365))});
                    end
                end
            end
        end
      else
        begin
          for (forvar442 = (1'h0); (forvar442 < (2'h3)); forvar442 = (forvar442 + (1'h1)))
            begin
              for (forvar443 = (1'h0); (forvar443 < (1'h0)); forvar443 = (forvar443 + (1'h1)))
                begin
                  for (forvar444 = (1'h0); (forvar444 < (1'h1)); forvar444 = (forvar444 + (1'h1)))
                    begin
                      reg445 <= $signed({(~|reg359)});
                      reg446 <= $signed((reg479 >>> reg367));
                      reg447 <= $signed(($unsigned({reg298}) ?
                          reg369 : (~reg269)));
                    end
                  for (forvar448 = (1'h0); (forvar448 < (1'h0)); forvar448 = (forvar448 + (1'h1)))
                    begin
                      reg449 <= $signed($signed(reg426));
                      reg450 <= {reg271[(1'h0):(1'h0)]};
                      reg451 <= $signed({$unsigned($signed(forvar442))});
                    end
                end
              for (forvar452 = (1'h0); (forvar452 < (2'h3)); forvar452 = (forvar452 + (1'h1)))
                begin
                  if ((reg260[(4'ha):(3'h6)] < forvar463[(2'h2):(1'h1)]))
                    begin
                      reg453 <= {wire234};
                      reg454 <= (reg424 >>> $signed($unsigned((~reg363))));
                    end
                  else
                    begin
                      reg453 <= reg466;
                      reg454 <= $signed(reg291);
                      reg455 <= reg273[(3'h7):(1'h1)];
                      reg456 <= $signed(reg353);
                    end
                end
              if ((reg388[(2'h2):(2'h2)] >= (reg262 ?
                  (~&forvar444) : reg453[(2'h3):(2'h3)])))
                begin
                  for (forvar457 = (1'h0); (forvar457 < (1'h0)); forvar457 = (forvar457 + (1'h1)))
                    begin
                      reg458 <= reg390[(3'h4):(1'h0)];
                      reg459 <= reg285;
                      reg460 <= (-$unsigned($signed((reg382 ?
                          reg390 : reg469))));
                      reg461 <= forvar370[(4'h8):(1'h0)];
                    end
                  if (($unsigned(reg306[(4'h9):(3'h7)]) ?
                      (({forvar398} ? (8'had) : (8'hb5)) != $unsigned((reg353 ?
                          reg353 : (8'hb3)))) : ($signed($signed(reg306)) ?
                          reg439[(4'ha):(3'h5)] : (((8'ha6) ? reg312 : reg452) ?
                              {reg260} : (forvar373 <<< wire346)))))
                    begin
                      reg462 <= reg343[(3'h7):(3'h5)];
                      reg463 <= $signed((8'hb7));
                    end
                  else
                    begin
                      reg462 <= $unsigned($unsigned((reg315 <= $unsigned(reg479))));
                      reg463 <= reg250;
                      reg464 <= ($unsigned(reg362) << (8'ha1));
                      reg465 <= (8'hb7);
                    end
                  if (((8'hb6) || reg479))
                    begin
                      reg466 <= $unsigned($unsigned($unsigned((reg468 ?
                          (8'hb1) : reg358))));
                      reg467 <= reg460[(1'h0):(1'h0)];
                      reg468 <= forvar447;
                    end
                  else
                    begin
                      reg466 <= ({{$signed((8'h9c))}} >> {reg323[(3'h5):(3'h5)]});
                      reg467 <= (!reg400);
                      reg468 <= $signed((reg451[(3'h7):(2'h3)] << (reg329 >= (8'ha6))));
                      reg469 <= (reg416[(2'h2):(1'h0)] ?
                          $unsigned($signed($signed((8'ha8)))) : reg300);
                    end
                  for (forvar470 = (1'h0); (forvar470 < (1'h1)); forvar470 = (forvar470 + (1'h1)))
                    begin
                      reg471 <= $unsigned(reg449);
                      reg472 <= ($signed({reg424}) * (~&(reg374 ~^ reg463[(1'h0):(1'h0)])));
                      reg473 <= $unsigned((reg363[(1'h1):(1'h1)] ^ (~$unsigned(reg415))));
                    end
                end
              else
                begin
                  reg457 <= ((~^(reg240 << reg280)) >>> reg236);
                end
            end
        end
    end
  assign wire488 = $signed(($signed((8'hba)) << $signed((wire346 ?
                       (8'hb5) : reg428))));
  assign wire489 = (($unsigned(reg438) ?
                           $unsigned((reg277 ? reg456 : reg466)) : ({reg460} ?
                               (8'hb1) : $unsigned(reg263))) ?
                       {reg358} : reg243[(3'h4):(2'h2)]);
  assign wire490 = reg320;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1186  (y, clk, wire1187, wire1188, wire1189, wire1190, wire1191);
  output wire [(32'h186e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire1187;
  input wire [(4'ha):(1'h0)] wire1188;
  input wire [(3'h7):(1'h0)] wire1189;
  input wire signed [(4'hd):(1'h0)] wire1190;
  input wire signed [(4'ha):(1'h0)] wire1191;
  wire signed [(4'ha):(1'h0)] wire3223;
  wire signed [(4'hb):(1'h0)] wire3021;
  wire [(4'ha):(1'h0)] wire2837;
  wire [(4'h8):(1'h0)] wire1192;
  wire signed [(3'h5):(1'h0)] wire1193;
  wire [(3'h5):(1'h0)] wire1241;
  wire [(4'h9):(1'h0)] wire2706;
  reg signed [(3'h4):(1'h0)] reg3222 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3221 = (1'h0);
  reg [(4'h9):(1'h0)] reg3209 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3218 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3217 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3216 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3215 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3214 = (1'h0);
  reg [(3'h6):(1'h0)] reg3213 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3212 = (1'h0);
  reg [(4'he):(1'h0)] reg3211 = (1'h0);
  reg [(4'hd):(1'h0)] reg3210 = (1'h0);
  reg [(3'h6):(1'h0)] reg3208 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3207 = (1'h0);
  reg [(5'h10):(1'h0)] reg3206 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3202 = (1'h0);
  reg [(4'h9):(1'h0)] reg3205 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3204 = (1'h0);
  reg [(4'h9):(1'h0)] reg3203 = (1'h0);
  reg [(3'h5):(1'h0)] reg3201 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3200 = (1'h0);
  reg [(5'h10):(1'h0)] reg3199 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3198 = (1'h0);
  reg [(4'hc):(1'h0)] reg3197 = (1'h0);
  reg [(4'hc):(1'h0)] reg3195 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3194 = (1'h0);
  reg [(4'hd):(1'h0)] reg3193 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3192 = (1'h0);
  reg [(2'h3):(1'h0)] reg3191 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3190 = (1'h0);
  reg [(4'h9):(1'h0)] reg3189 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3188 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3187 = (1'h0);
  reg [(4'hf):(1'h0)] reg3186 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3185 = (1'h0);
  reg [(4'h8):(1'h0)] reg3184 = (1'h0);
  reg [(4'hc):(1'h0)] reg3183 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3182 = (1'h0);
  reg [(4'hd):(1'h0)] reg3181 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3180 = (1'h0);
  reg [(2'h2):(1'h0)] reg3177 = (1'h0);
  reg [(3'h5):(1'h0)] reg3176 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3175 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3174 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3172 = (1'h0);
  reg [(4'hd):(1'h0)] reg3171 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3170 = (1'h0);
  reg [(3'h7):(1'h0)] reg3168 = (1'h0);
  reg [(4'hf):(1'h0)] reg3167 = (1'h0);
  reg [(3'h5):(1'h0)] reg3166 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3165 = (1'h0);
  reg [(4'h9):(1'h0)] reg3164 = (1'h0);
  reg [(4'hc):(1'h0)] reg3163 = (1'h0);
  reg [(3'h7):(1'h0)] reg3162 = (1'h0);
  reg [(4'h9):(1'h0)] reg3161 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3159 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3157 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3156 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3155 = (1'h0);
  reg [(4'ha):(1'h0)] reg3154 = (1'h0);
  reg [(2'h3):(1'h0)] reg3153 = (1'h0);
  reg [(2'h2):(1'h0)] reg3151 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3150 = (1'h0);
  reg [(2'h2):(1'h0)] reg3149 = (1'h0);
  reg [(4'hc):(1'h0)] reg3144 = (1'h0);
  reg [(4'h9):(1'h0)] reg3143 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3142 = (1'h0);
  reg [(4'ha):(1'h0)] reg3141 = (1'h0);
  reg [(4'hb):(1'h0)] reg3139 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3138 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3137 = (1'h0);
  reg [(4'hf):(1'h0)] reg3133 = (1'h0);
  reg [(3'h7):(1'h0)] reg3062 = (1'h0);
  reg [(4'h9):(1'h0)] reg3058 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3132 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3131 = (1'h0);
  reg [(3'h6):(1'h0)] reg3130 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3129 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3128 = (1'h0);
  reg [(4'hf):(1'h0)] reg3127 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3126 = (1'h0);
  reg [(2'h3):(1'h0)] reg3125 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3124 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3123 = (1'h0);
  reg [(4'h8):(1'h0)] reg3121 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3120 = (1'h0);
  reg [(4'h8):(1'h0)] reg3119 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3116 = (1'h0);
  reg [(4'hb):(1'h0)] reg3115 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3114 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3113 = (1'h0);
  reg [(3'h5):(1'h0)] reg3112 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3111 = (1'h0);
  reg [(4'hf):(1'h0)] reg3110 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3109 = (1'h0);
  reg [(3'h6):(1'h0)] reg3108 = (1'h0);
  reg [(5'h10):(1'h0)] reg3107 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3106 = (1'h0);
  reg [(2'h3):(1'h0)] reg3104 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3103 = (1'h0);
  reg [(4'ha):(1'h0)] reg3099 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3098 = (1'h0);
  reg [(4'h9):(1'h0)] reg3096 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3095 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3094 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3093 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3092 = (1'h0);
  reg [(4'hf):(1'h0)] reg3091 = (1'h0);
  reg [(5'h10):(1'h0)] reg3089 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3088 = (1'h0);
  reg [(4'hf):(1'h0)] reg3087 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3086 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3085 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3083 = (1'h0);
  reg [(4'hc):(1'h0)] reg3082 = (1'h0);
  reg [(2'h3):(1'h0)] reg3084 = (1'h0);
  reg [(3'h6):(1'h0)] reg3081 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3080 = (1'h0);
  reg [(3'h5):(1'h0)] reg3079 = (1'h0);
  reg [(2'h2):(1'h0)] reg3078 = (1'h0);
  reg [(4'h8):(1'h0)] reg3076 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3075 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3074 = (1'h0);
  reg [(3'h7):(1'h0)] reg3051 = (1'h0);
  reg [(4'he):(1'h0)] reg3071 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3069 = (1'h0);
  reg [(4'hd):(1'h0)] reg3073 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3072 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3070 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3068 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3067 = (1'h0);
  reg [(3'h4):(1'h0)] reg3066 = (1'h0);
  reg [(4'hd):(1'h0)] reg3065 = (1'h0);
  reg [(4'h9):(1'h0)] reg3064 = (1'h0);
  reg [(4'h8):(1'h0)] reg3063 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3061 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3060 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3059 = (1'h0);
  reg [(3'h7):(1'h0)] reg3057 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3056 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3055 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3054 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3053 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3052 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3050 = (1'h0);
  reg [(3'h5):(1'h0)] reg3049 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3048 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3043 = (1'h0);
  reg [(4'hf):(1'h0)] reg3042 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3036 = (1'h0);
  reg [(4'hd):(1'h0)] reg3023 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3038 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3035 = (1'h0);
  reg [(4'ha):(1'h0)] reg3033 = (1'h0);
  reg [(4'hd):(1'h0)] reg3047 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3046 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3045 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3044 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3041 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3040 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3039 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3037 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3034 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3032 = (1'h0);
  reg [(3'h6):(1'h0)] reg3024 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3031 = (1'h0);
  reg [(2'h3):(1'h0)] reg3030 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3029 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3028 = (1'h0);
  reg [(2'h2):(1'h0)] reg3027 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3026 = (1'h0);
  reg [(4'hd):(1'h0)] reg3025 = (1'h0);
  reg [(3'h5):(1'h0)] reg3022 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2996 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2995 = (1'h0);
  reg [(4'h9):(1'h0)] reg2984 = (1'h0);
  reg [(4'he):(1'h0)] reg2962 = (1'h0);
  reg [(4'he):(1'h0)] reg2977 = (1'h0);
  reg [(3'h6):(1'h0)] reg2965 = (1'h0);
  reg [(4'h8):(1'h0)] reg2964 = (1'h0);
  reg [(4'he):(1'h0)] reg3020 = (1'h0);
  reg [(3'h6):(1'h0)] reg2991 = (1'h0);
  reg [(4'hf):(1'h0)] reg3019 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3018 = (1'h0);
  reg [(4'hb):(1'h0)] reg3017 = (1'h0);
  reg [(4'hf):(1'h0)] reg3013 = (1'h0);
  reg [(4'hc):(1'h0)] reg3007 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3016 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3015 = (1'h0);
  reg [(4'hc):(1'h0)] reg3014 = (1'h0);
  reg [(3'h6):(1'h0)] reg3012 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3011 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3010 = (1'h0);
  reg [(2'h2):(1'h0)] reg3009 = (1'h0);
  reg [(4'hb):(1'h0)] reg3008 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3006 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3005 = (1'h0);
  reg [(2'h2):(1'h0)] reg3004 = (1'h0);
  reg [(4'h9):(1'h0)] reg3003 = (1'h0);
  reg [(4'he):(1'h0)] reg3002 = (1'h0);
  reg [(4'hf):(1'h0)] reg3001 = (1'h0);
  reg [(4'ha):(1'h0)] reg3000 = (1'h0);
  reg [(3'h5):(1'h0)] reg2999 = (1'h0);
  reg [(4'hc):(1'h0)] reg2998 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2997 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2994 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2993 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2992 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2987 = (1'h0);
  reg [(4'hf):(1'h0)] reg2990 = (1'h0);
  reg [(4'ha):(1'h0)] reg2989 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2988 = (1'h0);
  reg [(4'ha):(1'h0)] reg2986 = (1'h0);
  reg [(4'hd):(1'h0)] reg2985 = (1'h0);
  reg [(4'he):(1'h0)] reg2983 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2982 = (1'h0);
  reg [(4'ha):(1'h0)] reg2981 = (1'h0);
  reg [(4'hc):(1'h0)] reg2980 = (1'h0);
  reg [(4'h9):(1'h0)] reg2979 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2976 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2975 = (1'h0);
  reg [(3'h4):(1'h0)] reg2974 = (1'h0);
  reg [(2'h3):(1'h0)] reg2973 = (1'h0);
  reg [(4'hd):(1'h0)] reg2972 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2971 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2970 = (1'h0);
  reg [(4'hf):(1'h0)] reg2969 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2968 = (1'h0);
  reg [(4'hd):(1'h0)] reg2967 = (1'h0);
  reg [(3'h5):(1'h0)] reg2966 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2963 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2917 = (1'h0);
  reg [(2'h3):(1'h0)] reg2961 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2960 = (1'h0);
  reg [(4'ha):(1'h0)] reg2930 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2958 = (1'h0);
  reg [(4'h8):(1'h0)] reg2957 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2956 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2955 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2954 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2953 = (1'h0);
  reg [(5'h10):(1'h0)] reg2951 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2950 = (1'h0);
  reg [(3'h7):(1'h0)] reg2949 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2947 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2946 = (1'h0);
  reg [(3'h5):(1'h0)] reg2945 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2943 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2942 = (1'h0);
  reg [(4'ha):(1'h0)] reg2940 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2939 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2938 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2937 = (1'h0);
  reg [(4'he):(1'h0)] reg2936 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2935 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2934 = (1'h0);
  reg [(3'h5):(1'h0)] reg2931 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2918 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2929 = (1'h0);
  reg [(4'hc):(1'h0)] reg2928 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2927 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2926 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2925 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2924 = (1'h0);
  reg [(4'hb):(1'h0)] reg2923 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2922 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2921 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2920 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2919 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2916 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2915 = (1'h0);
  reg [(4'he):(1'h0)] reg2906 = (1'h0);
  reg [(4'hf):(1'h0)] reg2904 = (1'h0);
  reg [(4'hb):(1'h0)] reg2903 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2914 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2913 = (1'h0);
  reg [(4'h8):(1'h0)] reg2912 = (1'h0);
  reg [(4'hb):(1'h0)] reg2911 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2910 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2909 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2908 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2907 = (1'h0);
  reg [(4'hb):(1'h0)] reg2905 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2902 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2901 = (1'h0);
  reg [(4'h9):(1'h0)] reg2900 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2899 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2897 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2896 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2895 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2894 = (1'h0);
  reg [(4'h9):(1'h0)] reg2893 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2892 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2891 = (1'h0);
  reg [(4'hb):(1'h0)] reg2889 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2888 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2886 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2885 = (1'h0);
  reg [(4'h9):(1'h0)] reg2884 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2883 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2882 = (1'h0);
  reg [(4'h8):(1'h0)] reg2880 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2879 = (1'h0);
  reg [(4'hd):(1'h0)] reg2878 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2877 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2873 = (1'h0);
  reg [(3'h7):(1'h0)] reg2864 = (1'h0);
  reg [(4'hb):(1'h0)] reg2861 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2860 = (1'h0);
  reg [(4'hf):(1'h0)] reg2859 = (1'h0);
  reg [(4'hd):(1'h0)] reg2855 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2852 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2851 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2846 = (1'h0);
  reg [(3'h7):(1'h0)] reg2845 = (1'h0);
  reg [(3'h4):(1'h0)] reg2840 = (1'h0);
  reg [(5'h10):(1'h0)] reg2839 = (1'h0);
  reg [(2'h3):(1'h0)] reg2871 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2870 = (1'h0);
  reg [(2'h3):(1'h0)] reg2869 = (1'h0);
  reg [(2'h3):(1'h0)] reg2868 = (1'h0);
  reg [(3'h5):(1'h0)] reg2867 = (1'h0);
  reg [(4'ha):(1'h0)] reg2866 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2865 = (1'h0);
  reg [(3'h6):(1'h0)] reg2863 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2862 = (1'h0);
  reg [(2'h2):(1'h0)] reg2858 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2857 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2856 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2854 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2853 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2850 = (1'h0);
  reg [(2'h2):(1'h0)] reg2849 = (1'h0);
  reg [(4'hd):(1'h0)] reg2848 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2847 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2844 = (1'h0);
  reg [(4'h9):(1'h0)] reg2843 = (1'h0);
  reg [(4'h8):(1'h0)] reg2842 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2841 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2838 = (1'h0);
  reg [(3'h6):(1'h0)] reg2836 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2835 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2834 = (1'h0);
  reg [(4'he):(1'h0)] reg2833 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2831 = (1'h0);
  reg [(3'h7):(1'h0)] reg2830 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2829 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2825 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2821 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2819 = (1'h0);
  reg [(4'he):(1'h0)] reg2828 = (1'h0);
  reg [(2'h2):(1'h0)] reg2827 = (1'h0);
  reg [(2'h3):(1'h0)] reg2826 = (1'h0);
  reg [(4'hc):(1'h0)] reg2824 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2823 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2822 = (1'h0);
  reg [(4'hf):(1'h0)] reg2820 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2812 = (1'h0);
  reg [(4'hc):(1'h0)] reg2818 = (1'h0);
  reg [(3'h4):(1'h0)] reg2817 = (1'h0);
  reg [(3'h6):(1'h0)] reg2815 = (1'h0);
  reg [(5'h10):(1'h0)] reg2814 = (1'h0);
  reg [(3'h7):(1'h0)] reg2813 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2811 = (1'h0);
  reg [(4'hc):(1'h0)] reg2810 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2808 = (1'h0);
  reg [(2'h2):(1'h0)] reg2807 = (1'h0);
  reg [(4'hf):(1'h0)] reg2806 = (1'h0);
  reg [(4'hb):(1'h0)] reg2805 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2803 = (1'h0);
  reg [(2'h3):(1'h0)] reg2802 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2801 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2800 = (1'h0);
  reg [(4'h9):(1'h0)] reg2799 = (1'h0);
  reg [(4'ha):(1'h0)] reg2798 = (1'h0);
  reg [(4'h9):(1'h0)] reg2797 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2796 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2795 = (1'h0);
  reg [(4'hb):(1'h0)] reg2784 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2793 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2791 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2790 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2788 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2787 = (1'h0);
  reg [(2'h3):(1'h0)] reg2786 = (1'h0);
  reg [(4'he):(1'h0)] reg2785 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2783 = (1'h0);
  reg [(4'hb):(1'h0)] reg2781 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2780 = (1'h0);
  reg [(5'h10):(1'h0)] reg2779 = (1'h0);
  reg [(3'h6):(1'h0)] reg2778 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2777 = (1'h0);
  reg [(4'ha):(1'h0)] reg2775 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2725 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2716 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2772 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2771 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2770 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2769 = (1'h0);
  reg [(3'h7):(1'h0)] reg2768 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2766 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2765 = (1'h0);
  reg [(4'hf):(1'h0)] reg2764 = (1'h0);
  reg [(3'h6):(1'h0)] reg2763 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2762 = (1'h0);
  reg [(2'h2):(1'h0)] reg2755 = (1'h0);
  reg [(4'h9):(1'h0)] reg2753 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2761 = (1'h0);
  reg [(4'h8):(1'h0)] reg2760 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2759 = (1'h0);
  reg [(4'ha):(1'h0)] reg2758 = (1'h0);
  reg [(4'hc):(1'h0)] reg2757 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2756 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2754 = (1'h0);
  reg [(3'h4):(1'h0)] reg2752 = (1'h0);
  reg [(4'h8):(1'h0)] reg2751 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2750 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2749 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2748 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2747 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2746 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2744 = (1'h0);
  reg [(3'h5):(1'h0)] reg2743 = (1'h0);
  reg [(3'h7):(1'h0)] reg2742 = (1'h0);
  reg [(4'hb):(1'h0)] reg2740 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2739 = (1'h0);
  reg [(3'h5):(1'h0)] reg2738 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2737 = (1'h0);
  reg [(2'h3):(1'h0)] reg2735 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2734 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2733 = (1'h0);
  reg [(3'h6):(1'h0)] reg2732 = (1'h0);
  reg [(3'h7):(1'h0)] reg2731 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2709 = (1'h0);
  reg [(2'h3):(1'h0)] reg2708 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2729 = (1'h0);
  reg [(4'h9):(1'h0)] reg2728 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2727 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2726 = (1'h0);
  reg [(3'h6):(1'h0)] reg2724 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2723 = (1'h0);
  reg [(2'h3):(1'h0)] reg2722 = (1'h0);
  reg [(3'h7):(1'h0)] reg2721 = (1'h0);
  reg [(2'h3):(1'h0)] reg2720 = (1'h0);
  reg [(2'h2):(1'h0)] reg2719 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2718 = (1'h0);
  reg [(4'hf):(1'h0)] reg2717 = (1'h0);
  reg [(3'h5):(1'h0)] reg2715 = (1'h0);
  reg [(4'ha):(1'h0)] reg2714 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2713 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2712 = (1'h0);
  reg [(2'h2):(1'h0)] reg2711 = (1'h0);
  reg [(2'h3):(1'h0)] reg2710 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1197 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1198 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1199 = (1'h0);
  reg [(2'h3):(1'h0)] reg1200 = (1'h0);
  reg [(4'hb):(1'h0)] reg1202 = (1'h0);
  reg [(5'h10):(1'h0)] reg1203 = (1'h0);
  reg [(3'h6):(1'h0)] reg1205 = (1'h0);
  reg [(4'he):(1'h0)] reg1208 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1209 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1210 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1213 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1214 = (1'h0);
  reg [(3'h7):(1'h0)] reg1215 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1216 = (1'h0);
  reg [(4'hb):(1'h0)] reg1217 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1219 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1220 = (1'h0);
  reg [(4'h9):(1'h0)] reg1222 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1223 = (1'h0);
  reg [(3'h6):(1'h0)] reg1224 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1226 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1227 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1228 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1229 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1230 = (1'h0);
  reg [(3'h4):(1'h0)] reg1232 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1233 = (1'h0);
  reg [(3'h6):(1'h0)] reg1234 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1235 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1237 = (1'h0);
  reg [(3'h7):(1'h0)] reg1238 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1239 = (1'h0);
  reg [(4'hb):(1'h0)] reg1240 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3207 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3198 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3192 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3220 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3219 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3211 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3208 = (1'h0);
  reg [(4'he):(1'h0)] forvar3209 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3193 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3202 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3196 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3179 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3178 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3173 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3170 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3169 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3160 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3158 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3152 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3148 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3147 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3146 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3145 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3140 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3136 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3135 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3134 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3079 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3076 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3067 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3065 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3122 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3118 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3117 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3105 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3102 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3101 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3100 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3097 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3090 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3081 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3078 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3083 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3082 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3077 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3072 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3066 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3060 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3052 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3070 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3068 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3071 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3069 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3062 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3058 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3051 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3046 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3039 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3034 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3028 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3032 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3043 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3042 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3038 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3036 = (1'h0);
  reg [(4'he):(1'h0)] forvar3035 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3033 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3025 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3024 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3023 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2999 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2998 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3001 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3000 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2994 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2990 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2989 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2979 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2970 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2976 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2963 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3011 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3013 = (1'h0);
  reg [(4'he):(1'h0)] forvar3007 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2996 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2995 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2991 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2987 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2984 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2978 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2977 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2965 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2964 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2962 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2915 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2914 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2902 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2901 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2959 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2952 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2948 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2944 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2941 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2933 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2932 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2930 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2927 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2926 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2920 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2918 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2917 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2912 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2908 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2899 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2906 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2904 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2903 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2898 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2891 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2890 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2887 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2881 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2876 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2875 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2874 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2872 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2862 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2857 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2853 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2850 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2843 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2838 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2864 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2861 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2860 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2859 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2855 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2852 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2851 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2846 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2845 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2840 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2839 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2832 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2820 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2825 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2821 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2819 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2810 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2816 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2812 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2809 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2798 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2796 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2804 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2794 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2792 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2789 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2784 = (1'h0);
  reg [(4'he):(1'h0)] forvar2782 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2776 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2774 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2773 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2711 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2723 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2715 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2710 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2767 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2763 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2758 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2754 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2755 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2753 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2745 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2741 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2736 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2730 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2712 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2725 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2716 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2709 = (1'h0);
  reg [(4'he):(1'h0)] forvar2708 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1236 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1231 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1225 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1221 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1218 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1212 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1211 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1207 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1206 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1204 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1201 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1196 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1195 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1194 = (1'h0);
  assign y = {wire3223,
                 wire3021,
                 wire2837,
                 wire1192,
                 wire1193,
                 wire1241,
                 wire2706,
                 reg3222,
                 reg3221,
                 reg3209,
                 reg3218,
                 reg3217,
                 reg3216,
                 reg3215,
                 reg3214,
                 reg3213,
                 reg3212,
                 reg3211,
                 reg3210,
                 reg3208,
                 reg3207,
                 reg3206,
                 reg3202,
                 reg3205,
                 reg3204,
                 reg3203,
                 reg3201,
                 reg3200,
                 reg3199,
                 reg3198,
                 reg3197,
                 reg3195,
                 reg3194,
                 reg3193,
                 reg3192,
                 reg3191,
                 reg3190,
                 reg3189,
                 reg3188,
                 reg3187,
                 reg3186,
                 reg3185,
                 reg3184,
                 reg3183,
                 reg3182,
                 reg3181,
                 reg3180,
                 reg3177,
                 reg3176,
                 reg3175,
                 reg3174,
                 reg3172,
                 reg3171,
                 reg3170,
                 reg3168,
                 reg3167,
                 reg3166,
                 reg3165,
                 reg3164,
                 reg3163,
                 reg3162,
                 reg3161,
                 reg3159,
                 reg3157,
                 reg3156,
                 reg3155,
                 reg3154,
                 reg3153,
                 reg3151,
                 reg3150,
                 reg3149,
                 reg3144,
                 reg3143,
                 reg3142,
                 reg3141,
                 reg3139,
                 reg3138,
                 reg3137,
                 reg3133,
                 reg3062,
                 reg3058,
                 reg3132,
                 reg3131,
                 reg3130,
                 reg3129,
                 reg3128,
                 reg3127,
                 reg3126,
                 reg3125,
                 reg3124,
                 reg3123,
                 reg3121,
                 reg3120,
                 reg3119,
                 reg3116,
                 reg3115,
                 reg3114,
                 reg3113,
                 reg3112,
                 reg3111,
                 reg3110,
                 reg3109,
                 reg3108,
                 reg3107,
                 reg3106,
                 reg3104,
                 reg3103,
                 reg3099,
                 reg3098,
                 reg3096,
                 reg3095,
                 reg3094,
                 reg3093,
                 reg3092,
                 reg3091,
                 reg3089,
                 reg3088,
                 reg3087,
                 reg3086,
                 reg3085,
                 reg3083,
                 reg3082,
                 reg3084,
                 reg3081,
                 reg3080,
                 reg3079,
                 reg3078,
                 reg3076,
                 reg3075,
                 reg3074,
                 reg3051,
                 reg3071,
                 reg3069,
                 reg3073,
                 reg3072,
                 reg3070,
                 reg3068,
                 reg3067,
                 reg3066,
                 reg3065,
                 reg3064,
                 reg3063,
                 reg3061,
                 reg3060,
                 reg3059,
                 reg3057,
                 reg3056,
                 reg3055,
                 reg3054,
                 reg3053,
                 reg3052,
                 reg3050,
                 reg3049,
                 reg3048,
                 reg3043,
                 reg3042,
                 reg3036,
                 reg3023,
                 reg3038,
                 reg3035,
                 reg3033,
                 reg3047,
                 reg3046,
                 reg3045,
                 reg3044,
                 reg3041,
                 reg3040,
                 reg3039,
                 reg3037,
                 reg3034,
                 reg3032,
                 reg3024,
                 reg3031,
                 reg3030,
                 reg3029,
                 reg3028,
                 reg3027,
                 reg3026,
                 reg3025,
                 reg3022,
                 reg2996,
                 reg2995,
                 reg2984,
                 reg2962,
                 reg2977,
                 reg2965,
                 reg2964,
                 reg3020,
                 reg2991,
                 reg3019,
                 reg3018,
                 reg3017,
                 reg3013,
                 reg3007,
                 reg3016,
                 reg3015,
                 reg3014,
                 reg3012,
                 reg3011,
                 reg3010,
                 reg3009,
                 reg3008,
                 reg3006,
                 reg3005,
                 reg3004,
                 reg3003,
                 reg3002,
                 reg3001,
                 reg3000,
                 reg2999,
                 reg2998,
                 reg2997,
                 reg2994,
                 reg2993,
                 reg2992,
                 reg2987,
                 reg2990,
                 reg2989,
                 reg2988,
                 reg2986,
                 reg2985,
                 reg2983,
                 reg2982,
                 reg2981,
                 reg2980,
                 reg2979,
                 reg2976,
                 reg2975,
                 reg2974,
                 reg2973,
                 reg2972,
                 reg2971,
                 reg2970,
                 reg2969,
                 reg2968,
                 reg2967,
                 reg2966,
                 reg2963,
                 reg2917,
                 reg2961,
                 reg2960,
                 reg2930,
                 reg2958,
                 reg2957,
                 reg2956,
                 reg2955,
                 reg2954,
                 reg2953,
                 reg2951,
                 reg2950,
                 reg2949,
                 reg2947,
                 reg2946,
                 reg2945,
                 reg2943,
                 reg2942,
                 reg2940,
                 reg2939,
                 reg2938,
                 reg2937,
                 reg2936,
                 reg2935,
                 reg2934,
                 reg2931,
                 reg2918,
                 reg2929,
                 reg2928,
                 reg2927,
                 reg2926,
                 reg2925,
                 reg2924,
                 reg2923,
                 reg2922,
                 reg2921,
                 reg2920,
                 reg2919,
                 reg2916,
                 reg2915,
                 reg2906,
                 reg2904,
                 reg2903,
                 reg2914,
                 reg2913,
                 reg2912,
                 reg2911,
                 reg2910,
                 reg2909,
                 reg2908,
                 reg2907,
                 reg2905,
                 reg2902,
                 reg2901,
                 reg2900,
                 reg2899,
                 reg2897,
                 reg2896,
                 reg2895,
                 reg2894,
                 reg2893,
                 reg2892,
                 reg2891,
                 reg2889,
                 reg2888,
                 reg2886,
                 reg2885,
                 reg2884,
                 reg2883,
                 reg2882,
                 reg2880,
                 reg2879,
                 reg2878,
                 reg2877,
                 reg2873,
                 reg2864,
                 reg2861,
                 reg2860,
                 reg2859,
                 reg2855,
                 reg2852,
                 reg2851,
                 reg2846,
                 reg2845,
                 reg2840,
                 reg2839,
                 reg2871,
                 reg2870,
                 reg2869,
                 reg2868,
                 reg2867,
                 reg2866,
                 reg2865,
                 reg2863,
                 reg2862,
                 reg2858,
                 reg2857,
                 reg2856,
                 reg2854,
                 reg2853,
                 reg2850,
                 reg2849,
                 reg2848,
                 reg2847,
                 reg2844,
                 reg2843,
                 reg2842,
                 reg2841,
                 reg2838,
                 reg2836,
                 reg2835,
                 reg2834,
                 reg2833,
                 reg2831,
                 reg2830,
                 reg2829,
                 reg2825,
                 reg2821,
                 reg2819,
                 reg2828,
                 reg2827,
                 reg2826,
                 reg2824,
                 reg2823,
                 reg2822,
                 reg2820,
                 reg2812,
                 reg2818,
                 reg2817,
                 reg2815,
                 reg2814,
                 reg2813,
                 reg2811,
                 reg2810,
                 reg2808,
                 reg2807,
                 reg2806,
                 reg2805,
                 reg2803,
                 reg2802,
                 reg2801,
                 reg2800,
                 reg2799,
                 reg2798,
                 reg2797,
                 reg2796,
                 reg2795,
                 reg2784,
                 reg2793,
                 reg2791,
                 reg2790,
                 reg2788,
                 reg2787,
                 reg2786,
                 reg2785,
                 reg2783,
                 reg2781,
                 reg2780,
                 reg2779,
                 reg2778,
                 reg2777,
                 reg2775,
                 reg2725,
                 reg2716,
                 reg2772,
                 reg2771,
                 reg2770,
                 reg2769,
                 reg2768,
                 reg2766,
                 reg2765,
                 reg2764,
                 reg2763,
                 reg2762,
                 reg2755,
                 reg2753,
                 reg2761,
                 reg2760,
                 reg2759,
                 reg2758,
                 reg2757,
                 reg2756,
                 reg2754,
                 reg2752,
                 reg2751,
                 reg2750,
                 reg2749,
                 reg2748,
                 reg2747,
                 reg2746,
                 reg2744,
                 reg2743,
                 reg2742,
                 reg2740,
                 reg2739,
                 reg2738,
                 reg2737,
                 reg2735,
                 reg2734,
                 reg2733,
                 reg2732,
                 reg2731,
                 reg2709,
                 reg2708,
                 reg2729,
                 reg2728,
                 reg2727,
                 reg2726,
                 reg2724,
                 reg2723,
                 reg2722,
                 reg2721,
                 reg2720,
                 reg2719,
                 reg2718,
                 reg2717,
                 reg2715,
                 reg2714,
                 reg2713,
                 reg2712,
                 reg2711,
                 reg2710,
                 reg1197,
                 reg1198,
                 reg1199,
                 reg1200,
                 reg1202,
                 reg1203,
                 reg1205,
                 reg1208,
                 reg1209,
                 reg1210,
                 reg1213,
                 reg1214,
                 reg1215,
                 reg1216,
                 reg1217,
                 reg1219,
                 reg1220,
                 reg1222,
                 reg1223,
                 reg1224,
                 reg1226,
                 reg1227,
                 reg1228,
                 reg1229,
                 reg1230,
                 reg1232,
                 reg1233,
                 reg1234,
                 reg1235,
                 reg1237,
                 reg1238,
                 reg1239,
                 reg1240,
                 forvar3207,
                 forvar3198,
                 forvar3192,
                 forvar3220,
                 forvar3219,
                 forvar3211,
                 forvar3208,
                 forvar3209,
                 forvar3193,
                 forvar3202,
                 forvar3196,
                 forvar3179,
                 forvar3178,
                 forvar3173,
                 forvar3170,
                 forvar3169,
                 forvar3160,
                 forvar3158,
                 forvar3152,
                 forvar3148,
                 forvar3147,
                 forvar3146,
                 forvar3145,
                 forvar3140,
                 forvar3136,
                 forvar3135,
                 forvar3134,
                 forvar3079,
                 forvar3076,
                 forvar3067,
                 forvar3065,
                 forvar3122,
                 forvar3118,
                 forvar3117,
                 forvar3105,
                 forvar3102,
                 forvar3101,
                 forvar3100,
                 forvar3097,
                 forvar3090,
                 forvar3081,
                 forvar3078,
                 forvar3083,
                 forvar3082,
                 forvar3077,
                 forvar3072,
                 forvar3066,
                 forvar3060,
                 forvar3052,
                 forvar3070,
                 forvar3068,
                 forvar3071,
                 forvar3069,
                 forvar3062,
                 forvar3058,
                 forvar3051,
                 forvar3046,
                 forvar3039,
                 forvar3034,
                 forvar3028,
                 forvar3032,
                 forvar3043,
                 forvar3042,
                 forvar3038,
                 forvar3036,
                 forvar3035,
                 forvar3033,
                 forvar3025,
                 forvar3024,
                 forvar3023,
                 forvar2999,
                 forvar2998,
                 forvar3001,
                 forvar3000,
                 forvar2994,
                 forvar2990,
                 forvar2989,
                 forvar2979,
                 forvar2970,
                 forvar2976,
                 forvar2963,
                 forvar3011,
                 forvar3013,
                 forvar3007,
                 forvar2996,
                 forvar2995,
                 forvar2991,
                 forvar2987,
                 forvar2984,
                 forvar2978,
                 forvar2977,
                 forvar2965,
                 forvar2964,
                 forvar2962,
                 forvar2915,
                 forvar2914,
                 forvar2902,
                 forvar2901,
                 forvar2959,
                 forvar2952,
                 forvar2948,
                 forvar2944,
                 forvar2941,
                 forvar2933,
                 forvar2932,
                 forvar2930,
                 forvar2927,
                 forvar2926,
                 forvar2920,
                 forvar2918,
                 forvar2917,
                 forvar2912,
                 forvar2908,
                 forvar2899,
                 forvar2906,
                 forvar2904,
                 forvar2903,
                 forvar2898,
                 forvar2891,
                 forvar2890,
                 forvar2887,
                 forvar2881,
                 forvar2876,
                 forvar2875,
                 forvar2874,
                 forvar2872,
                 forvar2862,
                 forvar2857,
                 forvar2853,
                 forvar2850,
                 forvar2843,
                 forvar2838,
                 forvar2864,
                 forvar2861,
                 forvar2860,
                 forvar2859,
                 forvar2855,
                 forvar2852,
                 forvar2851,
                 forvar2846,
                 forvar2845,
                 forvar2840,
                 forvar2839,
                 forvar2832,
                 forvar2820,
                 forvar2825,
                 forvar2821,
                 forvar2819,
                 forvar2810,
                 forvar2816,
                 forvar2812,
                 forvar2809,
                 forvar2798,
                 forvar2796,
                 forvar2804,
                 forvar2794,
                 forvar2792,
                 forvar2789,
                 forvar2784,
                 forvar2782,
                 forvar2776,
                 forvar2774,
                 forvar2773,
                 forvar2711,
                 forvar2723,
                 forvar2715,
                 forvar2710,
                 forvar2767,
                 forvar2763,
                 forvar2758,
                 forvar2754,
                 forvar2755,
                 forvar2753,
                 forvar2745,
                 forvar2741,
                 forvar2736,
                 forvar2730,
                 forvar2712,
                 forvar2725,
                 forvar2716,
                 forvar2709,
                 forvar2708,
                 forvar1236,
                 forvar1231,
                 forvar1225,
                 forvar1221,
                 forvar1218,
                 forvar1212,
                 forvar1211,
                 forvar1207,
                 forvar1206,
                 forvar1204,
                 forvar1201,
                 forvar1196,
                 forvar1195,
                 forvar1194,
                 (1'h0)};
  assign wire1192 = (^({$unsigned(wire1191)} ?
                        {wire1187[(2'h2):(1'h0)]} : $signed((wire1187 ^~ wire1189))));
  assign wire1193 = wire1190[(3'h6):(3'h4)];
  always
    @(posedge clk) begin
      for (forvar1194 = (1'h0); (forvar1194 < (2'h2)); forvar1194 = (forvar1194 + (1'h1)))
        begin
          for (forvar1195 = (1'h0); (forvar1195 < (2'h2)); forvar1195 = (forvar1195 + (1'h1)))
            begin
              if ((((~|$signed((8'h9f))) ?
                      forvar1195[(4'h8):(1'h1)] : ((8'hae) ?
                          $unsigned(forvar1195) : {(8'hb1)})) ?
                  wire1193[(3'h4):(3'h4)] : wire1190[(4'hd):(2'h2)]))
                begin
                  for (forvar1196 = (1'h0); (forvar1196 < (1'h1)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 <= (wire1193 ?
                          wire1193[(2'h3):(1'h1)] : {({forvar1194} ?
                                  wire1191[(4'h9):(3'h4)] : (forvar1194 ?
                                      (8'ha8) : (8'ha7)))});
                      reg1198 <= ($signed(((wire1188 ?
                              reg1197 : (8'hb2)) && wire1191)) ?
                          (reg1197 ~^ (~^(forvar1195 - wire1189))) : $signed(reg1197));
                      reg1199 <= ($signed(($unsigned(wire1193) >> forvar1195[(1'h1):(1'h1)])) ?
                          $signed(((&wire1187) ?
                              forvar1196 : $unsigned(wire1188))) : wire1192[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar1196 = (1'h0); (forvar1196 < (1'h1)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 <= $unsigned({forvar1195[(1'h1):(1'h0)]});
                      reg1198 <= forvar1194[(4'h9):(3'h7)];
                      reg1199 <= $unsigned(((~forvar1195) ?
                          {$unsigned(wire1189)} : ({wire1188} ?
                              wire1193[(1'h1):(1'h1)] : (wire1193 ?
                                  wire1188 : reg1198))));
                      reg1200 <= (($signed($signed((8'ha4))) ?
                              ({forvar1196} ?
                                  ((8'hb7) || wire1193) : ((8'haf) ?
                                      wire1189 : reg1199)) : $signed(reg1198[(4'ha):(4'ha)])) ?
                          $signed({$unsigned((8'ha1))}) : (((wire1190 <= forvar1194) ^~ $unsigned((8'hac))) <<< forvar1196));
                    end
                  for (forvar1201 = (1'h0); (forvar1201 < (2'h3)); forvar1201 = (forvar1201 + (1'h1)))
                    begin
                      reg1202 <= forvar1195;
                      reg1203 <= (($signed((forvar1196 ?
                              reg1202 : wire1192)) ~^ {{forvar1194}}) ?
                          (^$signed(wire1193[(2'h2):(1'h0)])) : reg1197);
                    end
                  for (forvar1204 = (1'h0); (forvar1204 < (1'h1)); forvar1204 = (forvar1204 + (1'h1)))
                    begin
                      reg1205 <= forvar1196;
                    end
                end
              for (forvar1206 = (1'h0); (forvar1206 < (2'h2)); forvar1206 = (forvar1206 + (1'h1)))
                begin
                  for (forvar1207 = (1'h0); (forvar1207 < (1'h1)); forvar1207 = (forvar1207 + (1'h1)))
                    begin
                      reg1208 <= {reg1197[(3'h6):(2'h2)]};
                      reg1209 <= {$signed(reg1200[(1'h1):(1'h0)])};
                      reg1210 <= $signed({(8'hb7)});
                    end
                end
              for (forvar1211 = (1'h0); (forvar1211 < (1'h0)); forvar1211 = (forvar1211 + (1'h1)))
                begin
                  for (forvar1212 = (1'h0); (forvar1212 < (1'h1)); forvar1212 = (forvar1212 + (1'h1)))
                    begin
                      reg1213 <= $unsigned({forvar1206[(1'h0):(1'h0)]});
                    end
                  if ((8'hb5))
                    begin
                      reg1214 <= (~((!$signed((8'ha3))) ?
                          $signed((forvar1206 ?
                              forvar1206 : reg1203)) : $unsigned((wire1191 <<< forvar1206))));
                      reg1215 <= (~^$signed((+(forvar1212 ?
                          forvar1194 : (8'hb7)))));
                      reg1216 <= forvar1211[(4'h9):(4'h8)];
                      reg1217 <= ($signed(forvar1207[(2'h2):(1'h0)]) ?
                          $unsigned($signed($signed(forvar1212))) : reg1210[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg1214 <= wire1187[(1'h1):(1'h1)];
                      reg1215 <= (reg1203[(3'h4):(3'h4)] ?
                          (|$unsigned(forvar1195)) : $signed($unsigned((forvar1201 ?
                              reg1203 : forvar1196))));
                    end
                  for (forvar1218 = (1'h0); (forvar1218 < (1'h0)); forvar1218 = (forvar1218 + (1'h1)))
                    begin
                      reg1219 <= ((~&$unsigned($unsigned(forvar1195))) ?
                          (8'h9f) : (((reg1209 ?
                                  forvar1206 : reg1202) <= (8'h9d)) ?
                              (~|$signed(forvar1195)) : wire1188));
                      reg1220 <= reg1217[(2'h3):(2'h2)];
                    end
                  for (forvar1221 = (1'h0); (forvar1221 < (2'h2)); forvar1221 = (forvar1221 + (1'h1)))
                    begin
                      reg1222 <= $unsigned($unsigned((8'h9c)));
                      reg1223 <= $signed($unsigned(reg1209));
                      reg1224 <= reg1220;
                    end
                end
              for (forvar1225 = (1'h0); (forvar1225 < (1'h1)); forvar1225 = (forvar1225 + (1'h1)))
                begin
                  if ((~&(reg1200[(2'h2):(1'h0)] & {$unsigned((8'haf))})))
                    begin
                      reg1226 <= wire1189[(3'h6):(1'h1)];
                      reg1227 <= wire1190;
                      reg1228 <= $unsigned(wire1191[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg1226 <= wire1192;
                      reg1227 <= $signed(wire1188[(3'h7):(2'h3)]);
                    end
                  if ($signed({forvar1194[(2'h2):(1'h0)]}))
                    begin
                      reg1229 <= wire1191;
                      reg1230 <= (reg1198[(4'hd):(4'h8)] > (&$signed((8'hb3))));
                    end
                  else
                    begin
                      reg1229 <= $signed(((^~(8'hb2)) << $unsigned(reg1203[(3'h7):(3'h7)])));
                    end
                end
            end
          for (forvar1231 = (1'h0); (forvar1231 < (2'h2)); forvar1231 = (forvar1231 + (1'h1)))
            begin
              if (((~&$signed($signed(reg1219))) < $unsigned(($signed(forvar1218) ?
                  $unsigned(forvar1231) : (~|forvar1206)))))
                begin
                  if (reg1205[(3'h4):(2'h3)])
                    begin
                      reg1232 <= ($unsigned($signed(forvar1218)) ?
                          {forvar1231} : (^~(reg1215[(1'h1):(1'h1)] ?
                              $unsigned(reg1216) : (reg1227 ?
                                  wire1188 : reg1214))));
                    end
                  else
                    begin
                      reg1232 <= forvar1221[(4'hb):(4'h9)];
                      reg1233 <= $signed((8'ha6));
                      reg1234 <= (&$signed($signed($signed(reg1222))));
                    end
                end
              else
                begin
                  if (reg1203)
                    begin
                      reg1232 <= ($signed({$unsigned(forvar1231)}) ?
                          {reg1205[(2'h2):(1'h1)]} : (~^((reg1227 ?
                                  reg1219 : forvar1211) ?
                              reg1219 : ((8'hb2) ? forvar1206 : (8'hab)))));
                      reg1233 <= {(8'h9d)};
                    end
                  else
                    begin
                      reg1232 <= (8'hb0);
                      reg1233 <= $signed(((~&reg1217) ?
                          (!$signed(wire1190)) : (reg1232 & wire1187)));
                      reg1234 <= $unsigned($unsigned($signed($signed(wire1190))));
                      reg1235 <= $unsigned({reg1208[(4'h8):(1'h0)]});
                    end
                  for (forvar1236 = (1'h0); (forvar1236 < (1'h0)); forvar1236 = (forvar1236 + (1'h1)))
                    begin
                      reg1237 <= $signed($signed((reg1233[(2'h2):(1'h0)] ~^ $unsigned(reg1216))));
                    end
                  if (reg1203[(4'he):(4'h8)])
                    begin
                      reg1238 <= {forvar1225[(4'ha):(1'h1)]};
                    end
                  else
                    begin
                      reg1238 <= forvar1196;
                      reg1239 <= (8'had);
                    end
                  reg1240 <= $unsigned(forvar1201);
                end
            end
        end
    end
  assign wire1241 = (reg1198[(4'he):(3'h5)] - reg1203);
  module1242 #() modinst2707 (.wire1244(wire1190), .wire1246(reg1226), .clk(clk), .wire1245(reg1197), .y(wire2706), .wire1243(reg1240));
  always
    @(posedge clk) begin
      if ((($signed($signed(reg1227)) < wire1189[(3'h7):(3'h5)]) ?
          $signed(reg1214) : ({reg1199} >= reg1203[(4'he):(3'h7)])))
        begin
          if ($signed(reg1228[(1'h0):(1'h0)]))
            begin
              for (forvar2708 = (1'h0); (forvar2708 < (2'h3)); forvar2708 = (forvar2708 + (1'h1)))
                begin
                  for (forvar2709 = (1'h0); (forvar2709 < (2'h2)); forvar2709 = (forvar2709 + (1'h1)))
                    begin
                      reg2710 <= reg1232[(1'h1):(1'h0)];
                      reg2711 <= $unsigned(reg1202[(4'h9):(3'h7)]);
                    end
                  if ($unsigned($signed((+$unsigned(reg1210)))))
                    begin
                      reg2712 <= $unsigned({({reg1199} ?
                              (wire1193 ? (8'ha6) : reg1232) : (|reg1214))});
                      reg2713 <= reg1230;
                      reg2714 <= (~|(((8'hab) >> {wire1188}) ?
                          $signed($signed(wire1192)) : (!(reg1226 ?
                              (8'hb9) : forvar2708))));
                      reg2715 <= (~^(((8'hb0) ?
                              (reg1224 ?
                                  (8'hb0) : reg1223) : reg1199[(3'h4):(3'h4)]) ?
                          reg1226 : $signed(((8'haa) ^ reg1237))));
                    end
                  else
                    begin
                      reg2712 <= $unsigned(reg1228[(2'h2):(1'h1)]);
                      reg2713 <= (8'hba);
                      reg2714 <= reg1227;
                    end
                  for (forvar2716 = (1'h0); (forvar2716 < (2'h3)); forvar2716 = (forvar2716 + (1'h1)))
                    begin
                      reg2717 <= (-(reg1205 <= reg1217[(2'h2):(1'h1)]));
                      reg2718 <= (reg2713 ?
                          (8'hae) : $signed($unsigned((reg1209 >> reg1223))));
                      reg2719 <= reg2714[(3'h4):(2'h2)];
                      reg2720 <= $unsigned((!(reg1214 || {reg1213})));
                    end
                  if ($unsigned(wire1188))
                    begin
                      reg2721 <= (~^$signed((forvar2709 == wire2706[(1'h0):(1'h0)])));
                      reg2722 <= {reg1217[(3'h6):(2'h3)]};
                      reg2723 <= reg1208;
                      reg2724 <= (reg1215 ?
                          (^reg2710) : (~|((reg1232 ^~ (8'ha7)) ?
                              ((8'hb3) && reg1205) : {reg1219})));
                    end
                  else
                    begin
                      reg2721 <= reg2713;
                      reg2722 <= ({((wire1191 ? wire1188 : reg1227) ?
                                  $signed(forvar2709) : $signed(reg1203))} ?
                          $signed(((reg1227 ?
                              wire1192 : reg1210) ^ $unsigned(reg1202))) : {$signed((8'ha0))});
                    end
                end
              for (forvar2725 = (1'h0); (forvar2725 < (1'h1)); forvar2725 = (forvar2725 + (1'h1)))
                begin
                  if ((($signed(reg1234[(1'h0):(1'h0)]) ?
                      {wire1187} : ({(8'ha9)} >> (!(8'hae)))) | {((reg2712 ?
                          wire1189 : (8'hac)) >> (~&reg1198))}))
                    begin
                      reg2726 <= reg1228[(1'h0):(1'h0)];
                      reg2727 <= reg1202[(3'h6):(2'h3)];
                      reg2728 <= $unsigned({(reg1208[(1'h1):(1'h0)] | (wire1187 ?
                              reg1226 : reg1223))});
                      reg2729 <= (((((8'had) < (8'ha1)) ?
                                  $unsigned(reg1227) : {reg2718}) ?
                              $unsigned((8'h9d)) : ((|reg2727) <= reg1220[(2'h3):(1'h0)])) ?
                          (^$unsigned(reg1199[(3'h4):(2'h3)])) : reg1229[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg2726 <= {reg1219[(1'h1):(1'h0)]};
                      reg2727 <= (reg1234 ? reg2727[(2'h2):(2'h2)] : reg2714);
                      reg2728 <= $signed({wire1190});
                      reg2729 <= reg2711;
                    end
                end
            end
          else
            begin
              if ((+$signed(reg1209)))
                begin
                  if (forvar2725)
                    begin
                      reg2708 <= reg1209[(3'h4):(2'h2)];
                      reg2709 <= {((~^((8'hba) ^ reg1227)) ?
                              ((reg2723 ? reg2719 : reg1228) ?
                                  (reg1240 * reg1202) : (reg2711 ?
                                      wire2706 : reg1220)) : $unsigned((~^wire1188)))};
                      reg2710 <= $unsigned($unsigned($signed({reg1216})));
                    end
                  else
                    begin
                      reg2708 <= ((((wire1187 || reg1223) ?
                              reg2728[(3'h5):(2'h3)] : reg1226) ?
                          (reg2724 ?
                              reg2724 : (forvar2708 - (8'ha0))) : (~^{reg2727})) > reg2708);
                    end
                  reg2711 <= forvar2725[(3'h7):(3'h4)];
                end
              else
                begin
                  for (forvar2708 = (1'h0); (forvar2708 < (2'h2)); forvar2708 = (forvar2708 + (1'h1)))
                    begin
                      reg2709 <= $signed(($unsigned(reg2721[(2'h3):(2'h2)]) * wire1190[(2'h2):(1'h0)]));
                    end
                end
              if (reg1226)
                begin
                  for (forvar2712 = (1'h0); (forvar2712 < (2'h2)); forvar2712 = (forvar2712 + (1'h1)))
                    begin
                      reg2713 <= reg1213;
                    end
                end
              else
                begin
                  for (forvar2712 = (1'h0); (forvar2712 < (2'h3)); forvar2712 = (forvar2712 + (1'h1)))
                    begin
                      reg2713 <= reg2715;
                      reg2714 <= $unsigned(reg1234[(2'h2):(2'h2)]);
                    end
                end
            end
          for (forvar2730 = (1'h0); (forvar2730 < (2'h3)); forvar2730 = (forvar2730 + (1'h1)))
            begin
              if ({(^reg2721)})
                begin
                  if ($unsigned((8'hb9)))
                    begin
                      reg2731 <= (8'hb4);
                      reg2732 <= reg2719[(2'h2):(1'h1)];
                      reg2733 <= $unsigned(reg1205);
                    end
                  else
                    begin
                      reg2731 <= (~(($signed(wire1190) ?
                          $unsigned(reg2717) : reg1232[(2'h3):(1'h0)]) ^ forvar2725));
                      reg2732 <= {(~($unsigned(reg2728) ?
                              reg1224[(1'h1):(1'h1)] : (reg1222 ?
                                  reg2714 : wire1191)))};
                      reg2733 <= $signed({(~&(reg2711 ? wire1191 : reg1222))});
                    end
                end
              else
                begin
                  reg2731 <= reg1228;
                  if (((((~|reg1208) <= (reg1198 & (8'ha7))) ^ wire1241) < ($signed((reg1197 ?
                          (8'hb1) : (8'hb4))) ?
                      reg2723[(1'h1):(1'h1)] : reg1203)))
                    begin
                      reg2732 <= (8'hb9);
                    end
                  else
                    begin
                      reg2732 <= (|$unsigned(reg2724[(3'h5):(3'h5)]));
                      reg2733 <= $signed((-($signed(reg1224) ?
                          reg2711[(1'h1):(1'h1)] : $signed(reg1220))));
                      reg2734 <= (^~({((8'ha1) ?
                              wire1190 : reg2715)} >>> $unsigned((reg1234 <= wire1193))));
                      reg2735 <= (^(((reg1222 + wire1241) ~^ (reg1202 ?
                          (8'ha3) : forvar2725)) && $unsigned((reg1202 ?
                          (8'hba) : reg1205))));
                    end
                  for (forvar2736 = (1'h0); (forvar2736 < (1'h0)); forvar2736 = (forvar2736 + (1'h1)))
                    begin
                      reg2737 <= reg2710[(2'h3):(2'h3)];
                      reg2738 <= $signed($unsigned(reg1228));
                      reg2739 <= reg1223[(2'h3):(1'h0)];
                      reg2740 <= $signed((-({reg2712} >>> $unsigned(reg2726))));
                    end
                end
              for (forvar2741 = (1'h0); (forvar2741 < (2'h2)); forvar2741 = (forvar2741 + (1'h1)))
                begin
                  reg2742 <= $signed($signed(((^~reg2739) ?
                      $unsigned(wire1188) : $signed(reg1202))));
                  if ((((~|reg1232[(2'h3):(1'h0)]) <= ((wire1191 ?
                      reg2734 : wire1241) <= $signed(reg2712))) >>> reg1237[(2'h3):(2'h3)]))
                    begin
                      reg2743 <= (~|$signed(forvar2709));
                      reg2744 <= ((!wire1190[(4'ha):(2'h3)]) ?
                          {reg2738[(2'h3):(1'h0)]} : $unsigned($unsigned((reg2739 == reg2710))));
                    end
                  else
                    begin
                      reg2743 <= (&{wire1193[(2'h3):(1'h1)]});
                      reg2744 <= $unsigned((reg1237 ? reg2737 : (|reg2710)));
                    end
                  for (forvar2745 = (1'h0); (forvar2745 < (2'h2)); forvar2745 = (forvar2745 + (1'h1)))
                    begin
                      reg2746 <= reg2721;
                      reg2747 <= $unsigned((+$signed(reg2715)));
                      reg2748 <= (!$signed($unsigned((^~reg1197))));
                    end
                  if ((-reg1220))
                    begin
                      reg2749 <= (&(!reg2733[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg2749 <= reg1203;
                    end
                end
              reg2750 <= reg1229;
              reg2751 <= (($signed(reg1228[(3'h4):(2'h2)]) != {{forvar2716}}) ?
                  ((reg1223[(1'h1):(1'h1)] ?
                      (+reg2711) : (!(8'hb9))) || ($unsigned(reg1215) ?
                      (reg2739 ?
                          reg1208 : reg2721) : forvar2745[(1'h0):(1'h0)])) : (reg1238[(2'h2):(2'h2)] ?
                      (!$unsigned(reg2708)) : reg2738[(3'h5):(3'h5)]));
            end
          reg2752 <= (({reg2724} ?
              ($unsigned(reg2749) && $unsigned(reg2727)) : wire1189) || $signed($unsigned({forvar2708})));
          if ($unsigned((8'ha0)))
            begin
              for (forvar2753 = (1'h0); (forvar2753 < (2'h3)); forvar2753 = (forvar2753 + (1'h1)))
                begin
                  reg2754 <= ($signed($unsigned($unsigned((8'hb9)))) <<< ($unsigned((^reg1229)) ?
                      (reg2729 >>> (|wire1241)) : ((|reg1200) ?
                          {reg2738} : (!reg1205))));
                  for (forvar2755 = (1'h0); (forvar2755 < (1'h0)); forvar2755 = (forvar2755 + (1'h1)))
                    begin
                      reg2756 <= $signed($signed((forvar2716[(3'h4):(1'h0)] + $signed(reg2729))));
                      reg2757 <= $signed(reg1238);
                    end
                  if ((wire1189[(1'h0):(1'h0)] > forvar2741))
                    begin
                      reg2758 <= (~&reg2723);
                      reg2759 <= $signed($unsigned(((reg2733 ?
                          reg1210 : (8'ha0)) >>> $signed(reg2726))));
                      reg2760 <= (8'h9f);
                    end
                  else
                    begin
                      reg2758 <= reg1223[(1'h1):(1'h1)];
                      reg2759 <= (^(((reg1222 < reg1229) << ((8'hb5) ?
                              reg2752 : reg2750)) ?
                          (-{reg2733}) : reg2722));
                      reg2760 <= $signed((~&reg2749));
                      reg2761 <= ((($signed(wire1188) <= $unsigned(forvar2755)) ?
                              (forvar2709[(4'hd):(4'hc)] <<< $unsigned(reg1205)) : (!$unsigned((8'hb5)))) ?
                          $unsigned(forvar2725[(3'h7):(2'h2)]) : $signed({(&forvar2745)}));
                    end
                end
            end
          else
            begin
              reg2753 <= (~{({reg1228} <<< reg1237)});
              if ({($unsigned(reg2738) + (&{reg1234}))})
                begin
                  for (forvar2754 = (1'h0); (forvar2754 < (2'h2)); forvar2754 = (forvar2754 + (1'h1)))
                    begin
                      reg2755 <= reg2729[(1'h0):(1'h0)];
                      reg2756 <= $unsigned(reg1214[(3'h4):(1'h1)]);
                      reg2757 <= ($signed(((reg2750 < (8'h9f)) <= forvar2709)) ?
                          reg2717 : (reg2753[(2'h3):(1'h0)] ?
                              (reg2733[(1'h0):(1'h0)] ?
                                  (reg2758 ?
                                      (8'hba) : reg2709) : $unsigned(wire1192)) : reg2744[(2'h3):(1'h1)]));
                    end
                  if (forvar2736[(2'h2):(1'h0)])
                    begin
                      reg2758 <= $signed({$signed(reg1237)});
                    end
                  else
                    begin
                      reg2758 <= ((reg2709 << (reg2747 - reg2708[(2'h2):(2'h2)])) ?
                          $unsigned($signed(reg1200)) : ($signed($unsigned((8'ha8))) ?
                              ((reg1228 & reg2722) ^~ $unsigned(forvar2754)) : reg2731));
                      reg2759 <= reg1209[(3'h7):(3'h7)];
                      reg2760 <= (({(forvar2716 ?
                                  reg2761 : reg1237)} >> (reg2734 && ((8'ha1) ?
                              reg2734 : forvar2725))) ?
                          reg1228[(1'h1):(1'h0)] : {(((8'hb0) < reg2727) ?
                                  $signed(reg1233) : ((8'haa) || reg2743))});
                      reg2761 <= (-(8'hb8));
                    end
                  if ((+(reg1224[(3'h5):(2'h2)] <= {reg2744})))
                    begin
                      reg2762 <= ($signed($unsigned((^reg2760))) & reg2753);
                      reg2763 <= $unsigned((^(((8'hb9) ?
                          reg1222 : reg2711) ^ (reg2721 && reg2732))));
                    end
                  else
                    begin
                      reg2762 <= $signed((reg1215 ?
                          (((8'hb1) != reg2763) ?
                              (~(8'haf)) : {(8'ha1)}) : (~|(reg1235 ^~ reg1200))));
                      reg2763 <= ((((^~reg1210) >> reg1217) ^~ $signed((8'ha5))) ~^ (8'ha3));
                    end
                end
              else
                begin
                  if (reg2753[(4'h9):(1'h0)])
                    begin
                      reg2754 <= (reg2746[(3'h7):(2'h2)] && {reg1226});
                      reg2755 <= $signed(reg1197[(4'ha):(3'h5)]);
                    end
                  else
                    begin
                      reg2754 <= (reg1237 ?
                          ((+{reg2746}) ?
                              reg2708 : ($unsigned((8'ha1)) ?
                                  $unsigned(reg2723) : reg2717[(4'hb):(2'h3)])) : (~|((reg2711 + (8'hb2)) - $unsigned(forvar2754))));
                      reg2755 <= reg1240[(4'h8):(2'h2)];
                      reg2756 <= reg2756;
                      reg2757 <= $unsigned(($signed((reg1235 ?
                              reg1228 : (8'hac))) ?
                          (reg2715[(3'h5):(1'h0)] ?
                              (reg2721 <= reg2737) : reg2713) : (reg2723[(3'h6):(2'h2)] == (reg2724 ?
                              reg2737 : reg1214))));
                    end
                  for (forvar2758 = (1'h0); (forvar2758 < (1'h0)); forvar2758 = (forvar2758 + (1'h1)))
                    begin
                      reg2759 <= (wire1188[(1'h1):(1'h0)] != $signed({(reg1209 + reg2743)}));
                      reg2760 <= ((~$signed((~&reg1222))) >= $unsigned($unsigned($signed(reg2754))));
                      reg2761 <= $unsigned($signed(((reg1223 - forvar2758) >> (reg2763 && wire1193))));
                      reg2762 <= ((((~reg1203) << $signed(reg1208)) ?
                              (reg1219[(2'h2):(1'h0)] ?
                                  $signed(forvar2745) : (reg2748 & reg2715)) : reg2737) ?
                          reg2713 : (wire1241 && (-$unsigned((8'haf)))));
                    end
                  for (forvar2763 = (1'h0); (forvar2763 < (2'h2)); forvar2763 = (forvar2763 + (1'h1)))
                    begin
                      reg2764 <= $unsigned($unsigned({reg2714}));
                      reg2765 <= (+$signed((reg2756[(1'h1):(1'h0)] ~^ {(8'hb6)})));
                      reg2766 <= $unsigned($unsigned(reg1223[(2'h2):(1'h1)]));
                    end
                  for (forvar2767 = (1'h0); (forvar2767 < (1'h0)); forvar2767 = (forvar2767 + (1'h1)))
                    begin
                      reg2768 <= forvar2709[(5'h10):(1'h1)];
                      reg2769 <= (&reg2708);
                      reg2770 <= ($signed((^~forvar2730[(1'h0):(1'h0)])) ^~ $signed($unsigned($unsigned((8'haf)))));
                      reg2771 <= (reg1234 >> reg1198);
                    end
                end
              reg2772 <= {((~&$signed(reg1198)) - $unsigned($unsigned(reg2737)))};
            end
        end
      else
        begin
          reg2708 <= $unsigned(reg1216);
          reg2709 <= (-wire1191);
          if ($signed((!reg1213[(4'ha):(3'h4)])))
            begin
              for (forvar2710 = (1'h0); (forvar2710 < (1'h1)); forvar2710 = (forvar2710 + (1'h1)))
                begin
                  if (reg2770[(2'h3):(2'h2)])
                    begin
                      reg2711 <= (~^({(forvar2741 > reg1210)} ?
                          (8'hb3) : {reg1233}));
                      reg2712 <= reg1215[(1'h0):(1'h0)];
                      reg2713 <= (+reg2723);
                      reg2714 <= ($signed((~$unsigned(reg2755))) >>> (^~$signed($signed(reg2729))));
                    end
                  else
                    begin
                      reg2711 <= reg1239[(4'hc):(2'h3)];
                      reg2712 <= forvar2754;
                      reg2713 <= ($unsigned(((reg1226 ^~ reg1237) > reg2732)) >> reg2712);
                      reg2714 <= (~|{reg1235[(1'h0):(1'h0)]});
                    end
                end
              for (forvar2715 = (1'h0); (forvar2715 < (2'h2)); forvar2715 = (forvar2715 + (1'h1)))
                begin
                  if ($unsigned((-($signed(reg2764) ?
                      reg1220[(1'h0):(1'h0)] : $signed(reg2750)))))
                    begin
                      reg2716 <= ((^reg2768[(3'h4):(1'h0)]) >= $signed({(reg1200 < (8'hab))}));
                      reg2717 <= $unsigned(reg2718[(1'h0):(1'h0)]);
                      reg2718 <= ($signed(wire1241) ?
                          {((8'hb1) - (reg1216 < (8'hba)))} : reg1215);
                      reg2719 <= (($unsigned(((8'hb0) ~^ reg2709)) > (reg2714 >>> (reg2731 <= (8'hb7)))) ~^ (forvar2715[(4'h8):(3'h7)] + reg1213));
                    end
                  else
                    begin
                      reg2716 <= {(($unsigned(reg2752) ?
                              $signed(wire1241) : (reg2715 ?
                                  forvar2712 : wire2706)) >> ((|reg1203) ?
                              (|reg2750) : forvar2753[(3'h4):(2'h3)]))};
                      reg2717 <= reg1199;
                    end
                end
              if ((-reg2724))
                begin
                  reg2720 <= (~$signed($signed((wire1189 ?
                      reg1229 : reg1227))));
                  if ((reg1233[(2'h2):(1'h0)] == {((-reg2735) ?
                          reg2765[(1'h0):(1'h0)] : (wire1193 & reg2766))}))
                    begin
                      reg2721 <= ($unsigned($unsigned($signed(reg2755))) + reg2715[(1'h1):(1'h0)]);
                      reg2722 <= $signed({(forvar2715[(4'h8):(3'h6)] <= reg1230[(2'h2):(2'h2)])});
                      reg2723 <= $signed((^~(^~reg1200)));
                    end
                  else
                    begin
                      reg2721 <= (8'ha7);
                      reg2722 <= reg2722;
                      reg2723 <= reg2720[(1'h0):(1'h0)];
                    end
                  if (forvar2753)
                    begin
                      reg2724 <= $signed(reg1217[(3'h5):(1'h1)]);
                    end
                  else
                    begin
                      reg2724 <= ($unsigned({(reg2716 ^ forvar2754)}) ?
                          (~(forvar2712[(1'h0):(1'h0)] ?
                              (~(8'haa)) : (reg2769 ?
                                  (8'hb7) : forvar2741))) : (reg2754 ?
                              $unsigned(reg2761[(3'h6):(3'h5)]) : reg1220[(4'ha):(4'ha)]));
                      reg2725 <= $unsigned((8'hb7));
                    end
                  reg2726 <= {(({reg1234} >> (^reg2759)) ?
                          {reg2752} : {(^~reg1237)})};
                end
              else
                begin
                  if ((~reg2712[(1'h1):(1'h0)]))
                    begin
                      reg2720 <= (^~$unsigned((forvar2710 >= (~^reg2768))));
                      reg2721 <= reg1220;
                      reg2722 <= reg2748;
                    end
                  else
                    begin
                      reg2720 <= (&((^~forvar2715) ~^ (-reg2759)));
                      reg2721 <= ((!forvar2730) & (8'h9e));
                    end
                  for (forvar2723 = (1'h0); (forvar2723 < (1'h1)); forvar2723 = (forvar2723 + (1'h1)))
                    begin
                      reg2724 <= $signed($unsigned(reg2718[(1'h0):(1'h0)]));
                      reg2725 <= ($unsigned((reg2747[(5'h10):(4'h8)] ?
                              $unsigned(reg2760) : (reg2757 ?
                                  forvar2715 : (8'ha1)))) ?
                          (reg1209 ?
                              $signed(reg2708) : $signed((-forvar2763))) : ({(wire1191 ?
                                      (8'ha1) : forvar2712)} ?
                              ((-reg2719) ?
                                  (|reg1222) : (reg1210 ?
                                      forvar2708 : reg1234)) : reg2716[(2'h3):(2'h3)]));
                      reg2726 <= ($unsigned(forvar2730) > {forvar2736[(1'h1):(1'h1)]});
                      reg2727 <= $signed(forvar2755[(4'ha):(2'h3)]);
                    end
                end
            end
          else
            begin
              reg2710 <= $signed($signed(((reg2760 && reg2771) * reg1202)));
              for (forvar2711 = (1'h0); (forvar2711 < (1'h1)); forvar2711 = (forvar2711 + (1'h1)))
                begin
                  for (forvar2712 = (1'h0); (forvar2712 < (1'h1)); forvar2712 = (forvar2712 + (1'h1)))
                    begin
                      reg2713 <= reg1239[(4'hd):(4'h9)];
                    end
                end
              reg2714 <= (&reg1210[(4'hf):(1'h0)]);
            end
          reg2728 <= ($signed(($unsigned(reg2761) | (reg1234 ?
                  (8'hac) : reg2762))) ?
              forvar2754 : reg2761[(1'h0):(1'h0)]);
        end
      for (forvar2773 = (1'h0); (forvar2773 < (2'h2)); forvar2773 = (forvar2773 + (1'h1)))
        begin
          for (forvar2774 = (1'h0); (forvar2774 < (2'h2)); forvar2774 = (forvar2774 + (1'h1)))
            begin
              if (reg2721)
                begin
                  reg2775 <= reg2709[(2'h3):(1'h0)];
                end
              else
                begin
                  reg2775 <= $unsigned(reg1216[(3'h6):(3'h6)]);
                  for (forvar2776 = (1'h0); (forvar2776 < (2'h3)); forvar2776 = (forvar2776 + (1'h1)))
                    begin
                      reg2777 <= $unsigned($unsigned($unsigned({(8'hb7)})));
                      reg2778 <= $unsigned((^~reg2724));
                      reg2779 <= (-(((^reg2777) ? {reg2717} : (^reg2737)) ?
                          (8'hb0) : (forvar2708[(1'h1):(1'h0)] ?
                              reg2725[(3'h6):(1'h1)] : (reg2714 > reg2719))));
                      reg2780 <= ((reg2754[(1'h1):(1'h0)] ?
                              reg1224 : wire1190) ?
                          ((wire1192 ?
                              $signed(forvar2711) : reg1198) * (reg2779 <<< reg2744[(3'h7):(2'h2)])) : reg2726);
                    end
                  reg2781 <= $signed((|{(^~reg2746)}));
                  for (forvar2782 = (1'h0); (forvar2782 < (2'h2)); forvar2782 = (forvar2782 + (1'h1)))
                    begin
                      reg2783 <= ((&$unsigned((reg2768 != forvar2723))) > {(&(+(8'hb8)))});
                    end
                end
              if ((-(^~reg2762[(4'h9):(3'h7)])))
                begin
                  for (forvar2784 = (1'h0); (forvar2784 < (2'h2)); forvar2784 = (forvar2784 + (1'h1)))
                    begin
                      reg2785 <= forvar2710[(2'h2):(2'h2)];
                      reg2786 <= $signed($signed($unsigned({forvar2723})));
                      reg2787 <= (~$unsigned(reg2779));
                    end
                  reg2788 <= $unsigned(forvar2767[(4'he):(3'h7)]);
                  for (forvar2789 = (1'h0); (forvar2789 < (1'h1)); forvar2789 = (forvar2789 + (1'h1)))
                    begin
                      reg2790 <= forvar2710[(2'h2):(2'h2)];
                      reg2791 <= reg1223[(2'h2):(1'h1)];
                    end
                  for (forvar2792 = (1'h0); (forvar2792 < (2'h3)); forvar2792 = (forvar2792 + (1'h1)))
                    begin
                      reg2793 <= {reg2748[(3'h4):(1'h0)]};
                    end
                end
              else
                begin
                  reg2784 <= reg2732[(1'h1):(1'h0)];
                end
            end
          for (forvar2794 = (1'h0); (forvar2794 < (2'h3)); forvar2794 = (forvar2794 + (1'h1)))
            begin
              reg2795 <= forvar2709[(5'h10):(4'ha)];
              if ($unsigned($unsigned(($signed(reg2779) ?
                  (reg2723 ? reg2766 : reg2738) : $signed(reg2728)))))
                begin
                  if (reg2762[(1'h1):(1'h1)])
                    begin
                      reg2796 <= $unsigned($signed(reg2786[(1'h0):(1'h0)]));
                      reg2797 <= reg2790[(1'h1):(1'h1)];
                      reg2798 <= $unsigned($unsigned(reg2729[(4'h8):(2'h3)]));
                    end
                  else
                    begin
                      reg2796 <= (8'hb7);
                      reg2797 <= (($unsigned(reg2780[(4'h8):(1'h1)]) ?
                              $signed((~^reg2797)) : ($signed(reg2759) ?
                                  $signed((8'hb3)) : reg2764[(3'h5):(3'h5)])) ?
                          $unsigned({(&reg2796)}) : (8'hb8));
                      reg2798 <= forvar2774[(1'h1):(1'h0)];
                      reg2799 <= (|(($signed(reg1224) ?
                          (reg2785 ?
                              wire1191 : (8'hb5)) : $signed(reg1223)) + ($signed(reg2718) ?
                          (reg2729 > (8'hab)) : (~&reg2710))));
                    end
                  if ((|$signed(((~^reg1214) ?
                      (reg2770 + reg2770) : $signed(reg2746)))))
                    begin
                      reg2800 <= forvar2723[(2'h3):(2'h2)];
                      reg2801 <= $signed(reg2748);
                      reg2802 <= ((reg2708[(2'h3):(1'h1)] & reg1209) >> ($signed(reg1213[(4'ha):(4'h9)]) ?
                          $unsigned($signed(reg2754)) : ({reg2791} ?
                              (forvar2710 ?
                                  forvar2784 : reg2787) : $unsigned(forvar2708))));
                      reg2803 <= reg1203;
                    end
                  else
                    begin
                      reg2800 <= reg2735[(1'h0):(1'h0)];
                      reg2801 <= {$signed($unsigned((forvar2774 << (8'hb7))))};
                      reg2802 <= wire1190;
                    end
                  for (forvar2804 = (1'h0); (forvar2804 < (2'h3)); forvar2804 = (forvar2804 + (1'h1)))
                    begin
                      reg2805 <= $signed(reg1199[(3'h4):(2'h3)]);
                      reg2806 <= $signed(reg2755);
                      reg2807 <= (-($signed((|reg1217)) ?
                          ((reg2714 & forvar2774) ?
                              (forvar2755 & reg2752) : reg2748[(4'hc):(2'h2)]) : reg2762[(4'hc):(4'h9)]));
                      reg2808 <= reg2737[(3'h7):(3'h7)];
                    end
                end
              else
                begin
                  for (forvar2796 = (1'h0); (forvar2796 < (1'h0)); forvar2796 = (forvar2796 + (1'h1)))
                    begin
                      reg2797 <= (|((~&(reg2710 ? forvar2725 : reg2786)) ?
                          {$signed(reg2784)} : (~(reg2784 >>> reg2723))));
                    end
                  for (forvar2798 = (1'h0); (forvar2798 < (2'h3)); forvar2798 = (forvar2798 + (1'h1)))
                    begin
                      reg2799 <= (8'hb2);
                    end
                end
            end
          for (forvar2809 = (1'h0); (forvar2809 < (1'h1)); forvar2809 = (forvar2809 + (1'h1)))
            begin
              if (($signed(forvar2730[(3'h7):(2'h3)]) << $signed((-forvar2711))))
                begin
                  if (reg2720)
                    begin
                      reg2810 <= ($unsigned(($unsigned(reg1233) < (forvar2710 * reg2756))) ?
                          ((reg1220[(4'ha):(1'h0)] != (reg1235 ?
                              reg2708 : reg2739)) > reg2748) : $signed($unsigned($signed(reg2729))));
                      reg2811 <= reg2786;
                    end
                  else
                    begin
                      reg2810 <= (-reg1227);
                    end
                  for (forvar2812 = (1'h0); (forvar2812 < (2'h3)); forvar2812 = (forvar2812 + (1'h1)))
                    begin
                      reg2813 <= {$signed($unsigned($signed(reg2786)))};
                      reg2814 <= (8'hb4);
                      reg2815 <= (^(!(-(+forvar2725))));
                    end
                  for (forvar2816 = (1'h0); (forvar2816 < (1'h0)); forvar2816 = (forvar2816 + (1'h1)))
                    begin
                      reg2817 <= ({$signed((!reg2712))} - reg2725[(4'h8):(1'h1)]);
                      reg2818 <= reg2781[(3'h6):(3'h4)];
                    end
                end
              else
                begin
                  for (forvar2810 = (1'h0); (forvar2810 < (1'h1)); forvar2810 = (forvar2810 + (1'h1)))
                    begin
                      reg2811 <= ((8'had) >>> $signed((8'hb1)));
                      reg2812 <= (reg2780 ?
                          ((&$unsigned(reg2815)) ?
                              reg2781 : $signed($signed(reg2710))) : forvar2712[(1'h0):(1'h0)]);
                      reg2813 <= reg2735[(1'h1):(1'h1)];
                      reg2814 <= (~{((!reg2755) ?
                              (reg2725 ^~ reg1238) : reg2717[(3'h7):(1'h0)])});
                    end
                end
            end
          if (wire1193)
            begin
              for (forvar2819 = (1'h0); (forvar2819 < (1'h1)); forvar2819 = (forvar2819 + (1'h1)))
                begin
                  reg2820 <= ($signed(((!reg1224) & reg1208)) << {{forvar2798}});
                  for (forvar2821 = (1'h0); (forvar2821 < (2'h2)); forvar2821 = (forvar2821 + (1'h1)))
                    begin
                      reg2822 <= $unsigned({({(8'ha7)} ?
                              (reg2757 ?
                                  reg2800 : reg2807) : $signed((8'ha8)))});
                      reg2823 <= {$unsigned(forvar2716[(3'h7):(1'h1)])};
                      reg2824 <= (&$unsigned((reg2772[(2'h2):(2'h2)] | ((8'hb3) ?
                          reg2749 : wire1188))));
                    end
                  for (forvar2825 = (1'h0); (forvar2825 < (1'h0)); forvar2825 = (forvar2825 + (1'h1)))
                    begin
                      reg2826 <= (((reg1224 ? {reg1230} : reg2787) ?
                          $unsigned(forvar2754) : forvar2755[(1'h0):(1'h0)]) >>> (-$signed((reg2802 << reg2746))));
                      reg2827 <= reg1203[(4'hd):(1'h1)];
                      reg2828 <= reg2769[(2'h3):(1'h1)];
                    end
                end
            end
          else
            begin
              reg2819 <= $unsigned(forvar2794[(4'h9):(2'h3)]);
              if ($unsigned(($signed(reg1235[(1'h1):(1'h1)]) <<< reg2811[(1'h1):(1'h1)])))
                begin
                  if ($unsigned((-reg2714[(4'ha):(4'h9)])))
                    begin
                      reg2820 <= (({(8'hb6)} >> reg2768) ?
                          {$unsigned((reg2758 ?
                                  forvar2809 : reg2762))} : forvar2754[(4'hb):(3'h5)]);
                      reg2821 <= {((8'hb6) ?
                              reg2779 : $signed(forvar2715[(2'h3):(1'h1)]))};
                    end
                  else
                    begin
                      reg2820 <= ((-(~|(reg2788 ? reg2798 : reg1234))) ?
                          {$signed(forvar2776)} : reg2740);
                      reg2821 <= $signed($signed(reg2744[(1'h0):(1'h0)]));
                      reg2822 <= $signed((((reg2784 ?
                          (8'ha4) : reg2808) > reg2735) * $signed(forvar2825[(1'h0):(1'h0)])));
                    end
                  if ($signed(wire1191))
                    begin
                      reg2823 <= reg2735[(2'h2):(2'h2)];
                      reg2824 <= (((reg2766 ?
                          forvar2709[(5'h10):(5'h10)] : (forvar2792 >= forvar2730)) + $unsigned($signed(reg1232))) ~^ $unsigned(((&reg2722) ?
                          $signed((8'hae)) : reg2795[(3'h7):(2'h2)])));
                    end
                  else
                    begin
                      reg2823 <= $unsigned({$unsigned(forvar2782)});
                      reg2824 <= ($unsigned(((reg2756 ? reg1223 : forvar2755) ?
                          forvar2809 : $signed(reg2720))) | reg2815);
                      reg2825 <= (^(&((reg1230 * reg2752) ^ (reg2742 ?
                          wire1189 : reg2797))));
                      reg2826 <= (((reg2827[(2'h2):(2'h2)] ?
                          {reg2803} : (~forvar2792)) - $signed(reg2718)) <<< ($unsigned((reg2790 ?
                              reg1219 : forvar2792)) ?
                          reg2708 : (reg2802 ?
                              $unsigned(reg2751) : reg1228[(1'h0):(1'h0)])));
                    end
                  if (reg1217[(3'h4):(2'h2)])
                    begin
                      reg2827 <= (^~reg2754);
                      reg2828 <= (8'ha9);
                    end
                  else
                    begin
                      reg2827 <= ($unsigned(reg2813[(2'h3):(2'h2)]) + $unsigned(reg1205[(3'h4):(2'h3)]));
                      reg2828 <= reg2783;
                      reg2829 <= forvar2773[(2'h2):(1'h0)];
                    end
                  if (((reg2796 <= ($unsigned(forvar2758) ?
                      reg1230 : (+reg2779))) | $unsigned(forvar2809[(1'h0):(1'h0)])))
                    begin
                      reg2830 <= (~|$unsigned(reg2819[(3'h5):(2'h2)]));
                      reg2831 <= reg2754;
                    end
                  else
                    begin
                      reg2830 <= (|$unsigned((&(reg1216 ? reg2742 : reg2714))));
                    end
                end
              else
                begin
                  for (forvar2820 = (1'h0); (forvar2820 < (1'h0)); forvar2820 = (forvar2820 + (1'h1)))
                    begin
                      reg2821 <= ($signed(reg2712) & {(((8'ha6) && reg2720) ?
                              reg2826 : (~&reg1215))});
                      reg2822 <= (-$unsigned(($signed(reg2756) || {reg2725})));
                    end
                  if ($unsigned($unsigned($signed(forvar2710))))
                    begin
                      reg2823 <= ((8'h9f) ?
                          {($signed(forvar2715) ?
                                  (|reg2811) : (reg1230 ?
                                      reg2752 : reg1239))} : $unsigned(reg2720));
                      reg2824 <= $signed({forvar2825[(2'h3):(1'h1)]});
                      reg2825 <= (~&(-$unsigned($unsigned(reg1205))));
                    end
                  else
                    begin
                      reg2823 <= forvar2715;
                      reg2824 <= (($signed((+reg1205)) == $unsigned((reg2748 ?
                              reg2824 : reg2759))) ?
                          reg2786 : {(!(^~reg2717))});
                      reg2825 <= (~&(reg2769 ?
                          wire1192 : reg2808[(4'hf):(1'h0)]));
                      reg2826 <= ($unsigned(reg2739[(2'h3):(1'h0)]) ?
                          $unsigned((^~$signed(reg2766))) : $unsigned((~^(~|reg2793))));
                    end
                  reg2827 <= reg2807;
                end
              for (forvar2832 = (1'h0); (forvar2832 < (2'h3)); forvar2832 = (forvar2832 + (1'h1)))
                begin
                  if ((~^($signed((~reg1197)) ~^ ((reg1232 <<< reg2762) ?
                      reg2728 : $signed((8'ha9))))))
                    begin
                      reg2833 <= reg2723;
                      reg2834 <= (~forvar2809);
                      reg2835 <= ((^forvar2745[(3'h7):(1'h0)]) ?
                          $signed(($signed(reg1229) >>> $unsigned(reg2724))) : $unsigned(reg2834[(3'h4):(2'h3)]));
                      reg2836 <= wire1187;
                    end
                  else
                    begin
                      reg2833 <= (^~$signed($unsigned($unsigned(reg1215))));
                      reg2834 <= {(&($signed(wire1191) >> (forvar2796 ?
                              reg1208 : reg2710)))};
                      reg2835 <= reg1233[(2'h2):(1'h1)];
                    end
                end
            end
        end
    end
  assign wire2837 = reg1208[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      if (reg2760[(1'h0):(1'h0)])
        begin
          reg2838 <= (-(|$signed(reg2724)));
          if (reg2720[(1'h0):(1'h0)])
            begin
              for (forvar2839 = (1'h0); (forvar2839 < (1'h1)); forvar2839 = (forvar2839 + (1'h1)))
                begin
                  for (forvar2840 = (1'h0); (forvar2840 < (1'h1)); forvar2840 = (forvar2840 + (1'h1)))
                    begin
                      reg2841 <= $unsigned((((8'h9d) && $signed(reg2810)) ?
                          ((reg2757 ? reg2779 : reg2768) ~^ (reg2834 ?
                              reg1224 : reg2805)) : reg2716[(2'h2):(1'h1)]));
                      reg2842 <= wire1189[(1'h1):(1'h0)];
                      reg2843 <= reg1223[(2'h2):(1'h1)];
                    end
                end
            end
          else
            begin
              for (forvar2839 = (1'h0); (forvar2839 < (2'h2)); forvar2839 = (forvar2839 + (1'h1)))
                begin
                  for (forvar2840 = (1'h0); (forvar2840 < (1'h0)); forvar2840 = (forvar2840 + (1'h1)))
                    begin
                      reg2841 <= {(reg2760[(4'h8):(2'h3)] ?
                              reg2828[(4'hc):(3'h6)] : {((8'h9e) ?
                                      reg2770 : reg2727)})};
                    end
                  reg2842 <= wire1241[(1'h0):(1'h0)];
                  if (($unsigned(forvar2839) ?
                      ({(reg2750 ? reg2756 : wire1190)} ?
                          $unsigned((reg2841 ?
                              reg2797 : reg1215)) : reg2793[(1'h1):(1'h0)]) : $unsigned((~|{reg1226}))))
                    begin
                      reg2843 <= reg1220;
                    end
                  else
                    begin
                      reg2843 <= $signed(reg1223[(2'h3):(1'h1)]);
                      reg2844 <= (|$signed($signed($signed(reg2781))));
                    end
                end
              for (forvar2845 = (1'h0); (forvar2845 < (2'h2)); forvar2845 = (forvar2845 + (1'h1)))
                begin
                  for (forvar2846 = (1'h0); (forvar2846 < (2'h3)); forvar2846 = (forvar2846 + (1'h1)))
                    begin
                      reg2847 <= $unsigned(((reg2727[(3'h4):(2'h3)] ?
                          $signed(reg2748) : (^(8'ha4))) >= ((reg2822 + reg2793) || reg2752)));
                    end
                  if (reg2797)
                    begin
                      reg2848 <= ($unsigned(((reg2727 <= (8'hb7)) || reg2815)) ?
                          {$signed({reg2779})} : $unsigned(reg2818[(3'h5):(1'h1)]));
                      reg2849 <= reg2844;
                      reg2850 <= reg1200[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg2848 <= reg2735;
                      reg2849 <= reg2834;
                    end
                end
              for (forvar2851 = (1'h0); (forvar2851 < (1'h0)); forvar2851 = (forvar2851 + (1'h1)))
                begin
                  for (forvar2852 = (1'h0); (forvar2852 < (1'h1)); forvar2852 = (forvar2852 + (1'h1)))
                    begin
                      reg2853 <= $unsigned($signed($signed({reg2833})));
                      reg2854 <= (((8'ha3) ?
                          $unsigned((reg1217 ?
                              reg2853 : reg2783)) : (((8'ha7) - (8'ha0)) >>> ((8'hb8) - reg2830))) <<< ($unsigned((reg2735 < wire1188)) ^~ {{reg2800}}));
                    end
                  for (forvar2855 = (1'h0); (forvar2855 < (1'h1)); forvar2855 = (forvar2855 + (1'h1)))
                    begin
                      reg2856 <= reg2770;
                    end
                  if (({reg2731} ?
                      reg2849 : (forvar2852 ?
                          reg2783[(3'h7):(2'h2)] : $signed({reg2788}))))
                    begin
                      reg2857 <= {(-{reg2812[(2'h3):(2'h3)]})};
                    end
                  else
                    begin
                      reg2857 <= $unsigned($unsigned(reg2718));
                      reg2858 <= reg2812;
                    end
                end
            end
          for (forvar2859 = (1'h0); (forvar2859 < (1'h0)); forvar2859 = (forvar2859 + (1'h1)))
            begin
              for (forvar2860 = (1'h0); (forvar2860 < (1'h1)); forvar2860 = (forvar2860 + (1'h1)))
                begin
                  for (forvar2861 = (1'h0); (forvar2861 < (1'h1)); forvar2861 = (forvar2861 + (1'h1)))
                    begin
                      reg2862 <= (reg2785 >>> $signed($unsigned((reg2831 ?
                          (8'ha0) : reg2770))));
                      reg2863 <= reg1216;
                    end
                  for (forvar2864 = (1'h0); (forvar2864 < (2'h3)); forvar2864 = (forvar2864 + (1'h1)))
                    begin
                      reg2865 <= $unsigned($unsigned(reg1233[(1'h0):(1'h0)]));
                    end
                  if (((!(~$signed(reg1214))) == ({reg2709[(1'h1):(1'h0)]} != $unsigned(reg1213[(2'h3):(2'h3)]))))
                    begin
                      reg2866 <= ($signed((-(~^reg2856))) | {(((8'h9e) ^ reg1214) ?
                              (reg2778 ? reg2720 : reg2834) : {reg2823})});
                      reg2867 <= ((((reg2802 | reg2788) && reg2716[(2'h3):(2'h2)]) ?
                              $signed($unsigned(reg2827)) : reg2770) ?
                          ((reg1223[(2'h3):(2'h2)] && (reg2733 ?
                                  reg2810 : reg2850)) ?
                              reg1214[(4'h8):(2'h2)] : reg2847[(2'h2):(2'h2)]) : reg2850[(4'h9):(3'h7)]);
                      reg2868 <= (reg2769[(3'h6):(3'h6)] <= {reg2772[(2'h2):(1'h1)]});
                      reg2869 <= $signed($signed(reg2752));
                    end
                  else
                    begin
                      reg2866 <= (~^{reg2869});
                      reg2867 <= (!((-$signed(wire1189)) >= ($unsigned(reg2743) ?
                          $unsigned(forvar2860) : (reg2847 | reg2766))));
                      reg2868 <= (((8'had) ?
                          {reg2821} : ($signed(reg2833) ?
                              (^reg1197) : reg1210[(4'he):(2'h2)])) - ($signed({reg2731}) == {(&reg2764)}));
                    end
                end
              reg2870 <= $unsigned(($signed(reg2829[(1'h0):(1'h0)]) ?
                  {$signed(reg2833)} : {((8'hb8) ? reg2771 : reg2825)}));
            end
          reg2871 <= ($unsigned(reg2812[(4'h8):(2'h3)]) ?
              $signed(reg2711) : $signed(reg1235[(2'h3):(2'h2)]));
        end
      else
        begin
          for (forvar2838 = (1'h0); (forvar2838 < (1'h1)); forvar2838 = (forvar2838 + (1'h1)))
            begin
              if (reg2740)
                begin
                  if (reg2709[(3'h7):(3'h7)])
                    begin
                      reg2839 <= $signed(reg2742);
                      reg2840 <= ($unsigned(((!reg2828) ?
                          {reg1219} : reg2798[(1'h0):(1'h0)])) <= (8'ha5));
                      reg2841 <= (($signed(reg2716[(1'h1):(1'h1)]) ^ {(reg2796 <= (8'hb2))}) ?
                          (^(8'ha1)) : $signed((8'hb6)));
                    end
                  else
                    begin
                      reg2839 <= ({$unsigned({reg2759})} ?
                          reg2735[(2'h3):(2'h3)] : {$signed((reg2797 >= reg2769))});
                    end
                  reg2842 <= $unsigned($signed($unsigned($unsigned(reg1223))));
                  for (forvar2843 = (1'h0); (forvar2843 < (1'h0)); forvar2843 = (forvar2843 + (1'h1)))
                    begin
                      reg2844 <= reg2856[(3'h6):(2'h3)];
                      reg2845 <= {($unsigned(((8'hb1) | reg2765)) ?
                              $signed((&reg2715)) : $signed(reg1230))};
                      reg2846 <= $unsigned(wire1188[(3'h4):(2'h3)]);
                      reg2847 <= $unsigned({($signed(reg1214) + {reg2768})});
                    end
                  reg2848 <= $signed($signed(reg2717[(2'h2):(1'h1)]));
                end
              else
                begin
                  if (reg2835[(1'h0):(1'h0)])
                    begin
                      reg2839 <= reg1214[(2'h3):(1'h1)];
                      reg2840 <= reg2805;
                      reg2841 <= reg2713[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg2839 <= $signed($signed(reg2786));
                    end
                  if ($signed($signed({(^~forvar2840)})))
                    begin
                      reg2842 <= ($signed($signed((reg2783 ^ wire2706))) ?
                          (8'h9c) : wire1191);
                      reg2843 <= ((~^$unsigned($unsigned(reg2833))) & (reg2803[(2'h3):(2'h2)] >> $signed((reg2863 ?
                          reg2720 : reg2713))));
                    end
                  else
                    begin
                      reg2842 <= $unsigned((reg2829 * reg1222[(4'h8):(1'h1)]));
                      reg2843 <= $unsigned(((~&reg1224) ?
                          reg2805[(3'h7):(3'h5)] : $unsigned((~&reg2850))));
                      reg2844 <= ((~|$unsigned((!forvar2860))) || (8'hae));
                      reg2845 <= ((~|reg2759) - $unsigned(reg2790[(3'h6):(1'h1)]));
                    end
                end
              reg2849 <= (|$signed({(&reg2834)}));
              for (forvar2850 = (1'h0); (forvar2850 < (1'h1)); forvar2850 = (forvar2850 + (1'h1)))
                begin
                  if (reg2830)
                    begin
                      reg2851 <= reg2821;
                    end
                  else
                    begin
                      reg2851 <= reg1240;
                    end
                  reg2852 <= wire1241[(2'h3):(2'h2)];
                  for (forvar2853 = (1'h0); (forvar2853 < (2'h3)); forvar2853 = (forvar2853 + (1'h1)))
                    begin
                      reg2854 <= ({((reg2830 && reg2718) == $unsigned(reg1222))} != reg2775[(3'h4):(2'h2)]);
                      reg2855 <= ($signed((((8'hab) ?
                              (8'hb5) : reg2778) == (wire2837 ?
                              reg2830 : reg2763))) ?
                          (~|((~wire1188) ~^ reg1220)) : (^reg2849));
                      reg2856 <= {$unsigned((&$unsigned(reg2853)))};
                    end
                  for (forvar2857 = (1'h0); (forvar2857 < (1'h0)); forvar2857 = (forvar2857 + (1'h1)))
                    begin
                      reg2858 <= $unsigned((+$unsigned((reg2870 * (8'hac)))));
                      reg2859 <= (|(~|$unsigned($unsigned(reg1224))));
                      reg2860 <= reg2777;
                      reg2861 <= reg2831[(3'h4):(1'h0)];
                    end
                end
              for (forvar2862 = (1'h0); (forvar2862 < (1'h0)); forvar2862 = (forvar2862 + (1'h1)))
                begin
                  if (forvar2845[(4'hc):(1'h1)])
                    begin
                      reg2863 <= ($unsigned(((reg2835 >= reg2863) ?
                          (~^reg2871) : (reg2862 != reg2844))) >= reg2770[(3'h6):(1'h1)]);
                    end
                  else
                    begin
                      reg2863 <= {reg1219[(1'h1):(1'h0)]};
                      reg2864 <= reg2728;
                      reg2865 <= {reg2775[(3'h4):(2'h3)]};
                    end
                end
            end
        end
      for (forvar2872 = (1'h0); (forvar2872 < (2'h3)); forvar2872 = (forvar2872 + (1'h1)))
        begin
          reg2873 <= (~&({((8'had) << reg2807)} * reg2865[(1'h0):(1'h0)]));
          for (forvar2874 = (1'h0); (forvar2874 < (1'h0)); forvar2874 = (forvar2874 + (1'h1)))
            begin
              for (forvar2875 = (1'h0); (forvar2875 < (2'h3)); forvar2875 = (forvar2875 + (1'h1)))
                begin
                  for (forvar2876 = (1'h0); (forvar2876 < (2'h3)); forvar2876 = (forvar2876 + (1'h1)))
                    begin
                      reg2877 <= reg2802[(2'h3):(1'h1)];
                      reg2878 <= ($signed(($unsigned(reg1199) ?
                              $unsigned(reg2715) : (!reg2856))) ?
                          reg2734 : {reg2836[(2'h3):(2'h3)]});
                      reg2879 <= $unsigned((^reg2771[(4'hd):(4'hd)]));
                    end
                  reg2880 <= forvar2876;
                end
              for (forvar2881 = (1'h0); (forvar2881 < (1'h1)); forvar2881 = (forvar2881 + (1'h1)))
                begin
                  reg2882 <= $unsigned((~((~&(8'hb4)) == $unsigned(forvar2851))));
                  if ((~^(&reg2858)))
                    begin
                      reg2883 <= (reg2849[(2'h2):(2'h2)] || ((^~(&(8'had))) ?
                          $signed({(8'ha0)}) : reg2826));
                      reg2884 <= $unsigned(($signed(((8'hb8) ?
                              reg2825 : forvar2838)) ?
                          ((reg2755 & reg2765) ?
                              reg2828[(2'h2):(2'h2)] : reg2742[(2'h3):(1'h1)]) : reg2869[(1'h0):(1'h0)]));
                      reg2885 <= (&(&(reg2788 ?
                          (reg2823 ? forvar2859 : reg1238) : reg2847)));
                      reg2886 <= (({reg1210} < forvar2875) ?
                          $signed(((^~(8'ha5)) & (reg2806 - reg2807))) : reg1219);
                    end
                  else
                    begin
                      reg2883 <= {(^$unsigned(((8'ha5) ? reg2883 : reg1216)))};
                      reg2884 <= reg2738[(1'h1):(1'h1)];
                      reg2885 <= (^~reg2856);
                      reg2886 <= ({(+reg2790[(3'h5):(3'h5)])} ?
                          reg1228[(1'h1):(1'h0)] : $unsigned($unsigned((~|reg1228))));
                    end
                  for (forvar2887 = (1'h0); (forvar2887 < (1'h1)); forvar2887 = (forvar2887 + (1'h1)))
                    begin
                      reg2888 <= (^~(reg2772 ?
                          reg2849[(1'h0):(1'h0)] : $unsigned($signed((8'ha0)))));
                    end
                end
              reg2889 <= reg2846;
            end
          if ({reg2836[(3'h5):(3'h4)]})
            begin
              for (forvar2890 = (1'h0); (forvar2890 < (2'h3)); forvar2890 = (forvar2890 + (1'h1)))
                begin
                  if (reg2752)
                    begin
                      reg2891 <= reg2807[(1'h1):(1'h1)];
                      reg2892 <= (~&reg2858);
                    end
                  else
                    begin
                      reg2891 <= reg2891;
                      reg2892 <= reg1199;
                    end
                end
            end
          else
            begin
              for (forvar2890 = (1'h0); (forvar2890 < (2'h3)); forvar2890 = (forvar2890 + (1'h1)))
                begin
                  for (forvar2891 = (1'h0); (forvar2891 < (2'h3)); forvar2891 = (forvar2891 + (1'h1)))
                    begin
                      reg2892 <= (wire1188 || $unsigned((8'ha3)));
                    end
                  if ({({forvar2864} ~^ $unsigned(reg2748))})
                    begin
                      reg2893 <= reg2771;
                      reg2894 <= reg2775;
                    end
                  else
                    begin
                      reg2893 <= {(^~((~^forvar2887) >>> (reg2824 ?
                              reg1238 : reg2761)))};
                      reg2894 <= reg2886[(3'h7):(2'h2)];
                      reg2895 <= reg2791;
                      reg2896 <= (|(^{{reg2857}}));
                    end
                end
              reg2897 <= ((8'h9e) & (reg1223[(2'h2):(2'h2)] != $unsigned(((8'h9d) << reg2813))));
            end
        end
      if ((~|reg2712))
        begin
          if ((reg2787[(4'h8):(2'h3)] ?
              reg2778[(2'h2):(1'h0)] : ({reg2747[(5'h10):(3'h7)]} ?
                  {forvar2875} : reg2812[(4'hb):(2'h2)])))
            begin
              for (forvar2898 = (1'h0); (forvar2898 < (1'h0)); forvar2898 = (forvar2898 + (1'h1)))
                begin
                  if ({((^~(reg2867 << reg2746)) ^~ {(^wire1188)})})
                    begin
                      reg2899 <= $unsigned($unsigned(reg2737));
                      reg2900 <= (reg2896 ?
                          ((reg1234 >> reg2756[(4'ha):(1'h1)]) ?
                              reg2854 : (reg2833[(4'hb):(1'h1)] << $signed(reg2870))) : reg2756);
                      reg2901 <= (8'ha4);
                    end
                  else
                    begin
                      reg2899 <= ($unsigned({{forvar2864}}) ?
                          (reg2844[(3'h5):(3'h5)] != $unsigned((reg2895 >>> reg2883))) : (forvar2861 ~^ {(!reg2883)}));
                      reg2900 <= reg2725;
                    end
                  reg2902 <= (~$signed($unsigned($unsigned(reg2883))));
                end
              for (forvar2903 = (1'h0); (forvar2903 < (1'h1)); forvar2903 = (forvar2903 + (1'h1)))
                begin
                  for (forvar2904 = (1'h0); (forvar2904 < (2'h2)); forvar2904 = (forvar2904 + (1'h1)))
                    begin
                      reg2905 <= reg2724;
                    end
                end
              for (forvar2906 = (1'h0); (forvar2906 < (2'h3)); forvar2906 = (forvar2906 + (1'h1)))
                begin
                  if (reg2712)
                    begin
                      reg2907 <= reg2720;
                    end
                  else
                    begin
                      reg2907 <= (forvar2898 ?
                          (!(reg2757[(4'h8):(1'h0)] ?
                              (reg2743 ?
                                  reg2715 : reg2770) : $signed(reg2762))) : reg2877);
                      reg2908 <= ({reg2829} ?
                          forvar2890[(2'h3):(1'h0)] : (8'h9c));
                      reg2909 <= reg1208[(4'he):(3'h6)];
                      reg2910 <= reg2779[(4'hf):(2'h3)];
                    end
                  if ((~^$signed($signed((reg1216 ? (8'had) : reg2856)))))
                    begin
                      reg2911 <= ((reg2793[(1'h0):(1'h0)] ?
                          forvar2862[(2'h2):(2'h2)] : $unsigned($unsigned(reg2814))) << $signed(($signed((8'hb1)) <<< $signed(reg2735))));
                      reg2912 <= $unsigned(reg2822);
                    end
                  else
                    begin
                      reg2911 <= reg1202[(3'h7):(2'h2)];
                      reg2912 <= $unsigned({((reg2737 == reg2752) ?
                              reg2836[(2'h2):(1'h1)] : $unsigned(forvar2857))});
                    end
                  if (reg2714)
                    begin
                      reg2913 <= $signed($unsigned({$signed(reg2820)}));
                    end
                  else
                    begin
                      reg2913 <= {{(reg2892[(3'h4):(2'h2)] > {reg2907})}};
                      reg2914 <= (($unsigned($unsigned(reg1228)) ?
                              ($unsigned((8'hae)) | $signed(forvar2853)) : $signed((8'ha2))) ?
                          (8'ha2) : {((forvar2857 < reg1210) ?
                                  $signed((8'hb5)) : reg1223)});
                    end
                end
            end
          else
            begin
              for (forvar2898 = (1'h0); (forvar2898 < (2'h3)); forvar2898 = (forvar2898 + (1'h1)))
                begin
                  for (forvar2899 = (1'h0); (forvar2899 < (2'h3)); forvar2899 = (forvar2899 + (1'h1)))
                    begin
                      reg2900 <= reg2788;
                      reg2901 <= $signed($unsigned($signed((^~reg2799))));
                      reg2902 <= (reg1239[(4'h9):(1'h1)] ?
                          reg2790[(3'h4):(2'h3)] : $signed(reg2787[(2'h3):(2'h3)]));
                      reg2903 <= (|reg2709);
                    end
                  if (reg2871)
                    begin
                      reg2904 <= ((({reg2813} ?
                              forvar2875[(1'h0):(1'h0)] : (-(8'haf))) >> $unsigned((&forvar2891))) ?
                          ($signed($unsigned((8'ha0))) <<< $signed($signed(reg2857))) : $unsigned(reg2739[(3'h4):(2'h3)]));
                    end
                  else
                    begin
                      reg2904 <= (^(~^reg2857[(4'h9):(3'h5)]));
                      reg2905 <= forvar2904[(4'hb):(4'hb)];
                      reg2906 <= reg2732;
                      reg2907 <= $unsigned($signed((reg1198[(3'h4):(3'h4)] == $signed(reg2786))));
                    end
                  for (forvar2908 = (1'h0); (forvar2908 < (1'h1)); forvar2908 = (forvar2908 + (1'h1)))
                    begin
                      reg2909 <= reg2788;
                      reg2910 <= $unsigned(reg2751);
                      reg2911 <= (~reg2732[(1'h0):(1'h0)]);
                    end
                  for (forvar2912 = (1'h0); (forvar2912 < (1'h1)); forvar2912 = (forvar2912 + (1'h1)))
                    begin
                      reg2913 <= (reg2723 ?
                          (reg2719 ?
                              reg2831 : $unsigned((8'hae))) : forvar2860[(4'ha):(4'ha)]);
                      reg2914 <= $unsigned(((-(reg2902 || wire1191)) ?
                          $signed($signed((8'ha1))) : (reg2882[(1'h1):(1'h0)] ^ {reg2784})));
                      reg2915 <= $signed((-$signed($unsigned(reg2877))));
                      reg2916 <= (&(~(reg2729[(2'h3):(1'h0)] >>> {wire1187})));
                    end
                end
            end
          if (reg1213[(4'ha):(1'h0)])
            begin
              for (forvar2917 = (1'h0); (forvar2917 < (1'h1)); forvar2917 = (forvar2917 + (1'h1)))
                begin
                  for (forvar2918 = (1'h0); (forvar2918 < (1'h0)); forvar2918 = (forvar2918 + (1'h1)))
                    begin
                      reg2919 <= reg2756[(4'h9):(3'h5)];
                      reg2920 <= $unsigned(reg2754);
                      reg2921 <= reg2757[(3'h6):(3'h6)];
                    end
                  if ((($unsigned(reg2838) > reg2813[(1'h1):(1'h0)]) != $unsigned((reg2740[(2'h3):(1'h0)] ?
                      $unsigned(reg2760) : $unsigned(wire1191)))))
                    begin
                      reg2922 <= ($signed(wire1188[(3'h6):(3'h4)]) ?
                          $signed(reg2799[(1'h1):(1'h1)]) : $signed($unsigned((reg2709 >> reg1205))));
                    end
                  else
                    begin
                      reg2922 <= reg2834;
                      reg2923 <= {($unsigned(forvar2852[(3'h5):(1'h0)]) >= (-(forvar2906 <= forvar2874)))};
                      reg2924 <= {reg2723[(3'h7):(3'h5)]};
                      reg2925 <= $unsigned($signed({((8'hac) ?
                              forvar2862 : (8'ha6))}));
                    end
                  if ($signed($signed($signed($signed(reg2871)))))
                    begin
                      reg2926 <= (+(^~(((8'hb8) ?
                          reg2758 : reg2743) > (reg2739 ? reg2841 : reg2790))));
                    end
                  else
                    begin
                      reg2926 <= reg2889[(4'ha):(4'h9)];
                      reg2927 <= (($signed(reg1238) ?
                          $unsigned(reg2793[(1'h1):(1'h1)]) : (|$unsigned(reg2815))) & reg2760[(3'h5):(2'h3)]);
                      reg2928 <= $signed($unsigned($unsigned($unsigned(reg2711))));
                    end
                  reg2929 <= $unsigned(((reg2791 <<< $signed(reg2788)) ?
                      (forvar2881[(1'h1):(1'h1)] * ((8'hb3) ?
                          forvar2890 : (8'h9e))) : $signed(reg2896[(3'h4):(3'h4)])));
                end
            end
          else
            begin
              for (forvar2917 = (1'h0); (forvar2917 < (1'h1)); forvar2917 = (forvar2917 + (1'h1)))
                begin
                  reg2918 <= (reg2760 ?
                      ((reg2929[(3'h4):(1'h0)] > $signed(reg2805)) ^ (|$unsigned(reg2766))) : ($signed((reg2788 ^ reg2895)) <<< (&(reg2843 ?
                          reg2819 : reg1210))));
                  reg2919 <= $signed($signed((+((8'ha1) >= reg2902))));
                  for (forvar2920 = (1'h0); (forvar2920 < (2'h3)); forvar2920 = (forvar2920 + (1'h1)))
                    begin
                      reg2921 <= {(8'had)};
                      reg2922 <= (forvar2920[(1'h1):(1'h0)] || ($unsigned((reg2732 & (8'hb2))) ?
                          reg2928 : (|reg2768)));
                      reg2923 <= $unsigned(reg2833[(4'h9):(4'h9)]);
                      reg2924 <= (~|$unsigned(($signed(reg1214) | (reg2713 ?
                          reg2734 : reg2746))));
                    end
                  reg2925 <= $unsigned(reg2848);
                end
              for (forvar2926 = (1'h0); (forvar2926 < (1'h1)); forvar2926 = (forvar2926 + (1'h1)))
                begin
                  for (forvar2927 = (1'h0); (forvar2927 < (2'h2)); forvar2927 = (forvar2927 + (1'h1)))
                    begin
                      reg2928 <= {reg2721};
                    end
                end
            end
          if ((8'hb1))
            begin
              for (forvar2930 = (1'h0); (forvar2930 < (1'h0)); forvar2930 = (forvar2930 + (1'h1)))
                begin
                  reg2931 <= (~^forvar2839);
                end
              for (forvar2932 = (1'h0); (forvar2932 < (2'h2)); forvar2932 = (forvar2932 + (1'h1)))
                begin
                  for (forvar2933 = (1'h0); (forvar2933 < (2'h2)); forvar2933 = (forvar2933 + (1'h1)))
                    begin
                      reg2934 <= (forvar2872[(4'ha):(4'h8)] ?
                          forvar2918[(1'h1):(1'h1)] : {$signed((!reg2731))});
                      reg2935 <= (($signed(reg2732) ^ $unsigned((reg2721 ?
                          forvar2852 : reg2807))) <<< $signed((~$signed(forvar2872))));
                      reg2936 <= forvar2933;
                      reg2937 <= (($signed((reg2797 != forvar2920)) ?
                          reg2802 : $unsigned($unsigned(reg2923))) <= ((^~(reg2860 <<< reg2765)) ?
                          (!(reg2873 ? reg2805 : forvar2930)) : (8'haf)));
                    end
                  reg2938 <= $unsigned(($unsigned((8'ha2)) ?
                      reg2852 : $signed($unsigned(reg2867))));
                  reg2939 <= (forvar2843[(3'h7):(2'h3)] ?
                      reg2708[(1'h0):(1'h0)] : (^(^(-reg2859))));
                  reg2940 <= {(~^$signed(reg2909))};
                end
              if (forvar2851[(2'h2):(2'h2)])
                begin
                  for (forvar2941 = (1'h0); (forvar2941 < (2'h3)); forvar2941 = (forvar2941 + (1'h1)))
                    begin
                      reg2942 <= reg2848;
                      reg2943 <= ({$unsigned((!(8'ha2)))} ^~ (reg2895 + $signed((^~(8'hb5)))));
                    end
                end
              else
                begin
                  for (forvar2941 = (1'h0); (forvar2941 < (1'h1)); forvar2941 = (forvar2941 + (1'h1)))
                    begin
                      reg2942 <= {reg2812[(4'hb):(4'ha)]};
                      reg2943 <= reg1238;
                    end
                  for (forvar2944 = (1'h0); (forvar2944 < (1'h0)); forvar2944 = (forvar2944 + (1'h1)))
                    begin
                      reg2945 <= ((|{(^reg1224)}) + ((~^reg2851) >= (+(~&reg2770))));
                      reg2946 <= forvar2840[(3'h6):(1'h1)];
                      reg2947 <= $unsigned((!((reg2824 << reg2927) ?
                          reg2729[(1'h0):(1'h0)] : (reg2858 * reg2894))));
                    end
                end
              for (forvar2948 = (1'h0); (forvar2948 < (2'h2)); forvar2948 = (forvar2948 + (1'h1)))
                begin
                  if (reg2906[(2'h3):(1'h0)])
                    begin
                      reg2949 <= forvar2941;
                      reg2950 <= (8'h9f);
                      reg2951 <= ((8'h9e) >= reg2910[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg2949 <= ($signed(reg2759[(4'h8):(3'h4)]) << $signed((~(&reg1239))));
                      reg2950 <= $signed($unsigned(reg2818[(2'h3):(2'h2)]));
                      reg2951 <= ((+reg2758[(3'h4):(1'h0)]) ?
                          reg2836[(3'h5):(2'h3)] : $unsigned(($signed(reg2785) && $signed(reg1229))));
                    end
                  for (forvar2952 = (1'h0); (forvar2952 < (1'h1)); forvar2952 = (forvar2952 + (1'h1)))
                    begin
                      reg2953 <= reg2844[(3'h4):(1'h0)];
                      reg2954 <= ({{$unsigned((8'hb4))}} ?
                          {($unsigned(reg2733) ?
                                  (reg2713 ?
                                      reg2853 : reg2861) : reg2901[(2'h2):(1'h1)])} : reg2867);
                      reg2955 <= $signed(reg2909[(2'h2):(1'h0)]);
                      reg2956 <= reg2879;
                    end
                  if (reg2833)
                    begin
                      reg2957 <= forvar2851;
                      reg2958 <= $signed(reg2722[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2957 <= $signed(reg2957);
                    end
                end
            end
          else
            begin
              reg2930 <= ((8'hba) <<< (8'hb4));
            end
          for (forvar2959 = (1'h0); (forvar2959 < (2'h3)); forvar2959 = (forvar2959 + (1'h1)))
            begin
              reg2960 <= reg2947[(1'h1):(1'h1)];
              reg2961 <= reg2811[(2'h2):(1'h1)];
            end
        end
      else
        begin
          for (forvar2898 = (1'h0); (forvar2898 < (2'h2)); forvar2898 = (forvar2898 + (1'h1)))
            begin
              reg2899 <= {(8'ha6)};
              reg2900 <= $unsigned(((forvar2855 && forvar2839) && (8'hb1)));
              for (forvar2901 = (1'h0); (forvar2901 < (1'h1)); forvar2901 = (forvar2901 + (1'h1)))
                begin
                  for (forvar2902 = (1'h0); (forvar2902 < (2'h2)); forvar2902 = (forvar2902 + (1'h1)))
                    begin
                      reg2903 <= ((reg1216[(2'h3):(1'h1)] ?
                          reg1217 : (reg2842[(2'h2):(1'h1)] >> reg2726[(3'h5):(3'h5)])) < (reg1224[(2'h2):(1'h0)] ?
                          reg2724[(3'h4):(1'h1)] : (|$unsigned(forvar2861))));
                      reg2904 <= reg2830[(1'h0):(1'h0)];
                      reg2905 <= (wire1190[(3'h7):(2'h2)] ?
                          $unsigned(reg2844) : (($unsigned(reg2732) - (reg2841 ?
                                  reg2867 : reg2895)) ?
                              ((8'ha3) <<< reg1198[(1'h1):(1'h1)]) : $unsigned((reg2921 ?
                                  reg2913 : reg2779))));
                      reg2906 <= ((~(8'hb0)) ?
                          (reg2763[(3'h4):(1'h0)] != $signed($unsigned(reg2884))) : (((reg2812 <<< forvar2948) >> forvar2857[(4'ha):(2'h2)]) ?
                              reg1235 : ((forvar2862 ?
                                  reg2818 : reg2795) <= (reg2853 ?
                                  forvar2908 : reg2870))));
                    end
                  if ($signed((&{(~^reg2838)})))
                    begin
                      reg2907 <= $unsigned($signed($unsigned($unsigned(forvar2853))));
                      reg2908 <= $signed(($unsigned((forvar2875 ?
                          forvar2948 : (8'hb8))) + $unsigned((reg2918 | reg2750))));
                      reg2909 <= (reg2768[(1'h1):(1'h1)] >> (reg2764 << ({reg2744} - (~&forvar2845))));
                      reg2910 <= ((8'hb3) < $unsigned((~$signed(reg2927))));
                    end
                  else
                    begin
                      reg2907 <= reg2909;
                      reg2908 <= reg2711[(2'h2):(2'h2)];
                    end
                  if ($signed($signed($unsigned((forvar2875 ?
                      reg1217 : reg2926)))))
                    begin
                      reg2911 <= reg2788;
                      reg2912 <= (~^reg1202[(2'h2):(1'h1)]);
                      reg2913 <= $signed($signed($unsigned(((8'haa) <= forvar2941))));
                    end
                  else
                    begin
                      reg2911 <= $unsigned((forvar2876[(3'h5):(1'h0)] * (!$unsigned(reg2931))));
                      reg2912 <= (-{$signed(forvar2898[(3'h6):(3'h6)])});
                    end
                end
              for (forvar2914 = (1'h0); (forvar2914 < (2'h3)); forvar2914 = (forvar2914 + (1'h1)))
                begin
                  for (forvar2915 = (1'h0); (forvar2915 < (2'h2)); forvar2915 = (forvar2915 + (1'h1)))
                    begin
                      reg2916 <= (reg2716 ^~ {$unsigned((reg2847 >= forvar2914))});
                      reg2917 <= (forvar2875[(1'h0):(1'h0)] ?
                          (|{(reg2847 <= reg2748)}) : $unsigned($signed((&reg2740))));
                      reg2918 <= ($unsigned(forvar2903) ?
                          ($unsigned((reg2813 ? (8'ha0) : reg2805)) ?
                              ((^~forvar2855) >> (~wire1189)) : (~^(forvar2887 == (8'h9f)))) : (reg2849[(1'h0):(1'h0)] < {(reg2785 - reg2925)}));
                    end
                  if ($unsigned(reg2861))
                    begin
                      reg2919 <= (((8'haf) && (8'hae)) ?
                          reg2768[(3'h7):(3'h4)] : reg2844[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg2919 <= (^(~$signed((~&reg1220))));
                      reg2920 <= $signed((reg2947[(2'h2):(2'h2)] ?
                          forvar2932[(3'h7):(3'h7)] : reg2920));
                      reg2921 <= (($signed((reg2821 ? reg2923 : (8'hb9))) ?
                          (~|{forvar2930}) : $unsigned(reg2854[(4'h9):(3'h6)])) << reg2863[(3'h6):(3'h4)]);
                      reg2922 <= $unsigned((reg2922[(3'h4):(2'h3)] ?
                          (!$unsigned(reg2801)) : $unsigned($unsigned(reg2825))));
                    end
                end
            end
        end
      if ((~&reg2862))
        begin
          for (forvar2962 = (1'h0); (forvar2962 < (2'h2)); forvar2962 = (forvar2962 + (1'h1)))
            begin
              reg2963 <= (reg1237[(4'h8):(2'h2)] ^ {(forvar2850[(2'h3):(1'h0)] <= reg2822)});
              for (forvar2964 = (1'h0); (forvar2964 < (1'h1)); forvar2964 = (forvar2964 + (1'h1)))
                begin
                  for (forvar2965 = (1'h0); (forvar2965 < (1'h0)); forvar2965 = (forvar2965 + (1'h1)))
                    begin
                      reg2966 <= (($unsigned($unsigned((8'hb2))) != ($signed(reg2893) & $unsigned(reg2812))) * (reg2717[(1'h0):(1'h0)] < $signed($unsigned(forvar2902))));
                      reg2967 <= forvar2932;
                      reg2968 <= reg1228;
                    end
                  if ($signed((((~^reg2709) ?
                          $unsigned(wire1188) : reg2738[(2'h2):(2'h2)]) ?
                      $unsigned(reg2790[(3'h4):(3'h4)]) : ($signed(reg2894) ?
                          $unsigned(forvar2899) : reg2913))))
                    begin
                      reg2969 <= (forvar2898 + (^~($unsigned(reg2840) <= (8'hb0))));
                      reg2970 <= ({$signed((&reg2891))} ~^ (reg2927[(2'h3):(1'h1)] ?
                          ((8'ha2) - forvar2898) : {(+reg2848)}));
                    end
                  else
                    begin
                      reg2969 <= (((8'hb8) ?
                              $signed((forvar2876 ?
                                  reg2919 : forvar2930)) : reg2892) ?
                          $signed($signed(reg2935[(3'h7):(1'h0)])) : (reg2771[(3'h5):(1'h1)] <= $signed(reg2714[(2'h3):(2'h3)])));
                      reg2970 <= $unsigned(((^{reg2867}) <= ($signed((8'haa)) >= ((8'ha9) && reg2797))));
                      reg2971 <= $signed($signed($unsigned($unsigned(reg2755))));
                      reg2972 <= $signed($unsigned((&wire1190[(3'h6):(2'h2)])));
                    end
                  if ({$unsigned(reg1203)})
                    begin
                      reg2973 <= $signed(($signed($unsigned(reg2897)) + {$unsigned(reg2717)}));
                      reg2974 <= (8'haf);
                      reg2975 <= ((^$unsigned($signed((8'ha3)))) >>> ($unsigned($unsigned(reg2820)) != $signed($unsigned(forvar2965))));
                    end
                  else
                    begin
                      reg2973 <= {$unsigned((((8'hb6) >>> reg2923) ?
                              (^~reg2747) : reg2883))};
                      reg2974 <= {reg2884};
                      reg2975 <= $signed($signed($signed($signed(reg1238))));
                      reg2976 <= (+(reg2756 && $signed($signed(reg2899))));
                    end
                end
            end
          for (forvar2977 = (1'h0); (forvar2977 < (1'h1)); forvar2977 = (forvar2977 + (1'h1)))
            begin
              for (forvar2978 = (1'h0); (forvar2978 < (1'h1)); forvar2978 = (forvar2978 + (1'h1)))
                begin
                  if (((reg2860 << $unsigned(forvar2933)) + (reg2713 ?
                      (forvar2906[(2'h2):(1'h1)] != (reg2940 ?
                          reg1238 : reg2937)) : ((reg2740 ?
                          forvar2948 : reg1210) >>> reg2929[(1'h1):(1'h0)]))))
                    begin
                      reg2979 <= reg2733[(1'h0):(1'h0)];
                      reg2980 <= {(^~forvar2927[(4'he):(4'hc)])};
                      reg2981 <= (~^(reg2848[(4'hd):(3'h7)] ?
                          $unsigned({(8'hac)}) : reg2873));
                    end
                  else
                    begin
                      reg2979 <= reg2711[(1'h1):(1'h1)];
                      reg2980 <= forvar2850[(2'h3):(2'h3)];
                      reg2981 <= (!(^~(~&reg2733)));
                      reg2982 <= (reg2859[(4'hf):(4'ha)] ?
                          (&reg2734[(1'h1):(1'h0)]) : reg2938[(4'ha):(4'h8)]);
                    end
                  if ($signed(reg2728[(2'h2):(2'h2)]))
                    begin
                      reg2983 <= ((($unsigned(reg2815) ?
                              (reg2862 ?
                                  reg1239 : reg2947) : (8'hb6)) > wire1193) ?
                          (wire1189 > reg2827) : reg2982[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg2983 <= (reg2934[(1'h1):(1'h1)] ?
                          reg2934 : ($signed(reg1205) << {reg2760}));
                    end
                  for (forvar2984 = (1'h0); (forvar2984 < (1'h0)); forvar2984 = (forvar2984 + (1'h1)))
                    begin
                      reg2985 <= ((|$unsigned((reg2883 != forvar2927))) ?
                          (~((reg2824 ~^ reg2839) * (forvar2978 ?
                              forvar2933 : reg2975))) : ((+(reg2856 + reg2758)) ?
                              reg2719 : $unsigned(reg2726[(4'ha):(2'h2)])));
                      reg2986 <= ($signed({(reg2825 >= (8'ha4))}) | (-$signed({reg2712})));
                    end
                end
            end
          if (reg2815[(3'h4):(2'h2)])
            begin
              if (((~&(~{(8'h9d)})) == (((reg2937 ~^ forvar2977) ?
                      forvar2908[(2'h3):(2'h3)] : $signed(reg1235)) ?
                  reg2976[(4'hd):(1'h0)] : reg2821)))
                begin
                  for (forvar2987 = (1'h0); (forvar2987 < (1'h0)); forvar2987 = (forvar2987 + (1'h1)))
                    begin
                      reg2988 <= (forvar2932 != {$unsigned((reg2861 ?
                              reg2857 : reg2896))});
                      reg2989 <= reg2737[(4'hb):(1'h1)];
                      reg2990 <= $signed(reg2903);
                    end
                end
              else
                begin
                  if (reg1239[(4'hf):(2'h3)])
                    begin
                      reg2987 <= reg2967[(1'h0):(1'h0)];
                      reg2988 <= (^~({(-reg2966)} == $signed((!reg2878))));
                      reg2989 <= $signed($signed(forvar2887[(3'h7):(3'h5)]));
                      reg2990 <= $unsigned($signed(reg2742));
                    end
                  else
                    begin
                      reg2987 <= forvar2959[(3'h5):(2'h3)];
                      reg2988 <= (~^(8'hb7));
                      reg2989 <= (+(((~|reg2895) <<< reg2752) * $unsigned($signed(reg2893))));
                    end
                  for (forvar2991 = (1'h0); (forvar2991 < (2'h3)); forvar2991 = (forvar2991 + (1'h1)))
                    begin
                      reg2992 <= reg2813[(3'h6):(3'h4)];
                      reg2993 <= $unsigned($unsigned({reg2740[(2'h3):(2'h3)]}));
                      reg2994 <= reg2725[(3'h6):(2'h2)];
                    end
                end
              for (forvar2995 = (1'h0); (forvar2995 < (1'h0)); forvar2995 = (forvar2995 + (1'h1)))
                begin
                  for (forvar2996 = (1'h0); (forvar2996 < (1'h0)); forvar2996 = (forvar2996 + (1'h1)))
                    begin
                      reg2997 <= reg2788[(3'h6):(3'h4)];
                      reg2998 <= (^~reg2945);
                      reg2999 <= (~{(~reg2717)});
                      reg3000 <= {reg2724[(3'h4):(1'h1)]};
                    end
                  if (($unsigned((reg2731 ^~ ((8'ha8) ?
                      reg2985 : reg2953))) != (^~({(8'ha1)} & ((8'hb9) | forvar2917)))))
                    begin
                      reg3001 <= $signed(reg2942[(2'h2):(2'h2)]);
                      reg3002 <= ($unsigned($signed((reg2708 || forvar2838))) >> ((8'hac) ?
                          {reg1223} : reg2847));
                      reg3003 <= (8'hb1);
                    end
                  else
                    begin
                      reg3001 <= (^$unsigned(reg2956[(3'h6):(3'h4)]));
                      reg3002 <= ($unsigned(reg2715) ?
                          $unsigned($unsigned(reg2869)) : $unsigned(reg2979));
                      reg3003 <= reg2867;
                    end
                  if (($unsigned({(reg2795 >>> reg2836)}) ?
                      $unsigned((((8'ha8) ?
                          reg2826 : forvar2850) > (wire2837 >>> forvar2839))) : $unsigned($unsigned($unsigned(reg2829)))))
                    begin
                      reg3004 <= (8'ha5);
                      reg3005 <= $unsigned((reg2901[(1'h1):(1'h1)] ?
                          $signed((reg2716 ?
                              forvar2851 : reg2788)) : (((8'h9d) ?
                                  reg2848 : reg2795) ?
                              reg1199[(1'h0):(1'h0)] : reg2974[(2'h2):(1'h1)])));
                      reg3006 <= (reg2860[(3'h6):(2'h3)] ?
                          ((+$signed(reg2840)) ^~ {(|reg3000)}) : (reg2985[(4'hc):(4'ha)] ^ ($signed(reg2738) ?
                              {forvar2875} : ((8'had) ? reg2748 : reg2908))));
                    end
                  else
                    begin
                      reg3004 <= $unsigned(reg2911);
                      reg3005 <= ($unsigned({reg2826[(1'h1):(1'h1)]}) & $signed($signed((reg2922 ?
                          wire1189 : forvar2918))));
                      reg3006 <= ({reg2985[(3'h4):(2'h2)]} ?
                          {reg2762} : reg2751);
                    end
                end
              if (($unsigned(($signed(forvar2906) ?
                      (reg2920 ? reg2838 : reg2957) : $unsigned((8'hb5)))) ?
                  ((~|(reg2761 ?
                      forvar2891 : forvar2926)) << reg2708) : {{reg2972[(3'h5):(1'h0)]}}))
                begin
                  for (forvar3007 = (1'h0); (forvar3007 < (1'h0)); forvar3007 = (forvar3007 + (1'h1)))
                    begin
                      reg3008 <= ((!reg2738) ?
                          $unsigned(((&reg2780) ?
                              (reg1215 ^ reg2779) : reg2972[(3'h7):(3'h5)])) : $unsigned((-{(8'hb3)})));
                    end
                  if ((~(-reg2824[(4'h8):(4'h8)])))
                    begin
                      reg3009 <= $signed(reg1209[(4'ha):(2'h3)]);
                      reg3010 <= $unsigned(((&$unsigned(forvar2843)) ?
                          forvar2899 : {((8'haa) ? forvar2862 : reg2775)}));
                      reg3011 <= (+$signed(reg2791));
                    end
                  else
                    begin
                      reg3009 <= $signed((8'hab));
                      reg3010 <= $signed((reg1199[(2'h3):(2'h3)] != $signed(forvar2875[(3'h4):(1'h0)])));
                      reg3011 <= wire1190;
                      reg3012 <= (&(($signed(forvar2962) ?
                              {(8'hab)} : $signed((8'ha8))) ?
                          $unsigned($unsigned(reg2840)) : ((~^reg2729) ?
                              $signed(reg2911) : (~reg2812))));
                    end
                  for (forvar3013 = (1'h0); (forvar3013 < (2'h3)); forvar3013 = (forvar3013 + (1'h1)))
                    begin
                      reg3014 <= ((+(reg2914 <<< reg2973[(2'h3):(2'h3)])) != reg1228);
                      reg3015 <= reg2926;
                      reg3016 <= ($signed({(~|reg1234)}) ?
                          ({(^reg2903)} ?
                              reg2924 : forvar2862) : $signed((|$unsigned(reg2847))));
                    end
                end
              else
                begin
                  if ((|forvar2881))
                    begin
                      reg3007 <= {((~^$unsigned(reg1208)) > ($signed((8'hab)) ?
                              (reg2783 ?
                                  reg2859 : reg1198) : $unsigned(forvar2908)))};
                      reg3008 <= $unsigned(reg2979);
                      reg3009 <= ({$unsigned(forvar2978)} ?
                          ({(forvar2890 ? reg1200 : reg2777)} ?
                              {((8'h9e) * (8'ha7))} : ($unsigned(reg3002) <<< $unsigned(forvar2861))) : ({reg2811[(2'h3):(1'h1)]} ^ reg1205[(3'h6):(3'h6)]));
                      reg3010 <= (({$signed(reg2715)} & (reg2835 != (forvar2944 >>> forvar2860))) && forvar2933[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg3007 <= $unsigned(reg2924);
                      reg3008 <= $unsigned(reg2989[(1'h0):(1'h0)]);
                    end
                  for (forvar3011 = (1'h0); (forvar3011 < (2'h2)); forvar3011 = (forvar3011 + (1'h1)))
                    begin
                      reg3012 <= $unsigned((((|reg2783) | (reg2979 ?
                              reg2943 : reg2878)) ?
                          forvar2855[(1'h1):(1'h0)] : (|reg2970)));
                      reg3013 <= reg2749[(4'h9):(1'h0)];
                      reg3014 <= ($unsigned(forvar2899) >>> ((&(-(8'h9c))) ?
                          ((&reg2869) ?
                              ((8'h9f) ?
                                  reg2759 : reg2882) : (reg2757 & reg2926)) : ($signed(reg2708) ?
                              (reg2820 ?
                                  reg2926 : forvar2862) : reg2983[(2'h2):(1'h1)])));
                      reg3015 <= {$unsigned($signed(forvar2859[(4'h8):(1'h0)]))};
                    end
                  if ((^reg2957))
                    begin
                      reg3016 <= ($signed({{reg2824}}) ?
                          ((reg2716[(2'h3):(2'h3)] != forvar2962) ~^ ((reg3000 >= reg2946) ?
                              (reg2928 ?
                                  reg2895 : forvar2987) : (reg2908 | (8'hb3)))) : $signed(((reg2862 ^ reg2748) ?
                              {forvar2840} : $signed(reg2960))));
                      reg3017 <= (reg2720 & reg3008[(1'h0):(1'h0)]);
                      reg3018 <= forvar2859[(4'he):(4'he)];
                      reg3019 <= reg1233;
                    end
                  else
                    begin
                      reg3016 <= (~^$signed(((reg2899 >>> (8'ha5)) ?
                          $unsigned(wire1193) : {reg2945})));
                    end
                end
            end
          else
            begin
              if (reg2725)
                begin
                  for (forvar2987 = (1'h0); (forvar2987 < (1'h0)); forvar2987 = (forvar2987 + (1'h1)))
                    begin
                      reg2988 <= $signed(($signed(reg2979[(1'h1):(1'h1)]) ?
                          $signed((reg2712 ?
                              reg2742 : reg2761)) : forvar2920[(2'h2):(1'h1)]));
                      reg2989 <= (-(wire1190[(3'h7):(3'h4)] <<< reg2918[(3'h4):(2'h2)]));
                      reg2990 <= $signed(reg2778);
                      reg2991 <= forvar2901;
                    end
                  if ({$signed($unsigned((^reg2811)))})
                    begin
                      reg2992 <= reg2847;
                      reg2993 <= ({{(-reg2737)}} != $unsigned((!(reg2945 ?
                          reg1202 : reg2787))));
                      reg2994 <= ($unsigned((~&$signed(reg2910))) ?
                          reg1233 : ((reg2732[(2'h3):(2'h3)] <= $signed(reg2805)) ^~ $unsigned((~^reg2899))));
                    end
                  else
                    begin
                      reg2992 <= $unsigned((&{$unsigned(reg2779)}));
                    end
                end
              else
                begin
                  if (((&reg2807[(1'h0):(1'h0)]) >> $unsigned($signed((reg1202 ~^ forvar2977)))))
                    begin
                      reg2987 <= ($unsigned($signed(forvar2890[(3'h5):(2'h2)])) ?
                          $unsigned(reg1235) : (reg2937 ?
                              reg2725 : (((8'hb0) ? reg2721 : (8'ha1)) ?
                                  reg1230[(2'h2):(2'h2)] : $unsigned(reg2763))));
                      reg2988 <= wire1190;
                      reg2989 <= reg2979;
                      reg2990 <= ($signed(reg2922[(3'h5):(3'h5)]) ?
                          (-$signed((8'h9c))) : (((reg1234 < reg2993) ?
                                  $unsigned(reg2877) : reg1216) ?
                              (~(reg2840 ?
                                  reg2900 : forvar2839)) : ($unsigned(reg2864) <= {reg2999})));
                    end
                  else
                    begin
                      reg2987 <= $unsigned((reg2838[(4'h9):(2'h3)] ?
                          $unsigned(forvar2964[(4'ha):(3'h5)]) : (~$signed(reg2902))));
                      reg2988 <= $unsigned((-reg2953[(3'h4):(1'h0)]));
                      reg2989 <= $signed((({reg1226} >>> (reg2991 ?
                          reg2744 : reg2822)) && ($unsigned(reg2771) ?
                          {(8'ha8)} : $signed((8'hac)))));
                      reg2990 <= $unsigned(reg2914[(3'h4):(1'h1)]);
                    end
                  for (forvar2991 = (1'h0); (forvar2991 < (2'h2)); forvar2991 = (forvar2991 + (1'h1)))
                    begin
                      reg2992 <= reg2725[(3'h5):(1'h1)];
                    end
                end
            end
          reg3020 <= reg2879[(3'h7):(3'h7)];
        end
      else
        begin
          if ({(~|((reg2761 ? reg1239 : reg2800) ?
                  reg2991[(1'h1):(1'h1)] : {reg2966}))})
            begin
              for (forvar2962 = (1'h0); (forvar2962 < (1'h1)); forvar2962 = (forvar2962 + (1'h1)))
                begin
                  for (forvar2963 = (1'h0); (forvar2963 < (1'h1)); forvar2963 = (forvar2963 + (1'h1)))
                    begin
                      reg2964 <= (&$unsigned(($signed(wire1189) ?
                          $unsigned(reg2869) : (reg2908 || reg2757))));
                      reg2965 <= reg1229[(3'h5):(1'h0)];
                      reg2966 <= (~(^~$signed((reg2981 ? reg2814 : reg3016))));
                      reg2967 <= (~^($unsigned((reg2793 ?
                          reg1202 : forvar2959)) && (~^(&reg2951))));
                    end
                  if (reg2739[(2'h3):(2'h3)])
                    begin
                      reg2968 <= (+$signed((reg3012[(1'h0):(1'h0)] ?
                          (reg1197 >> reg3015) : (&(8'hb1)))));
                      reg2969 <= (8'hac);
                    end
                  else
                    begin
                      reg2968 <= (&$signed((8'ha0)));
                    end
                end
              if ($signed(($signed($unsigned(reg2888)) ?
                  (+(forvar2926 >> wire1189)) : ($signed(reg1222) ~^ $unsigned(reg2714)))))
                begin
                  if ($unsigned(((^reg2951[(4'ha):(4'ha)]) != {forvar2927[(3'h4):(1'h1)]})))
                    begin
                      reg2970 <= {(forvar2996 >= ($unsigned((8'hb3)) != (&reg2986)))};
                      reg2971 <= (~(!$unsigned(((8'hba) ^~ reg2923))));
                    end
                  else
                    begin
                      reg2970 <= reg2988;
                      reg2971 <= $unsigned((reg1220[(2'h3):(2'h3)] && $unsigned({(8'hb2)})));
                    end
                  if ((reg2831[(2'h2):(2'h2)] | {(^{reg2863})}))
                    begin
                      reg2972 <= ({(reg2801[(3'h5):(1'h0)] == $signed((8'ha9)))} ^ {reg2909});
                      reg2973 <= (|forvar2852);
                      reg2974 <= (reg2930[(4'h8):(3'h5)] ?
                          (forvar2890[(3'h5):(1'h1)] ^ forvar2912) : ((~&((8'ha5) ?
                                  reg2844 : wire1193)) ?
                              (|(8'ha9)) : {(forvar2926 ^ reg3001)}));
                      reg2975 <= reg2721;
                    end
                  else
                    begin
                      reg2972 <= {reg2968};
                    end
                  for (forvar2976 = (1'h0); (forvar2976 < (1'h1)); forvar2976 = (forvar2976 + (1'h1)))
                    begin
                      reg2977 <= wire2837[(3'h5):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar2970 = (1'h0); (forvar2970 < (2'h3)); forvar2970 = (forvar2970 + (1'h1)))
                    begin
                      reg2971 <= (|(|reg2971));
                      reg2972 <= ($signed($signed((+reg2834))) ?
                          {{reg2797}} : (^~($signed(forvar2965) ^ (reg2810 ?
                              reg2824 : reg1238))));
                    end
                end
            end
          else
            begin
              reg2962 <= ({$unsigned((~&reg2719))} ^~ $signed((reg2846[(1'h1):(1'h0)] ?
                  (~^(8'h9c)) : {forvar2976})));
              reg2963 <= $unsigned(reg1219);
            end
          for (forvar2978 = (1'h0); (forvar2978 < (1'h0)); forvar2978 = (forvar2978 + (1'h1)))
            begin
              for (forvar2979 = (1'h0); (forvar2979 < (1'h0)); forvar2979 = (forvar2979 + (1'h1)))
                begin
                  if (reg2820[(2'h3):(2'h2)])
                    begin
                      reg2980 <= reg2931[(1'h1):(1'h0)];
                      reg2981 <= $unsigned(reg2754[(2'h2):(1'h0)]);
                      reg2982 <= reg2756;
                      reg2983 <= {(((reg2808 >= forvar2853) + (~forvar2920)) && $unsigned(reg2945[(2'h3):(2'h2)]))};
                    end
                  else
                    begin
                      reg2980 <= forvar2987;
                    end
                  if ({$signed($signed($unsigned(reg1215)))})
                    begin
                      reg2984 <= {(({reg2833} ?
                              (~|(8'h9e)) : ((8'ha3) != forvar2915)) << (|(~^reg2974)))};
                      reg2985 <= ($signed(forvar2902[(3'h7):(3'h7)]) >= ((reg2711[(1'h0):(1'h0)] ?
                          reg2838[(4'hc):(3'h6)] : $signed(reg2849)) << $unsigned((wire2837 ~^ reg2873))));
                      reg2986 <= reg2960;
                      reg2987 <= $signed($unsigned({(|reg2851)}));
                    end
                  else
                    begin
                      reg2984 <= {reg2923[(3'h7):(2'h2)]};
                      reg2985 <= $unsigned($signed(({(8'hb7)} ?
                          (+reg2953) : forvar2845[(2'h2):(1'h1)])));
                      reg2986 <= {$signed($unsigned((reg2848 ?
                              (8'ha1) : reg2966)))};
                      reg2987 <= (!(-((reg2936 ? reg2802 : reg2956) ?
                          $unsigned(reg2977) : (reg2994 * forvar3011))));
                    end
                end
              reg2988 <= reg2840;
            end
          if ((~^$signed(reg2935)))
            begin
              for (forvar2989 = (1'h0); (forvar2989 < (1'h1)); forvar2989 = (forvar2989 + (1'h1)))
                begin
                  for (forvar2990 = (1'h0); (forvar2990 < (1'h0)); forvar2990 = (forvar2990 + (1'h1)))
                    begin
                      reg2991 <= reg2888;
                      reg2992 <= forvar2926;
                      reg2993 <= (~&((+((8'had) ?
                          reg2991 : reg2781)) <= forvar2920));
                    end
                  for (forvar2994 = (1'h0); (forvar2994 < (2'h3)); forvar2994 = (forvar2994 + (1'h1)))
                    begin
                      reg2995 <= ($signed((reg2829 ?
                          $signed(reg2921) : {reg2797})) | $signed({(|reg2939)}));
                    end
                  if ($signed(reg2842))
                    begin
                      reg2996 <= $signed($unsigned($unsigned($unsigned(reg2910))));
                      reg2997 <= (!(&((reg1222 > reg2993) ?
                          $signed((8'ha4)) : $signed(reg2798))));
                    end
                  else
                    begin
                      reg2996 <= (forvar2978 || $signed($unsigned(reg3017[(4'h9):(4'h9)])));
                      reg2997 <= ((reg2746 && reg2796) || $signed($unsigned($unsigned(reg2846))));
                      reg2998 <= ((~|((reg2860 && reg1217) ?
                          ((8'h9e) ?
                              reg2725 : reg1226) : (8'ha7))) * ((~^forvar2979) ?
                          {$signed((8'ha0))} : $signed(reg2925[(4'h8):(4'h8)])));
                      reg2999 <= (~|$unsigned((~^(reg2757 > forvar2994))));
                    end
                end
              for (forvar3000 = (1'h0); (forvar3000 < (2'h3)); forvar3000 = (forvar3000 + (1'h1)))
                begin
                  for (forvar3001 = (1'h0); (forvar3001 < (1'h0)); forvar3001 = (forvar3001 + (1'h1)))
                    begin
                      reg3002 <= (reg2796[(3'h5):(1'h0)] ?
                          (~forvar2920) : $unsigned((reg2770[(2'h3):(1'h1)] ?
                              (forvar2930 == reg2720) : forvar2994)));
                      reg3003 <= (-($signed(reg2908[(1'h1):(1'h1)]) ~^ (8'hb9)));
                      reg3004 <= reg2775[(4'h8):(1'h0)];
                      reg3005 <= reg2857[(4'ha):(2'h3)];
                    end
                  if (((($unsigned(reg2734) && (reg2739 ?
                      forvar2891 : reg2970)) - reg2802) << $unsigned($unsigned({forvar2850}))))
                    begin
                      reg3006 <= reg2946;
                      reg3007 <= $signed((~$signed(forvar2978)));
                    end
                  else
                    begin
                      reg3006 <= ($unsigned(reg2777) ~^ $unsigned({(reg2980 >>> reg2934)}));
                      reg3007 <= $unsigned(reg2866[(4'h8):(2'h3)]);
                    end
                  if (($signed(((reg2826 && forvar2851) == reg2769[(4'hd):(3'h7)])) <= reg2968[(1'h0):(1'h0)]))
                    begin
                      reg3008 <= $unsigned((reg2790[(2'h3):(1'h1)] ?
                          (8'hae) : reg2755[(2'h2):(1'h0)]));
                      reg3009 <= reg1216;
                    end
                  else
                    begin
                      reg3008 <= $unsigned(reg2928[(1'h0):(1'h0)]);
                      reg3009 <= $unsigned(forvar2857[(3'h5):(3'h5)]);
                      reg3010 <= reg1208[(4'hc):(4'h9)];
                    end
                  reg3011 <= (reg3012[(3'h6):(1'h0)] * ((~(~|reg2934)) >= reg2749[(1'h0):(1'h0)]));
                end
            end
          else
            begin
              if ($unsigned($unsigned({forvar2903[(4'hd):(4'h9)]})))
                begin
                  for (forvar2989 = (1'h0); (forvar2989 < (2'h3)); forvar2989 = (forvar2989 + (1'h1)))
                    begin
                      reg2990 <= reg2798;
                      reg2991 <= $signed($signed(($unsigned(reg3003) ?
                          (reg2732 ? reg1228 : reg2857) : reg2853)));
                      reg2992 <= ($signed((~(|(8'hb0)))) ?
                          $unsigned($unsigned(((8'h9f) > reg2867))) : reg2960[(2'h2):(1'h0)]);
                      reg2993 <= (~^(((reg3016 ? reg2842 : (8'hb9)) ?
                          reg2724[(3'h5):(1'h1)] : (~|reg2921)) < forvar3007));
                    end
                  if ((reg2805 <= reg2786))
                    begin
                      reg2994 <= ({(~$signed(reg1209))} ?
                          ($unsigned($unsigned(forvar2864)) * $unsigned(reg1228)) : (reg2719 | reg1226[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg2994 <= reg2931;
                    end
                  reg2995 <= $signed($unsigned(reg2783[(4'h9):(3'h4)]));
                end
              else
                begin
                  for (forvar2989 = (1'h0); (forvar2989 < (1'h0)); forvar2989 = (forvar2989 + (1'h1)))
                    begin
                      reg2990 <= $unsigned((forvar2996[(3'h4):(2'h2)] + forvar2970));
                      reg2991 <= ((8'hb9) > $unsigned(((8'hba) ~^ $signed(reg2836))));
                    end
                end
              if ((^forvar2927[(1'h0):(1'h0)]))
                begin
                  if ({reg1200[(1'h1):(1'h1)]})
                    begin
                      reg2996 <= (+reg2937);
                      reg2997 <= reg2993[(4'he):(3'h7)];
                    end
                  else
                    begin
                      reg2996 <= (reg1239 && ($signed((reg1202 ?
                              reg2834 : reg2957)) ?
                          {(reg1229 >> forvar2962)} : (reg2981 ~^ $unsigned(forvar2887))));
                      reg2997 <= ($unsigned(forvar2962[(2'h2):(2'h2)]) ?
                          (8'h9f) : $unsigned(((reg2954 ?
                                  reg2942 : forvar2881) ?
                              $signed((8'hb5)) : $signed(reg2929))));
                    end
                end
              else
                begin
                  reg2996 <= (reg2985 ?
                      ((~reg3018[(1'h0):(1'h0)]) ?
                          {reg2778[(3'h6):(1'h0)]} : $unsigned({reg2768})) : ($unsigned(reg2999[(1'h1):(1'h0)]) ?
                          ((forvar2874 != (8'hb0)) == (reg1227 != forvar2915)) : ((reg2982 >>> reg2865) ?
                              $unsigned(wire1193) : {reg2747})));
                end
              if ((({(8'ha4)} ~^ (&$unsigned(reg3005))) | (-forvar2984[(4'h8):(3'h5)])))
                begin
                  for (forvar2998 = (1'h0); (forvar2998 < (1'h1)); forvar2998 = (forvar2998 + (1'h1)))
                    begin
                      reg2999 <= ((((reg2897 << reg1230) ?
                              reg2841[(3'h4):(1'h1)] : $unsigned(forvar2952)) ~^ {$unsigned(forvar2941)}) ?
                          reg2749 : {{(&reg3017)}});
                      reg3000 <= reg2981;
                      reg3001 <= $unsigned($unsigned($unsigned((^~reg2819))));
                      reg3002 <= (|reg2848[(4'h9):(3'h6)]);
                    end
                  reg3003 <= $signed($signed(((^~(8'hac)) ?
                      {forvar2964} : (reg2724 * reg2973))));
                end
              else
                begin
                  if (reg2722[(1'h1):(1'h0)])
                    begin
                      reg2998 <= $unsigned((reg2993 ?
                          reg2737 : $signed((^~reg2739))));
                    end
                  else
                    begin
                      reg2998 <= {reg2744};
                    end
                  for (forvar2999 = (1'h0); (forvar2999 < (1'h1)); forvar2999 = (forvar2999 + (1'h1)))
                    begin
                      reg3000 <= $signed((~reg2926));
                      reg3001 <= (8'hb5);
                      reg3002 <= ((&($signed((8'haa)) || $unsigned(reg3010))) > ($signed($signed((8'h9c))) * reg2958));
                    end
                  if ({(!(((8'hac) ? forvar2930 : reg1237) <<< (reg2712 ?
                          reg3014 : reg2719)))})
                    begin
                      reg3003 <= (8'ha7);
                      reg3004 <= $unsigned({$unsigned((reg2966 ?
                              (8'ha3) : reg2943))});
                      reg3005 <= ((reg2958[(3'h4):(2'h2)] ?
                          ((~|reg2821) ^ reg2947[(1'h1):(1'h0)]) : forvar2838[(4'h9):(4'h8)]) && $signed($signed((reg1214 ?
                          reg2729 : forvar2906))));
                    end
                  else
                    begin
                      reg3003 <= ((~|($signed((8'ha0)) < (reg2709 < reg2882))) <<< reg2860);
                    end
                end
              if ({(^(|(reg3001 ? reg2756 : reg2935)))})
                begin
                  reg3006 <= reg2760;
                  for (forvar3007 = (1'h0); (forvar3007 < (1'h0)); forvar3007 = (forvar3007 + (1'h1)))
                    begin
                      reg3008 <= {(forvar2845[(4'hb):(3'h6)] <<< {$unsigned(reg2981)})};
                    end
                end
              else
                begin
                  if ((8'ha9))
                    begin
                      reg3006 <= ($unsigned($signed((^reg2710))) ?
                          ((~^reg1209) + ((reg2747 < (8'hb0)) ?
                              forvar3007[(1'h1):(1'h1)] : forvar2998[(2'h2):(2'h2)])) : forvar2875[(3'h7):(3'h5)]);
                      reg3007 <= $signed(($signed($signed(reg2899)) ^ (reg2976 ?
                          $unsigned((8'hae)) : $signed(reg2970))));
                    end
                  else
                    begin
                      reg3006 <= ((-((reg2830 ?
                              reg2735 : reg2986) ^~ (reg2963 & reg2835))) ?
                          (((~&reg2950) != reg2862[(1'h1):(1'h0)]) >= reg2925[(3'h7):(2'h2)]) : (~&$signed(forvar3000[(4'hf):(4'hf)])));
                      reg3007 <= reg2775;
                      reg3008 <= ((reg2801 >= reg2747) ^~ $unsigned($unsigned({(8'h9f)})));
                      reg3009 <= $signed({({reg2957} ?
                              {forvar2978} : (reg2970 ? reg2914 : (8'ha4)))});
                    end
                  if ($signed((({reg2780} ? (!reg2820) : $unsigned(reg2950)) ?
                      ((reg2849 ?
                          reg1237 : reg2835) || ((8'hb4) >> forvar2948)) : ((~&reg1227) | (reg2847 || reg2761)))))
                    begin
                      reg3010 <= $signed({$unsigned(reg2749[(3'h4):(1'h1)])});
                      reg3011 <= $signed((|{forvar2941[(3'h5):(1'h1)]}));
                      reg3012 <= {($signed((~&forvar2890)) ?
                              {reg2922} : ((!reg2719) ?
                                  forvar2977[(4'hc):(2'h2)] : $unsigned(reg2851)))};
                    end
                  else
                    begin
                      reg3010 <= {reg2795[(1'h1):(1'h1)]};
                      reg3011 <= (reg2891 ?
                          ($signed(forvar2930) != $unsigned(reg2882)) : $unsigned((forvar2998[(3'h5):(2'h2)] ?
                              $signed(reg2780) : reg2769)));
                      reg3012 <= reg1238[(1'h1):(1'h1)];
                    end
                  for (forvar3013 = (1'h0); (forvar3013 < (2'h3)); forvar3013 = (forvar3013 + (1'h1)))
                    begin
                      reg3014 <= reg1220;
                      reg3015 <= ($signed(reg3004) ?
                          (((reg3007 << reg2947) > (reg2909 >= reg1226)) >> ($unsigned(reg2854) ?
                              (reg2855 ?
                                  reg2709 : reg2738) : $signed(reg2746))) : ($unsigned(forvar2901[(1'h1):(1'h0)]) * forvar3007));
                    end
                end
            end
        end
    end
  assign wire3021 = reg2758[(4'h9):(1'h0)];
  always
    @(posedge clk) begin
      reg3022 <= $signed($unsigned(($signed(reg2878) <<< (reg2905 ?
          reg2859 : reg2907))));
      if ($signed(reg2972))
        begin
          for (forvar3023 = (1'h0); (forvar3023 < (2'h2)); forvar3023 = (forvar3023 + (1'h1)))
            begin
              if ($unsigned($unsigned({{reg3010}})))
                begin
                  for (forvar3024 = (1'h0); (forvar3024 < (2'h3)); forvar3024 = (forvar3024 + (1'h1)))
                    begin
                      reg3025 <= $signed(($unsigned(reg2753[(3'h6):(2'h2)]) ?
                          (~|(reg2999 ? reg2803 : (8'h9d))) : wire1241));
                      reg3026 <= $unsigned({(^~reg2894)});
                      reg3027 <= (^~(8'hb0));
                    end
                  if ((^~reg2859[(3'h6):(1'h1)]))
                    begin
                      reg3028 <= wire1192;
                    end
                  else
                    begin
                      reg3028 <= $unsigned(wire2706);
                      reg3029 <= reg2893;
                      reg3030 <= reg2820[(2'h2):(2'h2)];
                      reg3031 <= reg3003;
                    end
                end
              else
                begin
                  reg3024 <= (^reg2999[(1'h1):(1'h0)]);
                  for (forvar3025 = (1'h0); (forvar3025 < (1'h1)); forvar3025 = (forvar3025 + (1'h1)))
                    begin
                      reg3026 <= (($unsigned(((8'hab) ? reg2860 : reg1228)) ?
                          {$unsigned(reg2783)} : ($signed(reg1199) ^~ ((8'ha2) ?
                              reg2946 : reg2924))) ~^ reg2735[(2'h3):(2'h3)]);
                      reg3027 <= $unsigned(reg2796);
                      reg3028 <= $signed((^~reg2997));
                    end
                  reg3029 <= $unsigned((((^~reg2930) ?
                          $unsigned(reg1234) : (&reg2780)) ?
                      (~^(reg2916 | reg2871)) : $unsigned($signed(reg2883))));
                end
            end
          if ({(|$signed($signed(reg2966)))})
            begin
              reg3032 <= $unsigned(reg2908);
              for (forvar3033 = (1'h0); (forvar3033 < (2'h3)); forvar3033 = (forvar3033 + (1'h1)))
                begin
                  reg3034 <= ({$signed((~|reg2822))} ?
                      $signed(reg2908[(4'ha):(3'h6)]) : (reg2968 ?
                          (8'hb4) : $unsigned($signed(reg3019))));
                end
              for (forvar3035 = (1'h0); (forvar3035 < (2'h2)); forvar3035 = (forvar3035 + (1'h1)))
                begin
                  for (forvar3036 = (1'h0); (forvar3036 < (1'h0)); forvar3036 = (forvar3036 + (1'h1)))
                    begin
                      reg3037 <= reg2991;
                    end
                  for (forvar3038 = (1'h0); (forvar3038 < (2'h3)); forvar3038 = (forvar3038 + (1'h1)))
                    begin
                      reg3039 <= reg2864[(2'h3):(1'h1)];
                      reg3040 <= ($signed((reg2995 * (+reg2761))) ?
                          $unsigned($signed((reg2918 <<< (8'hac)))) : $signed(reg2964));
                      reg3041 <= $signed({reg2988[(3'h7):(3'h4)]});
                    end
                end
              for (forvar3042 = (1'h0); (forvar3042 < (2'h2)); forvar3042 = (forvar3042 + (1'h1)))
                begin
                  for (forvar3043 = (1'h0); (forvar3043 < (1'h1)); forvar3043 = (forvar3043 + (1'h1)))
                    begin
                      reg3044 <= $signed(reg2769[(4'he):(4'hc)]);
                      reg3045 <= (~$unsigned(((reg2828 ?
                          reg2788 : reg2829) ^~ reg2740[(1'h1):(1'h1)])));
                      reg3046 <= (($unsigned((^(8'hae))) | (reg2928[(2'h3):(1'h1)] != reg2779)) ?
                          {reg2871[(2'h3):(2'h3)]} : $signed(reg2833[(4'hc):(4'hc)]));
                      reg3047 <= $unsigned(((8'hab) == {$unsigned(reg2800)}));
                    end
                end
            end
          else
            begin
              if ($unsigned(reg2724[(1'h1):(1'h1)]))
                begin
                  if (forvar3038)
                    begin
                      reg3032 <= reg1238[(2'h2):(1'h1)];
                      reg3033 <= $signed($signed((+reg2815)));
                      reg3034 <= reg2905;
                      reg3035 <= (reg3022[(1'h0):(1'h0)] & reg2766[(4'hb):(4'h8)]);
                    end
                  else
                    begin
                      reg3032 <= $signed($signed({(reg2846 ?
                              reg2850 : reg2815)}));
                      reg3033 <= (8'ha4);
                      reg3034 <= ($signed($signed($unsigned(reg2738))) << $signed(reg2882[(1'h1):(1'h1)]));
                    end
                  for (forvar3036 = (1'h0); (forvar3036 < (2'h3)); forvar3036 = (forvar3036 + (1'h1)))
                    begin
                      reg3037 <= $unsigned(reg2735[(2'h2):(2'h2)]);
                      reg3038 <= $unsigned((|(~^$unsigned(reg2757))));
                      reg3039 <= (&reg2906[(3'h5):(3'h5)]);
                    end
                end
              else
                begin
                  for (forvar3032 = (1'h0); (forvar3032 < (2'h3)); forvar3032 = (forvar3032 + (1'h1)))
                    begin
                      reg3033 <= reg2714[(3'h6):(3'h6)];
                      reg3034 <= reg2839;
                    end
                end
            end
        end
      else
        begin
          reg3023 <= ((reg2785[(4'h8):(3'h6)] & reg2982) ?
              {(^~(8'hb1))} : {$signed(reg2712[(2'h2):(2'h2)])});
          if ($signed((+$unsigned($unsigned((8'h9e))))))
            begin
              reg3024 <= reg2757[(4'ha):(3'h6)];
              reg3025 <= forvar3042[(3'h5):(1'h0)];
            end
          else
            begin
              if (((+(+reg2975)) ? reg1208 : $unsigned({$signed(reg2747)})))
                begin
                  reg3024 <= $signed($unsigned($unsigned({(8'ha1)})));
                  reg3025 <= reg2957[(2'h2):(1'h0)];
                end
              else
                begin
                  if (reg2896)
                    begin
                      reg3024 <= ({$signed((reg3038 ? (8'hae) : reg3037))} ?
                          ((~^$signed(reg1228)) > reg2888[(1'h0):(1'h0)]) : ($signed((reg1198 && reg2740)) * (!reg3019)));
                      reg3025 <= reg3005[(4'h9):(3'h4)];
                      reg3026 <= ($unsigned($signed(reg2742[(3'h5):(3'h4)])) ?
                          reg2734[(3'h5):(2'h2)] : reg2896);
                      reg3027 <= reg2863;
                    end
                  else
                    begin
                      reg3024 <= reg2906;
                      reg3025 <= $signed(((reg2923[(3'h4):(2'h3)] ?
                              $signed(reg2757) : (reg2853 >>> reg2972)) ?
                          $unsigned($signed(reg3004)) : reg3017[(3'h5):(2'h3)]));
                      reg3026 <= reg2903;
                      reg3027 <= $signed((reg3002[(3'h5):(3'h5)] ?
                          $unsigned($unsigned(reg2921)) : reg2759));
                    end
                  for (forvar3028 = (1'h0); (forvar3028 < (2'h2)); forvar3028 = (forvar3028 + (1'h1)))
                    begin
                      reg3029 <= ({$signed((~|reg2969))} << reg2947);
                      reg3030 <= (wire2837[(2'h3):(1'h1)] ?
                          $unsigned((^reg3032[(2'h3):(1'h1)])) : $unsigned((reg1197[(3'h7):(1'h1)] & $signed((8'ha4)))));
                      reg3031 <= $unsigned((^$unsigned($signed(reg2979))));
                      reg3032 <= reg2754[(1'h0):(1'h0)];
                    end
                end
            end
          reg3033 <= ((({(8'hac)} ?
              (8'hb1) : wire2837[(1'h0):(1'h0)]) <<< $unsigned((reg2817 ~^ reg2974))) != (($signed((8'hb7)) | ((8'ha2) == reg2916)) ?
              {reg2894[(4'h8):(3'h4)]} : $signed($signed((8'hae)))));
          if ($signed({reg2971[(1'h0):(1'h0)]}))
            begin
              if ((reg2842[(3'h5):(1'h0)] ? (^(^~$signed(reg2814))) : (8'hb7)))
                begin
                  if (((reg2910[(1'h0):(1'h0)] ? reg2884 : $signed(reg2772)) ?
                      reg2934[(1'h1):(1'h0)] : (^((!reg2957) || (8'hb0)))))
                    begin
                      reg3034 <= reg2980[(4'h9):(4'h8)];
                    end
                  else
                    begin
                      reg3034 <= (|reg3011);
                      reg3035 <= ((((reg2731 & reg2918) ?
                              $unsigned(reg2966) : (^(8'haf))) ^~ reg2940) ?
                          ($signed((reg1224 ?
                              reg2801 : reg2852)) << $unsigned((+reg2738))) : (+$unsigned(reg2787)));
                      reg3036 <= reg3010[(3'h4):(1'h1)];
                    end
                  if ($signed($signed((^(~&reg2727)))))
                    begin
                      reg3037 <= reg2851;
                    end
                  else
                    begin
                      reg3037 <= reg3046;
                      reg3038 <= reg2838[(3'h5):(2'h2)];
                      reg3039 <= reg2740;
                      reg3040 <= ({{$unsigned(reg3006)}} ?
                          (((reg2722 << reg2829) ?
                                  (reg2935 ? reg2870 : reg2823) : (reg2750 ?
                                      reg2750 : reg2716)) ?
                              $signed(reg1224[(3'h6):(3'h4)]) : reg2830) : reg2963);
                    end
                  if ($unsigned($unsigned({$signed(reg2921)})))
                    begin
                      reg3041 <= {$unsigned((reg2714 - (reg2853 ?
                              reg2963 : reg2919)))};
                    end
                  else
                    begin
                      reg3041 <= {((reg2800[(4'h9):(3'h5)] ?
                                  (reg2722 >= reg1205) : (^~reg2893)) ?
                              ($unsigned(reg2825) ?
                                  (reg2864 || reg2746) : (~|reg3026)) : reg2891[(3'h4):(2'h3)])};
                      reg3042 <= forvar3035;
                    end
                end
              else
                begin
                  for (forvar3034 = (1'h0); (forvar3034 < (1'h1)); forvar3034 = (forvar3034 + (1'h1)))
                    begin
                      reg3035 <= reg2866;
                      reg3036 <= {($signed((^reg1227)) <= {reg2785[(1'h0):(1'h0)]})};
                      reg3037 <= $signed((^~(reg2996[(3'h5):(3'h5)] ?
                          (reg1214 ? reg2720 : forvar3034) : (reg2815 ?
                              reg3026 : reg2960))));
                      reg3038 <= (!($signed(reg2746[(2'h2):(1'h1)]) != {$signed(forvar3032)}));
                    end
                  for (forvar3039 = (1'h0); (forvar3039 < (1'h0)); forvar3039 = (forvar3039 + (1'h1)))
                    begin
                      reg3040 <= wire1193[(3'h4):(1'h1)];
                      reg3041 <= (|reg2969);
                      reg3042 <= (~&$unsigned((~^((8'had) <= reg2750))));
                      reg3043 <= (8'ha5);
                    end
                  reg3044 <= reg1203[(1'h0):(1'h0)];
                  reg3045 <= $unsigned($signed(((reg3014 ?
                      reg2867 : reg3029) <<< (reg2813 ? reg2993 : reg2799))));
                end
              for (forvar3046 = (1'h0); (forvar3046 < (1'h0)); forvar3046 = (forvar3046 + (1'h1)))
                begin
                  if ($signed($unsigned(reg2826[(2'h2):(1'h0)])))
                    begin
                      reg3047 <= (^((~reg2785) || ((reg2770 && reg2753) ?
                          (^reg2754) : (reg2937 ? reg3031 : reg2910))));
                      reg3048 <= $signed(reg3002[(2'h3):(2'h2)]);
                      reg3049 <= reg2878;
                      reg3050 <= $unsigned(((reg2814[(4'h9):(4'h9)] <<< reg2922) ^~ ($unsigned((8'hb0)) && (reg2828 ?
                          reg2822 : forvar3039))));
                    end
                  else
                    begin
                      reg3047 <= reg2825[(4'h9):(3'h6)];
                      reg3048 <= $signed(($unsigned($signed((8'hab))) ?
                          reg2807[(2'h2):(2'h2)] : reg2998[(4'hc):(4'hb)]));
                    end
                end
            end
          else
            begin
              reg3034 <= (!((~^$unsigned(reg1216)) & (reg2772[(2'h2):(1'h0)] > $signed(reg2916))));
            end
        end
      if ({$signed(reg2769)})
        begin
          if ((8'ha9))
            begin
              for (forvar3051 = (1'h0); (forvar3051 < (2'h2)); forvar3051 = (forvar3051 + (1'h1)))
                begin
                  if ($unsigned({($signed(reg2958) || $unsigned(reg2722))}))
                    begin
                      reg3052 <= $signed(reg2895[(2'h2):(1'h0)]);
                      reg3053 <= wire1191;
                    end
                  else
                    begin
                      reg3052 <= ({((forvar3023 ?
                              reg2871 : reg2846) > (reg3043 ~^ (8'hb5)))} * {$signed($signed((8'ha1)))});
                    end
                  if (($signed($signed(reg2718)) ~^ (8'ha8)))
                    begin
                      reg3054 <= reg3015;
                    end
                  else
                    begin
                      reg3054 <= reg2987;
                      reg3055 <= (8'hb4);
                      reg3056 <= $signed({((~&reg2723) ?
                              $unsigned(reg2936) : $unsigned(reg2897))});
                      reg3057 <= $signed(reg2883[(3'h5):(1'h0)]);
                    end
                  for (forvar3058 = (1'h0); (forvar3058 < (2'h3)); forvar3058 = (forvar3058 + (1'h1)))
                    begin
                      reg3059 <= ((($unsigned(reg1229) ?
                                  (reg3038 ?
                                      reg2883 : reg2961) : reg2958[(4'hc):(4'hb)]) ?
                              reg1222 : $signed({(8'haf)})) ?
                          $unsigned($unsigned(reg2877)) : (($signed(reg2865) ^~ $signed(reg2754)) ?
                              $unsigned({reg2921}) : (~&(wire1192 ?
                                  reg2739 : reg2901))));
                      reg3060 <= (~|((~^{reg3042}) ?
                          (~reg2842[(1'h0):(1'h0)]) : $unsigned((+reg2781))));
                    end
                end
              reg3061 <= $signed(reg2993[(4'he):(2'h3)]);
              if ($signed((((~^reg2827) ? {reg3033} : $unsigned(forvar3032)) ?
                  (8'ha5) : ({reg2928} ?
                      (wire1191 ^~ reg2723) : $unsigned(reg1229)))))
                begin
                  for (forvar3062 = (1'h0); (forvar3062 < (1'h1)); forvar3062 = (forvar3062 + (1'h1)))
                    begin
                      reg3063 <= {((-(reg2920 ? reg2723 : (8'hae))) ?
                              $unsigned($signed(reg2987)) : forvar3058)};
                      reg3064 <= (reg1239 ?
                          (+reg1237[(3'h6):(3'h6)]) : $signed((8'ha1)));
                    end
                  if ((reg2717 ? (^~$signed((!reg2710))) : reg2924))
                    begin
                      reg3065 <= ($unsigned(reg3042) ?
                          reg2980[(3'h7):(3'h7)] : $signed(((~&(8'ha2)) ?
                              $unsigned(reg3007) : reg2817[(1'h0):(1'h0)])));
                      reg3066 <= (reg2906 ~^ reg3029);
                      reg3067 <= (reg3045[(4'h8):(2'h2)] ~^ $unsigned($signed((reg2791 ~^ reg1197))));
                      reg3068 <= reg2815;
                    end
                  else
                    begin
                      reg3065 <= $unsigned((reg2738 + $signed(forvar3058)));
                    end
                  for (forvar3069 = (1'h0); (forvar3069 < (1'h0)); forvar3069 = (forvar3069 + (1'h1)))
                    begin
                      reg3070 <= ((($unsigned(reg2777) ?
                                  {reg2808} : (!reg2955)) ?
                              $signed((forvar3046 ?
                                  reg2765 : reg2996)) : $unsigned((reg3054 | reg2849))) ?
                          reg3063[(1'h0):(1'h0)] : $unsigned(reg2870[(3'h7):(3'h7)]));
                    end
                  for (forvar3071 = (1'h0); (forvar3071 < (2'h3)); forvar3071 = (forvar3071 + (1'h1)))
                    begin
                      reg3072 <= (($signed((reg2803 ^~ reg2712)) >> ($signed(reg1227) ?
                          $signed(reg2742) : $signed(reg2770))) | forvar3058);
                      reg3073 <= reg3015[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar3062 = (1'h0); (forvar3062 < (2'h2)); forvar3062 = (forvar3062 + (1'h1)))
                    begin
                      reg3063 <= $signed(($signed($signed(reg2856)) ?
                          ((reg2817 ?
                              reg3056 : (8'had)) < $signed(reg2769)) : {reg2970[(3'h7):(2'h3)]}));
                    end
                  if (($signed((^(~reg2960))) ?
                      $signed((&reg3012)) : reg3019[(4'he):(4'he)]))
                    begin
                      reg3064 <= (^~(~^(8'hb4)));
                      reg3065 <= reg2810[(1'h0):(1'h0)];
                      reg3066 <= forvar3024;
                      reg3067 <= (|reg3046);
                    end
                  else
                    begin
                      reg3064 <= $unsigned($unsigned($unsigned(reg2733[(2'h3):(2'h2)])));
                      reg3065 <= reg3020;
                      reg3066 <= reg1233;
                      reg3067 <= reg3045;
                    end
                  for (forvar3068 = (1'h0); (forvar3068 < (1'h1)); forvar3068 = (forvar3068 + (1'h1)))
                    begin
                      reg3069 <= {(8'haf)};
                    end
                  for (forvar3070 = (1'h0); (forvar3070 < (2'h2)); forvar3070 = (forvar3070 + (1'h1)))
                    begin
                      reg3071 <= reg2889[(1'h1):(1'h0)];
                      reg3072 <= reg3011;
                      reg3073 <= (-reg2817);
                    end
                end
            end
          else
            begin
              reg3051 <= (~&($unsigned((reg2927 ?
                  (8'hb8) : reg2723)) == reg2999));
              for (forvar3052 = (1'h0); (forvar3052 < (2'h2)); forvar3052 = (forvar3052 + (1'h1)))
                begin
                  reg3053 <= $signed((8'ha8));
                  if ((reg3004 & {((reg2760 ~^ reg3040) ?
                          reg2929[(3'h6):(3'h5)] : $signed(reg2991))}))
                    begin
                      reg3054 <= reg2799[(4'h8):(3'h5)];
                      reg3055 <= forvar3036[(4'ha):(4'h8)];
                      reg3056 <= reg2801;
                      reg3057 <= (reg1203 | $signed((+reg2734[(2'h3):(2'h3)])));
                    end
                  else
                    begin
                      reg3054 <= (!$signed(reg2823[(5'h10):(1'h1)]));
                      reg3055 <= (($signed((^reg3039)) || $unsigned(reg3059[(1'h0):(1'h0)])) ?
                          $signed(reg2889) : ($signed((!reg2734)) < $unsigned((forvar3052 != (8'ha1)))));
                      reg3056 <= (reg2986[(3'h7):(3'h6)] ?
                          {reg2791[(3'h6):(2'h2)]} : reg2889);
                    end
                  for (forvar3058 = (1'h0); (forvar3058 < (2'h3)); forvar3058 = (forvar3058 + (1'h1)))
                    begin
                      reg3059 <= reg1198[(4'hc):(2'h3)];
                    end
                  for (forvar3060 = (1'h0); (forvar3060 < (2'h3)); forvar3060 = (forvar3060 + (1'h1)))
                    begin
                      reg3061 <= ((!reg2785) >= (reg2970[(2'h3):(2'h3)] ?
                          ((reg2963 ^~ reg1220) != ((8'hb3) | reg2714)) : (~^$signed((8'haf)))));
                    end
                end
              for (forvar3062 = (1'h0); (forvar3062 < (2'h2)); forvar3062 = (forvar3062 + (1'h1)))
                begin
                  if ($unsigned($signed({{reg2845}})))
                    begin
                      reg3063 <= reg2850;
                      reg3064 <= ((~^($unsigned(reg2954) >>> (reg2842 ?
                          reg2963 : reg3073))) ^ (~&($unsigned(reg2775) ?
                          (reg2974 ^ reg1230) : (-forvar3025))));
                      reg3065 <= reg2900[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg3063 <= (~|reg1240[(1'h1):(1'h0)]);
                      reg3064 <= ((~&$signed(((8'ha5) ? reg2934 : (8'hb5)))) ?
                          ($signed((reg3063 < wire2837)) ?
                              ((8'ha8) && $unsigned(reg2739)) : ({(8'h9c)} != {reg3035})) : reg2863);
                      reg3065 <= (~&($signed((reg2968 ?
                          reg1226 : reg2768)) << (&(reg2895 << (8'hb7)))));
                    end
                  for (forvar3066 = (1'h0); (forvar3066 < (2'h2)); forvar3066 = (forvar3066 + (1'h1)))
                    begin
                      reg3067 <= forvar3032[(4'hb):(4'hb)];
                      reg3068 <= ((wire1191[(3'h5):(2'h3)] ^~ {(reg2985 + reg3025)}) ?
                          {reg2895} : (forvar3060[(2'h2):(1'h1)] << (reg2938 ?
                              reg2716 : $unsigned(reg3001))));
                      reg3069 <= {($signed($signed(reg2821)) ?
                              (~(|reg3008)) : reg2972)};
                      reg3070 <= $unsigned(reg3059);
                    end
                end
              if ((8'haa))
                begin
                  reg3071 <= $unsigned(reg3044);
                  for (forvar3072 = (1'h0); (forvar3072 < (1'h0)); forvar3072 = (forvar3072 + (1'h1)))
                    begin
                      reg3073 <= $signed($unsigned(((reg2793 >= reg2908) ?
                          reg2824 : $unsigned(reg2983))));
                      reg3074 <= $unsigned($unsigned(reg2967));
                      reg3075 <= (!(+$unsigned((-reg3074))));
                    end
                  reg3076 <= (reg2888[(1'h1):(1'h0)] > ($unsigned({(8'haa)}) ?
                      $signed($signed(reg2755)) : ($signed(reg2729) ?
                          $signed(reg2971) : (!reg1237))));
                end
              else
                begin
                  reg3071 <= (reg3006 ?
                      ((^~(reg2762 ? reg2851 : reg2947)) ?
                          $unsigned(((8'hba) != reg2880)) : (^reg3044)) : (^(~^{reg2860})));
                end
            end
          if (reg3050[(4'h8):(4'h8)])
            begin
              for (forvar3077 = (1'h0); (forvar3077 < (2'h3)); forvar3077 = (forvar3077 + (1'h1)))
                begin
                  if (reg2922[(4'h8):(2'h3)])
                    begin
                      reg3078 <= $unsigned(reg2928[(4'hb):(3'h6)]);
                      reg3079 <= (((8'hba) <<< ((reg2808 ?
                          reg2852 : forvar3039) == $signed(reg1200))) << reg2954);
                    end
                  else
                    begin
                      reg3078 <= $signed((!$signed($signed(reg2969))));
                      reg3079 <= (reg2868[(1'h1):(1'h1)] ?
                          reg3047[(4'hc):(3'h7)] : ($unsigned($unsigned(reg2936)) ?
                              (^(reg3051 >= reg2777)) : {forvar3028[(4'h8):(1'h0)]}));
                      reg3080 <= reg2729;
                      reg3081 <= $signed(forvar3025);
                    end
                end
              for (forvar3082 = (1'h0); (forvar3082 < (1'h1)); forvar3082 = (forvar3082 + (1'h1)))
                begin
                  for (forvar3083 = (1'h0); (forvar3083 < (1'h0)); forvar3083 = (forvar3083 + (1'h1)))
                    begin
                      reg3084 <= reg2955;
                    end
                end
            end
          else
            begin
              for (forvar3077 = (1'h0); (forvar3077 < (1'h1)); forvar3077 = (forvar3077 + (1'h1)))
                begin
                  for (forvar3078 = (1'h0); (forvar3078 < (1'h1)); forvar3078 = (forvar3078 + (1'h1)))
                    begin
                      reg3079 <= $unsigned($unsigned(((&reg2850) + $unsigned(reg2994))));
                      reg3080 <= reg2999;
                    end
                end
              for (forvar3081 = (1'h0); (forvar3081 < (1'h1)); forvar3081 = (forvar3081 + (1'h1)))
                begin
                  if ($signed((reg2848[(4'h8):(1'h0)] ?
                      $signed(forvar3083[(1'h1):(1'h1)]) : (reg1208[(4'ha):(4'ha)] && $unsigned(reg2946)))))
                    begin
                      reg3082 <= ((~|$signed({reg2723})) ?
                          (|$unsigned((~&reg2826))) : reg2714[(3'h4):(3'h4)]);
                      reg3083 <= (((reg3029[(1'h1):(1'h1)] ?
                          (-(8'h9e)) : (reg2920 ?
                              reg3043 : (8'ha7))) > $signed({reg2714})) | ({$unsigned((8'h9f))} ^ ({(8'hac)} ?
                          (reg3072 >= (8'hac)) : $signed(forvar3025))));
                      reg3084 <= reg3006;
                    end
                  else
                    begin
                      reg3082 <= (~&(8'haa));
                      reg3083 <= ($unsigned($signed($unsigned(reg2788))) ?
                          (!reg2803) : (|((reg3073 == reg2788) ?
                              reg2779 : (^~(8'hb6)))));
                      reg3084 <= reg2828;
                      reg3085 <= reg3011;
                    end
                  if ((+($unsigned((reg1205 + reg2905)) <<< (((8'ha1) ^ reg3007) << reg2970))))
                    begin
                      reg3086 <= (((8'ha1) ?
                          ({(8'ha1)} * $unsigned(reg2964)) : reg2975) != $unsigned(reg2897));
                      reg3087 <= $signed($signed((~|(reg2924 ?
                          reg2738 : (8'ha5)))));
                      reg3088 <= $signed((($unsigned(forvar3072) ?
                          (~^forvar3035) : (&reg3082)) | (reg1205 != $signed(reg3016))));
                      reg3089 <= {$signed(forvar3077[(5'h10):(4'hc)])};
                    end
                  else
                    begin
                      reg3086 <= {reg3080[(2'h3):(1'h1)]};
                    end
                  for (forvar3090 = (1'h0); (forvar3090 < (2'h2)); forvar3090 = (forvar3090 + (1'h1)))
                    begin
                      reg3091 <= (reg2852 + $signed(reg3074[(3'h5):(3'h4)]));
                      reg3092 <= $unsigned((8'ha1));
                      reg3093 <= ((|(+(~|reg3074))) ?
                          {$unsigned($signed(reg2818))} : ((-((8'hb2) || wire1191)) && ((reg2786 < (8'ha2)) ?
                              (reg2781 | reg2735) : (reg2989 | reg2833))));
                    end
                  if ($unsigned((reg2987[(2'h2):(1'h0)] > $unsigned($signed(reg3000)))))
                    begin
                      reg3094 <= $signed(($unsigned(((8'hae) | reg2919)) ?
                          ((~&reg2724) ?
                              $unsigned(reg2817) : (reg2787 ?
                                  reg3004 : reg2966)) : $unsigned($signed(reg3026))));
                      reg3095 <= $signed($unsigned($signed(((8'ha1) ?
                          reg3032 : reg3012))));
                      reg3096 <= $signed(reg2787);
                    end
                  else
                    begin
                      reg3094 <= $unsigned($signed(forvar3082[(1'h1):(1'h1)]));
                      reg3095 <= $signed((reg2717 <<< reg3006));
                      reg3096 <= reg2958[(4'h9):(4'h8)];
                    end
                end
              for (forvar3097 = (1'h0); (forvar3097 < (1'h0)); forvar3097 = (forvar3097 + (1'h1)))
                begin
                  reg3098 <= $signed((+($unsigned(reg3039) ?
                      $signed(reg2908) : {reg3034})));
                end
            end
          reg3099 <= reg2803;
          for (forvar3100 = (1'h0); (forvar3100 < (2'h3)); forvar3100 = (forvar3100 + (1'h1)))
            begin
              for (forvar3101 = (1'h0); (forvar3101 < (2'h3)); forvar3101 = (forvar3101 + (1'h1)))
                begin
                  for (forvar3102 = (1'h0); (forvar3102 < (1'h1)); forvar3102 = (forvar3102 + (1'h1)))
                    begin
                      reg3103 <= reg2988[(1'h0):(1'h0)];
                      reg3104 <= (^~reg2780);
                    end
                  for (forvar3105 = (1'h0); (forvar3105 < (2'h3)); forvar3105 = (forvar3105 + (1'h1)))
                    begin
                      reg3106 <= (!reg2751[(3'h4):(1'h0)]);
                      reg3107 <= ((8'hb5) ?
                          (reg2753 ?
                              (!reg2807) : reg2955[(4'h8):(3'h7)]) : reg2829);
                    end
                  if (reg3049[(3'h5):(3'h4)])
                    begin
                      reg3108 <= ((!$unsigned((reg3025 ^ reg2777))) ?
                          $unsigned((reg3042[(2'h3):(1'h0)] ?
                              (+reg2956) : reg3084)) : reg2869[(2'h3):(1'h0)]);
                      reg3109 <= ((((reg2973 ?
                              reg3059 : reg1216) << {reg3036}) != reg2772) ?
                          ($signed($signed(reg2870)) ?
                              $signed((reg2800 * (8'haf))) : (8'h9f)) : ((8'ha8) ^~ {{(8'ha0)}}));
                      reg3110 <= forvar3101[(2'h3):(2'h2)];
                      reg3111 <= (|$signed(((reg2896 || wire1188) ?
                          (forvar3071 && (8'hae)) : (reg2715 ?
                              reg2926 : reg3027))));
                    end
                  else
                    begin
                      reg3108 <= $signed(((~^reg2728[(2'h3):(2'h2)]) <<< reg2833));
                    end
                end
              if ($signed(({reg2732[(3'h4):(2'h2)]} ^ (-reg1220))))
                begin
                  if ($unsigned($signed({reg2954})))
                    begin
                      reg3112 <= ($unsigned(reg2931) - $signed($unsigned((8'ha7))));
                      reg3113 <= (~^reg2919);
                    end
                  else
                    begin
                      reg3112 <= ($unsigned((~&$signed(forvar3023))) & {$signed($unsigned(reg2967))});
                      reg3113 <= (reg2721[(2'h3):(1'h1)] ?
                          (~|{(reg3049 ?
                                  reg2957 : reg2731)}) : $unsigned($unsigned((reg3047 < reg2849))));
                      reg3114 <= {($signed((|forvar3062)) ?
                              ((reg2779 <<< forvar3036) ?
                                  $signed(reg2840) : reg2759[(4'hc):(3'h5)]) : reg2910)};
                      reg3115 <= ($unsigned($signed((|reg3038))) * reg2999[(2'h3):(2'h2)]);
                    end
                  reg3116 <= (reg3078[(1'h0):(1'h0)] || {forvar3102[(2'h2):(1'h1)]});
                end
              else
                begin
                  if ((($unsigned((!reg2790)) ?
                          (!reg3023[(4'ha):(2'h2)]) : reg2936) ?
                      reg2971[(3'h5):(2'h3)] : (reg2747 | $signed($signed((8'ha8))))))
                    begin
                      reg3112 <= (8'hab);
                      reg3113 <= (~|((-$signed(reg3033)) ?
                          $signed((reg2995 ?
                              reg3096 : forvar3070)) : $unsigned($unsigned(reg2919))));
                    end
                  else
                    begin
                      reg3112 <= reg3012;
                    end
                  if ({reg2861})
                    begin
                      reg3114 <= reg2985[(1'h0):(1'h0)];
                      reg3115 <= ($unsigned({(reg2962 ? reg3005 : reg2746)}) ?
                          $signed((~&(reg2740 & reg3044))) : $unsigned({reg2904[(1'h0):(1'h0)]}));
                      reg3116 <= (~&$unsigned($signed((reg2934 - (8'h9d)))));
                    end
                  else
                    begin
                      reg3114 <= $unsigned($unsigned($signed($signed(reg3061))));
                      reg3115 <= reg2975[(4'ha):(2'h2)];
                    end
                end
              for (forvar3117 = (1'h0); (forvar3117 < (1'h0)); forvar3117 = (forvar3117 + (1'h1)))
                begin
                  for (forvar3118 = (1'h0); (forvar3118 < (2'h3)); forvar3118 = (forvar3118 + (1'h1)))
                    begin
                      reg3119 <= $signed((+reg3043));
                      reg3120 <= (reg2873[(2'h2):(2'h2)] * (($signed(reg2744) ?
                              (-reg3112) : (reg2721 ? reg2813 : (8'h9c))) ?
                          $signed((reg2879 ?
                              reg2913 : (8'had))) : $signed($signed(reg1215))));
                      reg3121 <= {(((~^reg2880) ?
                                  (forvar3038 ?
                                      reg2998 : (8'ha3)) : $signed(reg2866)) ?
                              ((reg2844 ~^ reg2852) ?
                                  (reg3069 && reg2945) : reg2818) : $signed((reg3093 ?
                                  reg2913 : reg3042)))};
                    end
                  for (forvar3122 = (1'h0); (forvar3122 < (2'h3)); forvar3122 = (forvar3122 + (1'h1)))
                    begin
                      reg3123 <= $unsigned($unsigned(($signed(reg3023) ?
                          (wire1193 == reg2732) : reg2710)));
                      reg3124 <= $signed(((^$unsigned((8'hb1))) ?
                          ($unsigned(reg1213) ?
                              (~reg2738) : reg2819[(3'h7):(3'h4)]) : reg1228[(2'h2):(1'h1)]));
                      reg3125 <= $unsigned((reg2924[(2'h2):(1'h1)] ?
                          reg1229[(3'h4):(2'h3)] : $signed(reg2834[(3'h4):(1'h1)])));
                    end
                  if (reg2763[(1'h1):(1'h1)])
                    begin
                      reg3126 <= reg2899[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg3126 <= $signed(reg2857);
                      reg3127 <= (-reg2834);
                      reg3128 <= reg1216[(2'h2):(1'h1)];
                      reg3129 <= $unsigned({(~|$signed((8'hb7)))});
                    end
                  if ((^$signed($signed(((8'hb7) ? reg1205 : (8'hb5))))))
                    begin
                      reg3130 <= (~|($signed((^~reg2760)) ?
                          $signed($signed(forvar3072)) : (reg2897[(1'h1):(1'h1)] ?
                              reg1235 : (~(8'ha8)))));
                      reg3131 <= (&($signed(reg2997[(3'h7):(3'h5)]) * reg2831[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg3130 <= $signed($unsigned($signed(reg3086)));
                      reg3131 <= $unsigned(reg3045);
                      reg3132 <= (($unsigned($unsigned(reg2869)) ^ ((reg2770 >= reg1222) ?
                          $signed(reg2911) : $unsigned(reg2937))) ^~ reg2847);
                    end
                end
            end
        end
      else
        begin
          for (forvar3051 = (1'h0); (forvar3051 < (1'h0)); forvar3051 = (forvar3051 + (1'h1)))
            begin
              if (reg2965)
                begin
                  for (forvar3052 = (1'h0); (forvar3052 < (1'h0)); forvar3052 = (forvar3052 + (1'h1)))
                    begin
                      reg3053 <= (^~(+$unsigned((reg2899 ?
                          reg2713 : forvar3072))));
                      reg3054 <= (^~reg2709);
                      reg3055 <= (reg3113[(2'h3):(1'h1)] ?
                          reg1234 : $signed($unsigned($signed(reg3020))));
                      reg3056 <= (+$unsigned($signed((forvar3097 > reg2920))));
                    end
                  if ((|(reg2984 ?
                      reg2949[(1'h1):(1'h1)] : reg2791[(4'hd):(4'h8)])))
                    begin
                      reg3057 <= $signed($signed(((|reg3066) >= ((8'ha9) ?
                          reg2764 : (8'hb7)))));
                    end
                  else
                    begin
                      reg3057 <= ((reg2765 ?
                          {$unsigned(reg2735)} : (reg2821[(1'h1):(1'h0)] ?
                              (8'haa) : $unsigned(reg2879))) != reg2920);
                    end
                  if (({(^~(~^reg2856))} << reg2786[(2'h2):(2'h2)]))
                    begin
                      reg3058 <= {$unsigned((reg2995[(4'hb):(2'h2)] - ((8'hb5) ?
                              reg3009 : reg3028)))};
                      reg3059 <= $unsigned($unsigned(($unsigned(forvar3052) * reg3051)));
                    end
                  else
                    begin
                      reg3058 <= $unsigned((((^reg3110) ?
                              reg3110[(3'h4):(1'h0)] : (~&reg1216)) ?
                          ($unsigned(reg1222) - $signed(reg3075)) : reg3006[(3'h6):(3'h6)]));
                      reg3059 <= reg1199;
                      reg3060 <= $unsigned(((~(reg2762 ?
                          reg2838 : reg1213)) << $unsigned(reg2894)));
                      reg3061 <= $unsigned((reg2857 ?
                          $signed((reg1205 ?
                              forvar3101 : reg2739)) : $signed((reg3110 <= reg3092))));
                    end
                end
              else
                begin
                  for (forvar3052 = (1'h0); (forvar3052 < (2'h3)); forvar3052 = (forvar3052 + (1'h1)))
                    begin
                      reg3053 <= $unsigned($signed(reg2759[(2'h2):(1'h0)]));
                      reg3054 <= $unsigned(reg3086);
                    end
                end
              if (reg2904)
                begin
                  if (((~|(~&$unsigned(reg2765))) ?
                      (reg2940 << $signed(reg1229)) : reg2926))
                    begin
                      reg3062 <= {(forvar3032[(3'h7):(3'h5)] << ((forvar3034 ?
                                  (8'hb3) : reg2815) ?
                              ((8'h9e) ?
                                  reg2977 : reg2961) : $signed((8'hb7))))};
                    end
                  else
                    begin
                      reg3062 <= reg2888;
                      reg3063 <= ($signed($signed({reg2968})) - (({reg3062} ?
                              forvar3069 : $unsigned(reg2958)) ?
                          (~|((8'haf) == reg3043)) : $unsigned(reg3017)));
                      reg3064 <= $signed(($unsigned((!reg2892)) || (reg3010 <<< {wire1192})));
                    end
                end
              else
                begin
                  reg3062 <= ($signed($signed(reg2972)) ?
                      $signed(($unsigned((8'ha6)) || (reg2919 ?
                          reg2996 : reg3051))) : reg2822[(1'h1):(1'h1)]);
                end
            end
          for (forvar3065 = (1'h0); (forvar3065 < (2'h3)); forvar3065 = (forvar3065 + (1'h1)))
            begin
              reg3066 <= (+{reg2923});
              for (forvar3067 = (1'h0); (forvar3067 < (1'h0)); forvar3067 = (forvar3067 + (1'h1)))
                begin
                  if ((reg2778[(1'h1):(1'h0)] ?
                      (reg3119[(4'h8):(1'h1)] << ((~&(8'h9f)) ?
                          $unsigned(reg2914) : reg2795)) : (&reg2755[(2'h2):(2'h2)])))
                    begin
                      reg3068 <= ((reg2827[(1'h1):(1'h1)] | ($unsigned(reg2997) ?
                          $signed(reg3058) : {reg2906})) >> $unsigned({((8'had) ?
                              (8'ha4) : reg2807)}));
                    end
                  else
                    begin
                      reg3068 <= $unsigned({(|$signed(reg2859))});
                    end
                  for (forvar3069 = (1'h0); (forvar3069 < (1'h0)); forvar3069 = (forvar3069 + (1'h1)))
                    begin
                      reg3070 <= reg2917[(2'h2):(1'h0)];
                      reg3071 <= (((reg3088 > reg3103[(1'h1):(1'h1)]) - (reg1209 == (reg2991 ?
                          forvar3071 : reg3123))) ^ $unsigned((|(&reg2984))));
                      reg3072 <= $signed(reg2802[(2'h3):(1'h0)]);
                      reg3073 <= (+(reg2998 ^~ $unsigned($unsigned(reg1230))));
                    end
                  if (($unsigned(((^reg2842) <<< {reg2848})) ?
                      {reg2895[(2'h2):(1'h1)]} : (8'h9e)))
                    begin
                      reg3074 <= (($signed($signed(reg2994)) == reg3071) ?
                          $unsigned($signed(reg2710)) : {$signed((reg3049 ?
                                  reg2869 : reg2869))});
                      reg3075 <= {((^reg3119[(3'h4):(1'h0)]) ?
                              (+$unsigned((8'hae))) : {(~&reg1235)})};
                    end
                  else
                    begin
                      reg3074 <= $signed($unsigned({reg2936}));
                      reg3075 <= (|reg2873[(4'hf):(4'he)]);
                    end
                end
            end
          for (forvar3076 = (1'h0); (forvar3076 < (2'h2)); forvar3076 = (forvar3076 + (1'h1)))
            begin
              if ((~$signed((~|reg2950))))
                begin
                  for (forvar3077 = (1'h0); (forvar3077 < (2'h3)); forvar3077 = (forvar3077 + (1'h1)))
                    begin
                      reg3078 <= $signed(reg3016);
                      reg3079 <= forvar3023[(4'hc):(3'h6)];
                      reg3080 <= reg2810;
                      reg3081 <= reg2909[(5'h10):(3'h6)];
                    end
                  for (forvar3082 = (1'h0); (forvar3082 < (1'h0)); forvar3082 = (forvar3082 + (1'h1)))
                    begin
                      reg3083 <= {{$signed(reg3029[(2'h3):(1'h1)])}};
                    end
                  if ((8'ha6))
                    begin
                      reg3084 <= ({$unsigned({reg3083})} ?
                          reg3022[(1'h1):(1'h1)] : $unsigned(((~reg3113) ?
                              $signed(reg2879) : reg2977[(4'h8):(3'h5)])));
                      reg3085 <= (&((((8'ha8) ?
                              reg2796 : reg2765) == $unsigned(forvar3118)) ?
                          ($unsigned(reg3060) << (reg2984 ?
                              reg3044 : reg2994)) : (^(reg2930 ^ reg2813))));
                    end
                  else
                    begin
                      reg3084 <= (~&$signed($unsigned($signed(reg2961))));
                    end
                end
              else
                begin
                  for (forvar3077 = (1'h0); (forvar3077 < (1'h1)); forvar3077 = (forvar3077 + (1'h1)))
                    begin
                      reg3078 <= {$unsigned($unsigned($unsigned(reg2739)))};
                    end
                  for (forvar3079 = (1'h0); (forvar3079 < (2'h2)); forvar3079 = (forvar3079 + (1'h1)))
                    begin
                      reg3080 <= (reg2928[(4'hc):(4'hc)] >>> (&(((8'hb6) == reg2949) ?
                          (8'ha8) : $signed(reg2771))));
                      reg3081 <= (~&$signed(($signed(wire1191) ?
                          $unsigned((8'haf)) : {reg2980})));
                      reg3082 <= (reg2983 ?
                          $signed((!$unsigned(reg2725))) : reg2892[(2'h2):(1'h0)]);
                    end
                end
              reg3086 <= $unsigned($signed($signed((forvar3071 ?
                  reg3127 : reg2715))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg3133 <= {((~|wire1193) + reg2798)};
      for (forvar3134 = (1'h0); (forvar3134 < (2'h2)); forvar3134 = (forvar3134 + (1'h1)))
        begin
          for (forvar3135 = (1'h0); (forvar3135 < (1'h0)); forvar3135 = (forvar3135 + (1'h1)))
            begin
              for (forvar3136 = (1'h0); (forvar3136 < (1'h0)); forvar3136 = (forvar3136 + (1'h1)))
                begin
                  if (reg2930[(3'h4):(1'h1)])
                    begin
                      reg3137 <= ((!{(reg2768 >>> reg3132)}) ?
                          reg2958 : (!reg2766));
                      reg3138 <= $unsigned({((reg2958 ?
                              reg2917 : reg3104) << reg2725[(1'h1):(1'h1)])});
                    end
                  else
                    begin
                      reg3137 <= $unsigned(($unsigned(reg2817[(1'h0):(1'h0)]) << reg2803));
                      reg3138 <= {reg2727};
                      reg3139 <= $unsigned($signed({((8'hb7) ?
                              reg2733 : reg2998)}));
                    end
                  for (forvar3140 = (1'h0); (forvar3140 < (2'h2)); forvar3140 = (forvar3140 + (1'h1)))
                    begin
                      reg3141 <= (reg2731[(3'h6):(1'h0)] ?
                          reg2857[(3'h7):(3'h6)] : $unsigned(((reg2919 * reg2899) ?
                              $unsigned(reg3039) : (reg2826 ^ reg2712))));
                      reg3142 <= ((reg3059 ?
                          reg2930[(1'h0):(1'h0)] : reg3096[(2'h2):(1'h1)]) & (~|((reg3011 ?
                              reg1199 : reg2919) ?
                          reg2988[(2'h3):(2'h2)] : reg2985)));
                    end
                  reg3143 <= ($signed((!(reg2845 ? reg3060 : (8'ha0)))) ?
                      ($unsigned(reg2888) ?
                          $unsigned({(8'hab)}) : $unsigned(reg2980[(4'h8):(1'h1)])) : reg2907[(3'h6):(1'h1)]);
                end
              reg3144 <= (reg2915 < $signed((reg2826[(1'h1):(1'h0)] != (&reg2724))));
            end
        end
      for (forvar3145 = (1'h0); (forvar3145 < (2'h3)); forvar3145 = (forvar3145 + (1'h1)))
        begin
          for (forvar3146 = (1'h0); (forvar3146 < (2'h2)); forvar3146 = (forvar3146 + (1'h1)))
            begin
              for (forvar3147 = (1'h0); (forvar3147 < (2'h3)); forvar3147 = (forvar3147 + (1'h1)))
                begin
                  for (forvar3148 = (1'h0); (forvar3148 < (2'h3)); forvar3148 = (forvar3148 + (1'h1)))
                    begin
                      reg3149 <= ((reg3062[(1'h0):(1'h0)] < $unsigned($signed(wire1241))) * $signed(($unsigned((8'hb5)) ?
                          reg2762 : {reg2777})));
                      reg3150 <= $unsigned((^~reg3095));
                      reg3151 <= $unsigned(reg2726[(1'h1):(1'h0)]);
                    end
                end
              for (forvar3152 = (1'h0); (forvar3152 < (1'h0)); forvar3152 = (forvar3152 + (1'h1)))
                begin
                  if ((reg1239[(4'hc):(3'h5)] ? reg2853 : $signed((^reg2970))))
                    begin
                      reg3153 <= ($signed($signed($signed(reg3144))) & (-{$unsigned(reg2904)}));
                      reg3154 <= (($signed((reg2763 ? (8'hb2) : (8'ha8))) ?
                              (~|reg2737[(3'h7):(3'h4)]) : $signed((reg2732 ^ reg3123))) ?
                          (8'ha8) : (-((reg3040 < (8'hb9)) && reg2883[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg3153 <= ($unsigned(($unsigned(reg2908) & reg2859[(2'h2):(1'h0)])) >>> $signed(($signed(reg2962) ?
                          (reg3001 > reg2708) : $unsigned((8'h9c)))));
                      reg3154 <= reg3150[(4'hb):(3'h5)];
                      reg3155 <= (8'ha5);
                      reg3156 <= reg3051;
                    end
                end
              reg3157 <= reg2831[(1'h1):(1'h1)];
            end
          for (forvar3158 = (1'h0); (forvar3158 < (1'h1)); forvar3158 = (forvar3158 + (1'h1)))
            begin
              reg3159 <= (~|reg3058[(3'h6):(3'h6)]);
              for (forvar3160 = (1'h0); (forvar3160 < (1'h1)); forvar3160 = (forvar3160 + (1'h1)))
                begin
                  if ($unsigned(reg2967))
                    begin
                      reg3161 <= $signed(($signed($signed(reg2806)) ?
                          (reg2769 + $signed(reg2742)) : (^~$signed(reg3074))));
                      reg3162 <= reg2807[(2'h2):(2'h2)];
                      reg3163 <= (8'hac);
                      reg3164 <= {(((reg3156 * reg2847) == $signed(reg2784)) ?
                              ((~|reg2931) ^~ reg2710[(2'h2):(1'h0)]) : reg3050[(2'h2):(1'h0)])};
                    end
                  else
                    begin
                      reg3161 <= {$signed(reg3073[(1'h1):(1'h0)])};
                    end
                  if ((~$unsigned($signed((reg2749 == reg2732)))))
                    begin
                      reg3165 <= $signed(reg2892[(3'h5):(1'h1)]);
                      reg3166 <= reg3113;
                      reg3167 <= ((~^((reg2840 ? (8'ha1) : reg3026) ?
                          (|reg2740) : $unsigned(reg3111))) != ($signed($signed(reg2849)) * $unsigned((reg2914 >> (8'haf)))));
                      reg3168 <= $signed({(^~(|(8'had)))});
                    end
                  else
                    begin
                      reg3165 <= reg3164[(4'h8):(2'h2)];
                    end
                end
            end
        end
      for (forvar3169 = (1'h0); (forvar3169 < (2'h2)); forvar3169 = (forvar3169 + (1'h1)))
        begin
          if ($unsigned(reg2715))
            begin
              reg3170 <= reg2806[(1'h0):(1'h0)];
            end
          else
            begin
              for (forvar3170 = (1'h0); (forvar3170 < (2'h3)); forvar3170 = (forvar3170 + (1'h1)))
                begin
                  reg3171 <= reg3082;
                  reg3172 <= reg2780[(1'h1):(1'h1)];
                  for (forvar3173 = (1'h0); (forvar3173 < (2'h2)); forvar3173 = (forvar3173 + (1'h1)))
                    begin
                      reg3174 <= {$signed(((reg3127 ? reg2766 : (8'ha4)) ?
                              reg2780[(1'h1):(1'h0)] : (8'h9c)))};
                      reg3175 <= ((+((reg2962 ? reg2778 : reg3088) ?
                              {(8'hb0)} : reg3058)) ?
                          reg3020[(2'h3):(1'h1)] : ($unsigned((reg1198 >= (8'hb0))) ?
                              reg2806 : reg3071));
                      reg3176 <= reg2902;
                    end
                  reg3177 <= (!reg2902);
                end
            end
          for (forvar3178 = (1'h0); (forvar3178 < (1'h0)); forvar3178 = (forvar3178 + (1'h1)))
            begin
              for (forvar3179 = (1'h0); (forvar3179 < (2'h3)); forvar3179 = (forvar3179 + (1'h1)))
                begin
                  if (({(^(8'ha0))} ~^ {{(reg2999 - reg3076)}}))
                    begin
                      reg3180 <= ($signed((reg2802[(1'h1):(1'h1)] ?
                          (reg3159 ?
                              reg3151 : (8'haf)) : $unsigned(reg2843))) > reg3025);
                    end
                  else
                    begin
                      reg3180 <= {({reg2842[(1'h0):(1'h0)]} >>> $unsigned(reg2940[(3'h6):(3'h6)]))};
                      reg3181 <= reg3049;
                      reg3182 <= $signed(reg3165[(1'h1):(1'h0)]);
                    end
                  if ($signed($signed((&$unsigned(reg3170)))))
                    begin
                      reg3183 <= (&reg3080[(1'h0):(1'h0)]);
                      reg3184 <= {(!reg2986)};
                      reg3185 <= ($unsigned({(~&reg2899)}) ?
                          (((reg2709 != (8'haf)) ^~ (^~reg3073)) && $unsigned(reg3085)) : $unsigned(($unsigned(reg2800) >>> (reg2846 ?
                              reg2716 : (8'ha5)))));
                      reg3186 <= ($unsigned((~|{reg1235})) <<< reg3068);
                    end
                  else
                    begin
                      reg3183 <= ((!$signed($unsigned(reg2963))) == reg3082[(1'h0):(1'h0)]);
                    end
                  if ((($signed($signed(reg2709)) <<< $signed(reg1217[(4'h8):(3'h7)])) ?
                      ((^~(~&reg2950)) | reg2992[(3'h6):(2'h3)]) : reg1202))
                    begin
                      reg3187 <= $unsigned((~(((8'ha6) ?
                          (8'hb3) : reg2958) << reg3126)));
                      reg3188 <= $unsigned($signed($signed($unsigned(reg2910))));
                      reg3189 <= reg2712;
                      reg3190 <= reg2961[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3187 <= {(^reg1213)};
                      reg3188 <= $unsigned(reg3172[(4'ha):(4'h8)]);
                      reg3189 <= (~^reg1202);
                    end
                end
              reg3191 <= wire1241[(2'h2):(1'h0)];
            end
          if ($signed(reg3177))
            begin
              reg3192 <= reg2866[(4'h9):(4'h8)];
              if ({reg3143})
                begin
                  if ((reg2752 ? reg2797 : $unsigned($signed({reg3096}))))
                    begin
                      reg3193 <= reg2970[(3'h6):(1'h1)];
                      reg3194 <= (~&(reg2927[(1'h1):(1'h0)] || $signed((~^reg2734))));
                      reg3195 <= ($unsigned(($unsigned(reg2824) || $unsigned(reg2857))) != $signed(reg2788));
                    end
                  else
                    begin
                      reg3193 <= reg2761[(3'h4):(2'h3)];
                      reg3194 <= ((reg2905[(3'h4):(1'h1)] & reg3153) ?
                          reg2815[(3'h4):(2'h3)] : (8'hb2));
                    end
                  for (forvar3196 = (1'h0); (forvar3196 < (2'h3)); forvar3196 = (forvar3196 + (1'h1)))
                    begin
                      reg3197 <= $signed((reg2756[(3'h5):(2'h3)] != ($unsigned(reg2906) ?
                          (reg2970 + reg2771) : reg2977[(3'h6):(2'h3)])));
                    end
                  if ({$signed(reg3074[(1'h0):(1'h0)])})
                    begin
                      reg3198 <= {{(reg3156 ?
                                  $unsigned(reg3001) : reg2943[(1'h1):(1'h1)])}};
                      reg3199 <= $signed($signed(reg2708));
                      reg3200 <= reg2758[(4'h8):(4'h8)];
                      reg3201 <= $signed(reg2768[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg3198 <= (^~((reg2912 >>> (reg2918 ?
                              reg2991 : reg2843)) ?
                          $signed(reg2780[(4'h9):(1'h0)]) : $signed((reg2863 ?
                              reg3007 : reg3017))));
                      reg3199 <= reg2963;
                      reg3200 <= ($unsigned((-$signed(reg2728))) ?
                          (-((|reg3086) || reg1229)) : ($signed($signed(reg3056)) ?
                              (reg2967 > $unsigned(reg2861)) : reg3055[(1'h0):(1'h0)]));
                    end
                  for (forvar3202 = (1'h0); (forvar3202 < (1'h1)); forvar3202 = (forvar3202 + (1'h1)))
                    begin
                      reg3203 <= (reg2966[(2'h3):(2'h3)] >>> ((8'hb2) ?
                          (&wire2837) : (reg3085 >>> reg2949)));
                      reg3204 <= $unsigned((((~&reg3131) ?
                          $unsigned(reg3155) : $signed(reg2947)) && {(8'hb1)}));
                      reg3205 <= forvar3134[(2'h3):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar3193 = (1'h0); (forvar3193 < (1'h1)); forvar3193 = (forvar3193 + (1'h1)))
                    begin
                      reg3194 <= (reg3041 ?
                          (reg2775 ?
                              reg1235 : $signed((reg2970 ?
                                  reg2908 : reg2795))) : (reg3041 >= $signed($unsigned(forvar3136))));
                      reg3195 <= (8'hb6);
                    end
                  for (forvar3196 = (1'h0); (forvar3196 < (1'h0)); forvar3196 = (forvar3196 + (1'h1)))
                    begin
                      reg3197 <= forvar3147;
                      reg3198 <= $signed($signed((8'hb2)));
                      reg3199 <= ((((reg2841 ? reg3085 : reg2770) ?
                              (8'hb9) : reg2923) ?
                          (~|(8'hba)) : $unsigned($unsigned(reg2747))) != reg2942);
                      reg3200 <= (8'ha5);
                    end
                  if ($unsigned((^~((reg3078 + reg2962) >= $signed(reg2827)))))
                    begin
                      reg3201 <= ((~{reg1232}) != $unsigned(($unsigned(reg2962) ?
                          reg2970 : $unsigned(reg3006))));
                      reg3202 <= {(^~(~&reg2953[(1'h1):(1'h1)]))};
                    end
                  else
                    begin
                      reg3201 <= reg3194[(4'hf):(3'h6)];
                      reg3202 <= $signed(($unsigned((forvar3196 || reg2735)) << ((reg2807 << (8'ha3)) ?
                          $signed(reg3170) : reg2819[(3'h7):(2'h2)])));
                      reg3203 <= $signed((~{((8'hba) ? reg3112 : reg2723)}));
                      reg3204 <= (reg3115[(4'h8):(1'h1)] ?
                          $signed($signed($signed(forvar3193))) : $signed(($signed(reg2867) - $signed(reg3141))));
                    end
                  if ($signed(((8'hb1) > (~&(reg2854 ? reg2928 : (8'ha8))))))
                    begin
                      reg3205 <= ($signed((&(reg3072 ? reg2857 : reg1208))) ?
                          ((!reg3086) >>> reg2838) : ((8'hb1) <<< {forvar3136[(3'h4):(2'h3)]}));
                      reg3206 <= reg2840;
                    end
                  else
                    begin
                      reg3205 <= reg1222[(2'h3):(2'h3)];
                      reg3206 <= reg3060;
                      reg3207 <= reg2919;
                    end
                end
              if (reg2983)
                begin
                  reg3208 <= reg2780;
                  for (forvar3209 = (1'h0); (forvar3209 < (2'h2)); forvar3209 = (forvar3209 + (1'h1)))
                    begin
                      reg3210 <= reg2810;
                      reg3211 <= $unsigned({($unsigned((8'h9c)) ?
                              $signed(reg2937) : (&reg3110))});
                      reg3212 <= $signed((&$signed((reg3130 ?
                          reg3138 : (8'ha7)))));
                      reg3213 <= reg3034;
                    end
                  if ($unsigned(reg2851))
                    begin
                      reg3214 <= (~|(8'ha7));
                    end
                  else
                    begin
                      reg3214 <= (8'hae);
                      reg3215 <= reg3201;
                    end
                  if ((reg3067 ?
                      reg2969[(4'hc):(3'h4)] : {$signed(forvar3193[(4'he):(4'hc)])}))
                    begin
                      reg3216 <= $signed(reg2851[(3'h5):(2'h2)]);
                      reg3217 <= reg3063[(3'h7):(2'h3)];
                      reg3218 <= ($signed((~(forvar3136 ^~ reg2749))) > $signed($unsigned(((8'h9f) ?
                          reg1222 : (8'ha4)))));
                    end
                  else
                    begin
                      reg3216 <= (~|(&(~|reg3020[(4'h9):(3'h7)])));
                      reg3217 <= reg2970;
                      reg3218 <= reg3188;
                    end
                end
              else
                begin
                  for (forvar3208 = (1'h0); (forvar3208 < (1'h1)); forvar3208 = (forvar3208 + (1'h1)))
                    begin
                      reg3209 <= reg3011;
                    end
                  reg3210 <= ((($unsigned(reg2910) ?
                      (reg2850 ?
                          reg2817 : reg3064) : reg2829) || $unsigned(reg2719[(2'h2):(1'h1)])) <<< $unsigned($signed(reg1210[(4'hd):(4'h8)])));
                  for (forvar3211 = (1'h0); (forvar3211 < (2'h2)); forvar3211 = (forvar3211 + (1'h1)))
                    begin
                      reg3212 <= reg2954[(2'h3):(2'h2)];
                      reg3213 <= ((^~$signed(reg3143)) ?
                          (((reg3109 ?
                              (8'ha9) : reg3113) != reg2765[(4'h8):(1'h1)]) & $signed((~reg1240))) : $signed(reg2947));
                      reg3214 <= ({reg3211[(3'h7):(3'h5)]} ?
                          {($signed((8'hb7)) ?
                                  {reg2917} : $signed(reg2713))} : {$unsigned((reg3110 ?
                                  reg2951 : reg3175))});
                    end
                  reg3215 <= $signed(reg2936[(4'he):(2'h3)]);
                end
              for (forvar3219 = (1'h0); (forvar3219 < (2'h3)); forvar3219 = (forvar3219 + (1'h1)))
                begin
                  for (forvar3220 = (1'h0); (forvar3220 < (1'h0)); forvar3220 = (forvar3220 + (1'h1)))
                    begin
                      reg3221 <= {reg2972[(2'h2):(2'h2)]};
                      reg3222 <= (+($unsigned($signed(reg2921)) <<< $signed((8'ha8))));
                    end
                end
            end
          else
            begin
              for (forvar3192 = (1'h0); (forvar3192 < (2'h3)); forvar3192 = (forvar3192 + (1'h1)))
                begin
                  if (reg2969)
                    begin
                      reg3193 <= reg3035[(1'h1):(1'h0)];
                      reg3194 <= {$signed((~^reg2768[(1'h0):(1'h0)]))};
                      reg3195 <= ((&reg2760[(2'h2):(2'h2)]) ?
                          reg2827[(2'h2):(1'h0)] : (((reg2960 <<< reg3027) <<< reg2761[(3'h7):(3'h7)]) | $signed(reg2847)));
                    end
                  else
                    begin
                      reg3193 <= reg3044[(1'h1):(1'h1)];
                    end
                  for (forvar3196 = (1'h0); (forvar3196 < (2'h2)); forvar3196 = (forvar3196 + (1'h1)))
                    begin
                      reg3197 <= reg2945;
                    end
                end
              if (($signed((reg2848 ? {reg2880} : $signed(reg3014))) ?
                  ({{reg2763}} ?
                      {reg3184} : reg2716) : {($signed(reg2748) <= wire1241)}))
                begin
                  for (forvar3198 = (1'h0); (forvar3198 < (2'h3)); forvar3198 = (forvar3198 + (1'h1)))
                    begin
                      reg3199 <= (^~(^~$unsigned((reg2916 ?
                          reg3166 : reg1220))));
                      reg3200 <= (-(^~({reg3087} ?
                          forvar3192 : reg3022[(3'h5):(1'h0)])));
                      reg3201 <= reg3193;
                      reg3202 <= $signed($unsigned($unsigned(reg3057)));
                    end
                  if (reg2979[(3'h4):(2'h3)])
                    begin
                      reg3203 <= $signed((^~{reg2928[(2'h2):(2'h2)]}));
                      reg3204 <= (+$signed($unsigned($signed((8'ha4)))));
                      reg3205 <= {(~|((reg2943 ? reg2925 : reg3086) ?
                              (~|reg2733) : (reg2740 ? (8'ha2) : (8'ha4))))};
                      reg3206 <= $signed($unsigned($signed($signed(reg2813))));
                    end
                  else
                    begin
                      reg3203 <= ((reg2861[(3'h5):(2'h2)] ?
                              ($signed(reg3034) ?
                                  (reg2903 && reg2810) : (reg3157 >> (8'hb5))) : ({reg2739} ?
                                  $signed((8'hab)) : (forvar3160 ?
                                      (8'hb5) : reg2940))) ?
                          $signed(reg2845) : $signed((^~$signed(reg2841))));
                      reg3204 <= reg3113[(3'h4):(2'h2)];
                    end
                end
              else
                begin
                  if ($signed($unsigned(reg3096)))
                    begin
                      reg3198 <= $unsigned((reg2820[(3'h6):(3'h6)] ?
                          $unsigned(reg2917[(4'h8):(1'h0)]) : reg3128[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg3198 <= (+reg2739[(1'h0):(1'h0)]);
                    end
                  if ((reg2748 ? reg3027 : reg2942[(3'h6):(1'h1)]))
                    begin
                      reg3199 <= (reg3218 ?
                          reg3195[(1'h0):(1'h0)] : (reg2902[(3'h5):(2'h3)] ^ ($signed(reg2733) ?
                              reg2744 : reg2818[(3'h5):(3'h5)])));
                      reg3200 <= reg2884[(3'h7):(1'h1)];
                    end
                  else
                    begin
                      reg3199 <= (^($signed(reg2969) ?
                          $signed((reg3149 ? reg3053 : (8'hb4))) : (reg3183 ?
                              reg2834 : (reg2878 ? reg2924 : reg2831))));
                      reg3200 <= ($unsigned(reg3046) ?
                          $signed($signed($unsigned(reg1238))) : $signed((+{reg2935})));
                      reg3201 <= ((((reg2743 ? reg2903 : reg2744) ?
                              (reg3048 | (8'hb5)) : $signed(reg3188)) ?
                          ((reg2802 ?
                              reg2935 : reg2977) <<< reg3110[(4'hc):(4'hb)]) : ((reg3198 + reg2973) == reg3168)) >> (8'had));
                    end
                end
              for (forvar3207 = (1'h0); (forvar3207 < (2'h3)); forvar3207 = (forvar3207 + (1'h1)))
                begin
                  reg3208 <= $unsigned(({(^reg1216)} >= ((-reg1200) << (reg2968 == reg2763))));
                  reg3209 <= (($unsigned(reg2833) ?
                          reg3081 : $signed($signed(reg3175))) ?
                      (^~((reg2843 << reg3144) ?
                          reg2907 : $unsigned(reg3106))) : forvar3169);
                end
            end
        end
    end
  assign wire3223 = ($unsigned($unsigned($unsigned(reg2919))) ^~ reg3116[(4'h9):(3'h4)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1242
#(parameter param2705 = (((((8'h9d) ~^ (8'hb8)) ? (&(8'hb4)) : ((8'hb2) | (8'ha6))) ? (((8'hb7) || (8'ha0)) >> (~|(8'hae))) : (-((8'hba) ^~ (8'ha0)))) >> {{(~|(8'hae))}}))
(y, clk, wire1246, wire1245, wire1244, wire1243);
  output wire [(32'hc1c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire1246;
  input wire [(4'hb):(1'h0)] wire1245;
  input wire [(3'h7):(1'h0)] wire1244;
  input wire signed [(4'hb):(1'h0)] wire1243;
  wire signed [(3'h6):(1'h0)] wire2704;
  wire [(2'h2):(1'h0)] wire2703;
  wire signed [(3'h6):(1'h0)] wire2638;
  wire [(3'h5):(1'h0)] wire2586;
  wire [(2'h2):(1'h0)] wire1410;
  wire signed [(3'h7):(1'h0)] wire1409;
  wire signed [(3'h6):(1'h0)] wire1355;
  reg [(4'hd):(1'h0)] reg2702 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2701 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2700 = (1'h0);
  reg [(3'h7):(1'h0)] reg2699 = (1'h0);
  reg [(5'h10):(1'h0)] reg2698 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2695 = (1'h0);
  reg [(4'h9):(1'h0)] reg2694 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2693 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2691 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2690 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2689 = (1'h0);
  reg [(4'ha):(1'h0)] reg2687 = (1'h0);
  reg [(4'h8):(1'h0)] reg2686 = (1'h0);
  reg [(4'h8):(1'h0)] reg2685 = (1'h0);
  reg [(4'h8):(1'h0)] reg2683 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2682 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2680 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2678 = (1'h0);
  reg [(3'h5):(1'h0)] reg2677 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2676 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2675 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2674 = (1'h0);
  reg [(4'h8):(1'h0)] reg2673 = (1'h0);
  reg [(3'h7):(1'h0)] reg2672 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2671 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2670 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2666 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2661 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2667 = (1'h0);
  reg [(2'h2):(1'h0)] reg2665 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2664 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2663 = (1'h0);
  reg [(3'h7):(1'h0)] reg2662 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2660 = (1'h0);
  reg [(4'h9):(1'h0)] reg2659 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2658 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2657 = (1'h0);
  reg [(5'h10):(1'h0)] reg2656 = (1'h0);
  reg [(4'h8):(1'h0)] reg2655 = (1'h0);
  reg [(4'h9):(1'h0)] reg2651 = (1'h0);
  reg [(4'h9):(1'h0)] reg2650 = (1'h0);
  reg [(4'hb):(1'h0)] reg2649 = (1'h0);
  reg [(4'h8):(1'h0)] reg2648 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2647 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2646 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2644 = (1'h0);
  reg [(3'h7):(1'h0)] reg2643 = (1'h0);
  reg [(2'h3):(1'h0)] reg2637 = (1'h0);
  reg [(4'hb):(1'h0)] reg2636 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2634 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2633 = (1'h0);
  reg [(4'hb):(1'h0)] reg2616 = (1'h0);
  reg [(5'h10):(1'h0)] reg2632 = (1'h0);
  reg [(3'h5):(1'h0)] reg2631 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2630 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2628 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2625 = (1'h0);
  reg [(3'h7):(1'h0)] reg2624 = (1'h0);
  reg [(2'h2):(1'h0)] reg2623 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2622 = (1'h0);
  reg [(2'h2):(1'h0)] reg2621 = (1'h0);
  reg [(3'h7):(1'h0)] reg2620 = (1'h0);
  reg [(3'h5):(1'h0)] reg2619 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2618 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2617 = (1'h0);
  reg [(3'h5):(1'h0)] reg2615 = (1'h0);
  reg [(4'h9):(1'h0)] reg2614 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2612 = (1'h0);
  reg [(4'hd):(1'h0)] reg2611 = (1'h0);
  reg [(4'hd):(1'h0)] reg2610 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2609 = (1'h0);
  reg [(3'h7):(1'h0)] reg2607 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2606 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2605 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2604 = (1'h0);
  reg [(4'hd):(1'h0)] reg2603 = (1'h0);
  reg [(3'h5):(1'h0)] reg2602 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2601 = (1'h0);
  reg [(2'h3):(1'h0)] reg2596 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2594 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2592 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2600 = (1'h0);
  reg [(4'hf):(1'h0)] reg2599 = (1'h0);
  reg [(3'h4):(1'h0)] reg2598 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2597 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2595 = (1'h0);
  reg [(3'h6):(1'h0)] reg2593 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2591 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2590 = (1'h0);
  reg [(4'ha):(1'h0)] reg1388 = (1'h0);
  reg [(3'h4):(1'h0)] reg1373 = (1'h0);
  reg [(4'hc):(1'h0)] reg1372 = (1'h0);
  reg [(5'h10):(1'h0)] reg1369 = (1'h0);
  reg [(3'h7):(1'h0)] reg1366 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1358 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1356 = (1'h0);
  reg [(4'h9):(1'h0)] reg1357 = (1'h0);
  reg [(3'h7):(1'h0)] reg1404 = (1'h0);
  reg [(5'h10):(1'h0)] reg1399 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1408 = (1'h0);
  reg [(4'he):(1'h0)] reg1395 = (1'h0);
  reg [(3'h7):(1'h0)] reg1407 = (1'h0);
  reg [(5'h10):(1'h0)] reg1406 = (1'h0);
  reg [(4'ha):(1'h0)] reg1405 = (1'h0);
  reg [(3'h6):(1'h0)] reg1403 = (1'h0);
  reg [(3'h7):(1'h0)] reg1402 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1401 = (1'h0);
  reg [(4'hf):(1'h0)] reg1400 = (1'h0);
  reg [(2'h2):(1'h0)] reg1398 = (1'h0);
  reg [(5'h10):(1'h0)] reg1397 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1396 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1394 = (1'h0);
  reg [(3'h6):(1'h0)] reg1384 = (1'h0);
  reg [(5'h10):(1'h0)] reg1393 = (1'h0);
  reg [(3'h6):(1'h0)] reg1392 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1391 = (1'h0);
  reg [(4'hf):(1'h0)] reg1390 = (1'h0);
  reg [(3'h7):(1'h0)] reg1389 = (1'h0);
  reg [(3'h6):(1'h0)] reg1387 = (1'h0);
  reg [(3'h5):(1'h0)] reg1386 = (1'h0);
  reg [(2'h3):(1'h0)] reg1385 = (1'h0);
  reg [(4'hf):(1'h0)] reg1379 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1383 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1382 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1381 = (1'h0);
  reg [(4'ha):(1'h0)] reg1380 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1378 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1377 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1376 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1375 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1374 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1371 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1370 = (1'h0);
  reg [(4'h8):(1'h0)] reg1368 = (1'h0);
  reg [(4'h8):(1'h0)] reg1367 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1365 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1364 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1362 = (1'h0);
  reg [(4'he):(1'h0)] reg1361 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1360 = (1'h0);
  reg [(3'h5):(1'h0)] reg1359 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1354 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1353 = (1'h0);
  reg [(3'h6):(1'h0)] reg1331 = (1'h0);
  reg [(3'h5):(1'h0)] reg1352 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1351 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1350 = (1'h0);
  reg [(4'hd):(1'h0)] reg1348 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1347 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1346 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1345 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1343 = (1'h0);
  reg [(4'hd):(1'h0)] reg1342 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1341 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1339 = (1'h0);
  reg [(4'h8):(1'h0)] reg1338 = (1'h0);
  reg [(4'ha):(1'h0)] reg1337 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1336 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1335 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1334 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1333 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1332 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1328 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1330 = (1'h0);
  reg [(5'h10):(1'h0)] reg1329 = (1'h0);
  reg [(3'h5):(1'h0)] reg1327 = (1'h0);
  reg [(3'h6):(1'h0)] reg1326 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1325 = (1'h0);
  reg [(4'he):(1'h0)] reg1324 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1323 = (1'h0);
  reg [(3'h7):(1'h0)] reg1322 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1321 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1320 = (1'h0);
  reg [(2'h3):(1'h0)] reg1319 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1317 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1315 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1314 = (1'h0);
  reg [(3'h5):(1'h0)] reg1313 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1312 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1299 = (1'h0);
  reg [(3'h4):(1'h0)] reg1310 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1309 = (1'h0);
  reg [(4'hd):(1'h0)] reg1308 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1307 = (1'h0);
  reg [(3'h4):(1'h0)] reg1303 = (1'h0);
  reg [(4'he):(1'h0)] reg1293 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1287 = (1'h0);
  reg [(2'h2):(1'h0)] reg1306 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1305 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1304 = (1'h0);
  reg [(5'h10):(1'h0)] reg1302 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1301 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1300 = (1'h0);
  reg [(3'h4):(1'h0)] reg1298 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1297 = (1'h0);
  reg [(4'h8):(1'h0)] reg1296 = (1'h0);
  reg [(2'h3):(1'h0)] reg1295 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1294 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1292 = (1'h0);
  reg [(2'h3):(1'h0)] reg1291 = (1'h0);
  reg [(4'hf):(1'h0)] reg1290 = (1'h0);
  reg [(4'hc):(1'h0)] reg1289 = (1'h0);
  reg [(4'hc):(1'h0)] reg1288 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1286 = (1'h0);
  reg [(4'ha):(1'h0)] reg1285 = (1'h0);
  reg [(3'h6):(1'h0)] reg1275 = (1'h0);
  reg [(5'h10):(1'h0)] reg1271 = (1'h0);
  reg [(3'h4):(1'h0)] reg1270 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1255 = (1'h0);
  reg [(3'h6):(1'h0)] reg1284 = (1'h0);
  reg [(5'h10):(1'h0)] reg1283 = (1'h0);
  reg [(4'h9):(1'h0)] reg1282 = (1'h0);
  reg [(4'hb):(1'h0)] reg1281 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1280 = (1'h0);
  reg [(3'h5):(1'h0)] reg1279 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1278 = (1'h0);
  reg [(4'h9):(1'h0)] reg1277 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1276 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1274 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1273 = (1'h0);
  reg [(2'h2):(1'h0)] reg1272 = (1'h0);
  reg [(4'h9):(1'h0)] reg1266 = (1'h0);
  reg [(4'h8):(1'h0)] reg1269 = (1'h0);
  reg [(3'h5):(1'h0)] reg1268 = (1'h0);
  reg [(4'h8):(1'h0)] reg1267 = (1'h0);
  reg [(3'h7):(1'h0)] reg1265 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1264 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1263 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1262 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1261 = (1'h0);
  reg [(4'hf):(1'h0)] reg1260 = (1'h0);
  reg [(4'hb):(1'h0)] reg1259 = (1'h0);
  reg [(4'hd):(1'h0)] reg1258 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1257 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1256 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1249 = (1'h0);
  reg [(3'h4):(1'h0)] reg1254 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1253 = (1'h0);
  reg [(4'hd):(1'h0)] reg1252 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1251 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1250 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1247 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2697 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2696 = (1'h0);
  reg [(4'he):(1'h0)] forvar2692 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2688 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2684 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2681 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2679 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2669 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2668 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2663 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2666 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2661 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2654 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2653 = (1'h0);
  reg [(4'he):(1'h0)] forvar2652 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2645 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2642 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2641 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2640 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2639 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2635 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2614 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2629 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2627 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2626 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2616 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2613 = (1'h0);
  reg [(4'he):(1'h0)] forvar2602 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2608 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2593 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2590 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2596 = (1'h0);
  reg [(4'he):(1'h0)] forvar2594 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2592 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2589 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2588 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1387 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1386 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1380 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1378 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1375 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1370 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1371 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1367 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1360 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1403 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1402 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1398 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1404 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1399 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1395 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1388 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1384 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1377 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1379 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1373 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1372 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1369 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1366 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1363 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1358 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1357 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1356 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1326 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1325 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1349 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1344 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1340 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1331 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1328 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1318 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1316 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1311 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1306 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1303 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1299 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1293 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1287 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1268 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1259 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1254 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1282 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1278 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1272 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1269 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1264 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1260 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1257 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1253 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1252 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1275 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1271 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1270 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1266 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1255 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1249 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1248 = (1'h0);
  assign y = {wire2704,
                 wire2703,
                 wire2638,
                 wire2586,
                 wire1410,
                 wire1409,
                 wire1355,
                 reg2702,
                 reg2701,
                 reg2700,
                 reg2699,
                 reg2698,
                 reg2695,
                 reg2694,
                 reg2693,
                 reg2691,
                 reg2690,
                 reg2689,
                 reg2687,
                 reg2686,
                 reg2685,
                 reg2683,
                 reg2682,
                 reg2680,
                 reg2678,
                 reg2677,
                 reg2676,
                 reg2675,
                 reg2674,
                 reg2673,
                 reg2672,
                 reg2671,
                 reg2670,
                 reg2666,
                 reg2661,
                 reg2667,
                 reg2665,
                 reg2664,
                 reg2663,
                 reg2662,
                 reg2660,
                 reg2659,
                 reg2658,
                 reg2657,
                 reg2656,
                 reg2655,
                 reg2651,
                 reg2650,
                 reg2649,
                 reg2648,
                 reg2647,
                 reg2646,
                 reg2644,
                 reg2643,
                 reg2637,
                 reg2636,
                 reg2634,
                 reg2633,
                 reg2616,
                 reg2632,
                 reg2631,
                 reg2630,
                 reg2628,
                 reg2625,
                 reg2624,
                 reg2623,
                 reg2622,
                 reg2621,
                 reg2620,
                 reg2619,
                 reg2618,
                 reg2617,
                 reg2615,
                 reg2614,
                 reg2612,
                 reg2611,
                 reg2610,
                 reg2609,
                 reg2607,
                 reg2606,
                 reg2605,
                 reg2604,
                 reg2603,
                 reg2602,
                 reg2601,
                 reg2596,
                 reg2594,
                 reg2592,
                 reg2600,
                 reg2599,
                 reg2598,
                 reg2597,
                 reg2595,
                 reg2593,
                 reg2591,
                 reg2590,
                 reg1388,
                 reg1373,
                 reg1372,
                 reg1369,
                 reg1366,
                 reg1358,
                 reg1356,
                 reg1357,
                 reg1404,
                 reg1399,
                 reg1408,
                 reg1395,
                 reg1407,
                 reg1406,
                 reg1405,
                 reg1403,
                 reg1402,
                 reg1401,
                 reg1400,
                 reg1398,
                 reg1397,
                 reg1396,
                 reg1394,
                 reg1384,
                 reg1393,
                 reg1392,
                 reg1391,
                 reg1390,
                 reg1389,
                 reg1387,
                 reg1386,
                 reg1385,
                 reg1379,
                 reg1383,
                 reg1382,
                 reg1381,
                 reg1380,
                 reg1378,
                 reg1377,
                 reg1376,
                 reg1375,
                 reg1374,
                 reg1371,
                 reg1370,
                 reg1368,
                 reg1367,
                 reg1365,
                 reg1364,
                 reg1362,
                 reg1361,
                 reg1360,
                 reg1359,
                 reg1354,
                 reg1353,
                 reg1331,
                 reg1352,
                 reg1351,
                 reg1350,
                 reg1348,
                 reg1347,
                 reg1346,
                 reg1345,
                 reg1343,
                 reg1342,
                 reg1341,
                 reg1339,
                 reg1338,
                 reg1337,
                 reg1336,
                 reg1335,
                 reg1334,
                 reg1333,
                 reg1332,
                 reg1328,
                 reg1330,
                 reg1329,
                 reg1327,
                 reg1326,
                 reg1325,
                 reg1324,
                 reg1323,
                 reg1322,
                 reg1321,
                 reg1320,
                 reg1319,
                 reg1317,
                 reg1315,
                 reg1314,
                 reg1313,
                 reg1312,
                 reg1299,
                 reg1310,
                 reg1309,
                 reg1308,
                 reg1307,
                 reg1303,
                 reg1293,
                 reg1287,
                 reg1306,
                 reg1305,
                 reg1304,
                 reg1302,
                 reg1301,
                 reg1300,
                 reg1298,
                 reg1297,
                 reg1296,
                 reg1295,
                 reg1294,
                 reg1292,
                 reg1291,
                 reg1290,
                 reg1289,
                 reg1288,
                 reg1286,
                 reg1285,
                 reg1275,
                 reg1271,
                 reg1270,
                 reg1255,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1281,
                 reg1280,
                 reg1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 reg1274,
                 reg1273,
                 reg1272,
                 reg1266,
                 reg1269,
                 reg1268,
                 reg1267,
                 reg1265,
                 reg1264,
                 reg1263,
                 reg1262,
                 reg1261,
                 reg1260,
                 reg1259,
                 reg1258,
                 reg1257,
                 reg1256,
                 reg1249,
                 reg1254,
                 reg1253,
                 reg1252,
                 reg1251,
                 reg1250,
                 reg1247,
                 forvar2697,
                 forvar2696,
                 forvar2692,
                 forvar2688,
                 forvar2684,
                 forvar2681,
                 forvar2679,
                 forvar2669,
                 forvar2668,
                 forvar2663,
                 forvar2666,
                 forvar2661,
                 forvar2654,
                 forvar2653,
                 forvar2652,
                 forvar2645,
                 forvar2642,
                 forvar2641,
                 forvar2640,
                 forvar2639,
                 forvar2635,
                 forvar2614,
                 forvar2629,
                 forvar2627,
                 forvar2626,
                 forvar2616,
                 forvar2613,
                 forvar2602,
                 forvar2608,
                 forvar2593,
                 forvar2590,
                 forvar2596,
                 forvar2594,
                 forvar2592,
                 forvar2589,
                 forvar2588,
                 forvar1387,
                 forvar1386,
                 forvar1380,
                 forvar1378,
                 forvar1375,
                 forvar1370,
                 forvar1371,
                 forvar1367,
                 forvar1360,
                 forvar1403,
                 forvar1402,
                 forvar1398,
                 forvar1404,
                 forvar1399,
                 forvar1395,
                 forvar1388,
                 forvar1384,
                 forvar1377,
                 forvar1379,
                 forvar1373,
                 forvar1372,
                 forvar1369,
                 forvar1366,
                 forvar1363,
                 forvar1358,
                 forvar1357,
                 forvar1356,
                 forvar1326,
                 forvar1325,
                 forvar1349,
                 forvar1344,
                 forvar1340,
                 forvar1331,
                 forvar1328,
                 forvar1318,
                 forvar1316,
                 forvar1311,
                 forvar1306,
                 forvar1303,
                 forvar1299,
                 forvar1293,
                 forvar1287,
                 forvar1268,
                 forvar1259,
                 forvar1254,
                 forvar1282,
                 forvar1278,
                 forvar1272,
                 forvar1269,
                 forvar1264,
                 forvar1260,
                 forvar1257,
                 forvar1253,
                 forvar1252,
                 forvar1275,
                 forvar1271,
                 forvar1270,
                 forvar1266,
                 forvar1255,
                 forvar1249,
                 forvar1248,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1247 <= ((8'hac) ?
          {({(8'ha3)} ?
                  wire1246 : $unsigned((8'hb2)))} : wire1243[(2'h2):(2'h2)]);
      if ((+(8'hb8)))
        begin
          for (forvar1248 = (1'h0); (forvar1248 < (2'h3)); forvar1248 = (forvar1248 + (1'h1)))
            begin
              if (wire1245)
                begin
                  for (forvar1249 = (1'h0); (forvar1249 < (2'h3)); forvar1249 = (forvar1249 + (1'h1)))
                    begin
                      reg1250 <= $unsigned(forvar1249);
                      reg1251 <= ($unsigned($signed((wire1245 + reg1247))) > {forvar1248[(3'h4):(3'h4)]});
                      reg1252 <= wire1243;
                      reg1253 <= ((reg1252 <= ($unsigned(wire1246) >> (~&wire1245))) & ($signed($signed(reg1247)) ?
                          (~&forvar1249) : (^~(reg1250 ? reg1250 : wire1246))));
                    end
                  reg1254 <= $unsigned(wire1246[(2'h2):(2'h2)]);
                end
              else
                begin
                  if ($signed((reg1254 ?
                      ((+wire1243) ^ (wire1245 ?
                          reg1253 : reg1252)) : $signed((reg1247 ?
                          reg1254 : reg1253)))))
                    begin
                      reg1249 <= (~^(~^$unsigned(wire1245)));
                      reg1250 <= $signed(reg1247);
                    end
                  else
                    begin
                      reg1249 <= (-(8'haa));
                      reg1250 <= ($signed(wire1244) - $unsigned($unsigned($unsigned(wire1246))));
                    end
                  if ($signed((wire1246 > ({wire1245} <<< (reg1254 ?
                      wire1246 : reg1254)))))
                    begin
                      reg1251 <= ($signed(((!(8'h9c)) << wire1244)) || $signed(forvar1249[(4'hd):(4'ha)]));
                      reg1252 <= $unsigned($unsigned(reg1253));
                      reg1253 <= (((reg1253 + $unsigned(reg1247)) | $unsigned((forvar1248 ~^ wire1243))) + (+((reg1250 >= reg1252) ?
                          $signed(forvar1249) : (^forvar1249))));
                      reg1254 <= $signed((|(wire1244 ?
                          (reg1249 ? reg1253 : reg1247) : $signed(reg1247))));
                    end
                  else
                    begin
                      reg1251 <= ((~&(-$unsigned(reg1253))) == $unsigned(reg1253));
                    end
                  for (forvar1255 = (1'h0); (forvar1255 < (1'h1)); forvar1255 = (forvar1255 + (1'h1)))
                    begin
                      reg1256 <= (forvar1248[(4'hf):(4'he)] ^~ $unsigned({{forvar1248}}));
                      reg1257 <= $signed($unsigned(reg1249));
                      reg1258 <= $unsigned(((~&(forvar1255 << (8'ha8))) || ($unsigned(wire1244) ~^ $signed(wire1243))));
                      reg1259 <= reg1249[(1'h0):(1'h0)];
                    end
                  reg1260 <= wire1243;
                end
              if ((!(reg1247 >>> $unsigned(reg1258))))
                begin
                  reg1261 <= wire1243;
                  if (($signed((~wire1244[(1'h1):(1'h1)])) ?
                      reg1256[(1'h1):(1'h0)] : (~&{(forvar1248 ?
                              reg1258 : (8'ha9))})))
                    begin
                      reg1262 <= $unsigned((!$signed(reg1249[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg1262 <= $unsigned((((reg1251 ? reg1254 : reg1253) ?
                          reg1247 : (~&reg1257)) & $signed((reg1250 ?
                          forvar1255 : reg1262))));
                    end
                  if ((reg1258 & ((&$signed((8'hab))) ?
                      (~$unsigned(reg1249)) : {wire1243})))
                    begin
                      reg1263 <= ((|reg1257[(3'h6):(3'h5)]) & reg1254);
                      reg1264 <= $signed($signed($unsigned((reg1253 ?
                          reg1260 : wire1245))));
                      reg1265 <= (~reg1252);
                    end
                  else
                    begin
                      reg1263 <= forvar1255;
                    end
                  for (forvar1266 = (1'h0); (forvar1266 < (1'h0)); forvar1266 = (forvar1266 + (1'h1)))
                    begin
                      reg1267 <= (~^(reg1254[(1'h0):(1'h0)] ^~ $signed(reg1260)));
                      reg1268 <= reg1260[(4'hc):(4'hc)];
                      reg1269 <= (-$signed((^~$signed(wire1243))));
                    end
                end
              else
                begin
                  if ((|(~^(reg1254[(3'h4):(1'h0)] < $signed(reg1265)))))
                    begin
                      reg1261 <= (~((!reg1252[(3'h6):(3'h4)]) ?
                          (((8'ha0) <= reg1258) * (+reg1250)) : forvar1248[(4'he):(2'h2)]));
                      reg1262 <= wire1243[(2'h2):(1'h0)];
                      reg1263 <= $unsigned(reg1268);
                    end
                  else
                    begin
                      reg1261 <= $unsigned($signed(reg1252[(3'h6):(3'h5)]));
                      reg1262 <= $unsigned({reg1261[(4'hb):(1'h1)]});
                      reg1263 <= $unsigned(($unsigned($unsigned((8'ha4))) ^ $signed((forvar1266 << reg1261))));
                      reg1264 <= (^~$unsigned(reg1269));
                    end
                  if (((|wire1245) ?
                      $signed((^~((8'hb1) ?
                          reg1252 : reg1254))) : ($signed(((8'h9e) >= wire1245)) ~^ $signed(reg1254[(2'h3):(1'h1)]))))
                    begin
                      reg1265 <= {((-reg1258) ?
                              reg1258[(4'hd):(3'h5)] : $unsigned($unsigned(reg1251)))};
                    end
                  else
                    begin
                      reg1265 <= $unsigned($unsigned(reg1247[(1'h1):(1'h0)]));
                      reg1266 <= reg1263;
                      reg1267 <= wire1246[(1'h1):(1'h1)];
                      reg1268 <= $unsigned(reg1250[(4'hb):(1'h1)]);
                    end
                end
              for (forvar1270 = (1'h0); (forvar1270 < (1'h1)); forvar1270 = (forvar1270 + (1'h1)))
                begin
                  for (forvar1271 = (1'h0); (forvar1271 < (2'h3)); forvar1271 = (forvar1271 + (1'h1)))
                    begin
                      reg1272 <= reg1253[(2'h2):(1'h1)];
                      reg1273 <= reg1262[(3'h4):(2'h2)];
                      reg1274 <= reg1257[(4'h8):(2'h2)];
                    end
                end
              if (((($unsigned(reg1257) ?
                      (reg1260 ?
                          reg1266 : (8'hac)) : reg1259[(3'h7):(2'h2)]) ^ $signed($signed(reg1253))) ?
                  reg1261 : $unsigned(((~|reg1259) >>> $unsigned(reg1247)))))
                begin
                  for (forvar1275 = (1'h0); (forvar1275 < (1'h1)); forvar1275 = (forvar1275 + (1'h1)))
                    begin
                      reg1276 <= $signed(reg1273);
                      reg1277 <= ($unsigned($signed($unsigned(reg1265))) || ((~(+forvar1255)) >> $signed((forvar1266 * wire1246))));
                      reg1278 <= reg1256;
                      reg1279 <= (~|reg1257);
                    end
                end
              else
                begin
                  for (forvar1275 = (1'h0); (forvar1275 < (1'h1)); forvar1275 = (forvar1275 + (1'h1)))
                    begin
                      reg1276 <= (reg1247[(1'h0):(1'h0)] ?
                          ($unsigned((~(8'h9c))) < ($unsigned(reg1274) ?
                              reg1267 : reg1265)) : ((|(reg1268 << reg1259)) | $unsigned({forvar1271})));
                      reg1277 <= ($signed($unsigned($unsigned((8'h9c)))) ?
                          (&($unsigned((8'ha1)) >= (reg1273 >> reg1247))) : (&((reg1251 ?
                              forvar1270 : reg1262) < $unsigned(reg1256))));
                    end
                  if (($signed(($unsigned(reg1253) > $unsigned((8'hb8)))) ?
                      (reg1278[(3'h5):(3'h5)] ?
                          ((reg1256 >>> reg1262) ?
                              $signed((8'hb2)) : $signed(forvar1266)) : (~|$unsigned(reg1267))) : $unsigned($unsigned((forvar1248 ?
                          reg1253 : (8'hb1))))))
                    begin
                      reg1278 <= ($unsigned((^(forvar1266 >> reg1269))) <<< (&(forvar1249[(3'h4):(2'h2)] ?
                          (!reg1266) : (forvar1255 ? wire1245 : reg1274))));
                      reg1279 <= ((^~{(reg1261 <= reg1265)}) ?
                          forvar1248[(4'ha):(3'h6)] : ((reg1272[(2'h2):(1'h0)] <= $signed(reg1278)) <<< (forvar1248 ?
                              $signed(reg1247) : (forvar1249 ?
                                  reg1254 : forvar1270))));
                      reg1280 <= $unsigned((($signed(wire1245) ?
                          reg1251[(2'h3):(2'h3)] : $signed((8'haf))) >= reg1266));
                      reg1281 <= (reg1264 > reg1280);
                    end
                  else
                    begin
                      reg1278 <= $unsigned($unsigned($signed($signed(reg1274))));
                      reg1279 <= (8'h9f);
                      reg1280 <= (^$unsigned($signed((reg1263 ?
                          reg1280 : forvar1266))));
                      reg1281 <= (+{reg1249});
                    end
                  if (reg1260)
                    begin
                      reg1282 <= ({(((8'hb7) >= forvar1249) ?
                                  $signed(reg1261) : (reg1254 >>> forvar1249))} ?
                          $unsigned($signed($signed(wire1245))) : reg1274[(3'h5):(1'h1)]);
                      reg1283 <= (&$signed($unsigned(((8'hb7) ?
                          reg1267 : reg1266))));
                      reg1284 <= {$unsigned(((|reg1279) ?
                              $unsigned(forvar1271) : (8'hb4)))};
                    end
                  else
                    begin
                      reg1282 <= $signed((reg1266[(1'h0):(1'h0)] > (((8'hb9) ?
                          forvar1248 : forvar1248) != reg1262)));
                      reg1283 <= $unsigned($signed((8'ha6)));
                      reg1284 <= (~reg1257);
                    end
                end
            end
        end
      else
        begin
          if (($signed(((reg1265 <<< reg1257) ?
              {reg1269} : reg1272[(1'h0):(1'h0)])) <<< reg1257))
            begin
              for (forvar1248 = (1'h0); (forvar1248 < (1'h0)); forvar1248 = (forvar1248 + (1'h1)))
                begin
                  for (forvar1249 = (1'h0); (forvar1249 < (2'h3)); forvar1249 = (forvar1249 + (1'h1)))
                    begin
                      reg1250 <= $unsigned(reg1282);
                      reg1251 <= (($signed(reg1273) ?
                          (!$unsigned(forvar1248)) : $unsigned((~|forvar1271))) + {(+$unsigned(reg1269))});
                    end
                end
              for (forvar1252 = (1'h0); (forvar1252 < (2'h3)); forvar1252 = (forvar1252 + (1'h1)))
                begin
                  for (forvar1253 = (1'h0); (forvar1253 < (1'h1)); forvar1253 = (forvar1253 + (1'h1)))
                    begin
                      reg1254 <= {$signed($unsigned((reg1278 ?
                              forvar1255 : reg1259)))};
                    end
                  if (reg1251)
                    begin
                      reg1255 <= $signed(reg1273[(4'h9):(3'h4)]);
                      reg1256 <= reg1280[(4'hd):(3'h7)];
                    end
                  else
                    begin
                      reg1255 <= forvar1248;
                      reg1256 <= $signed({reg1256[(4'hc):(4'h8)]});
                    end
                  for (forvar1257 = (1'h0); (forvar1257 < (1'h1)); forvar1257 = (forvar1257 + (1'h1)))
                    begin
                      reg1258 <= ($signed((~(!forvar1275))) >>> ($signed((8'hab)) ?
                          $unsigned($signed(reg1256)) : (8'hb7)));
                      reg1259 <= (^{(^~$signed(reg1282))});
                    end
                end
              for (forvar1260 = (1'h0); (forvar1260 < (1'h0)); forvar1260 = (forvar1260 + (1'h1)))
                begin
                  if ($signed($signed((+(~forvar1248)))))
                    begin
                      reg1261 <= (($signed((8'ha5)) ?
                          $signed(reg1279) : $signed((^forvar1266))) >= forvar1266);
                      reg1262 <= {forvar1257[(2'h3):(1'h0)]};
                    end
                  else
                    begin
                      reg1261 <= (wire1245[(4'h8):(4'h8)] <= $signed(reg1261[(4'ha):(2'h3)]));
                      reg1262 <= (+$unsigned(reg1274));
                    end
                  reg1263 <= $unsigned($unsigned((^$signed(reg1272))));
                  for (forvar1264 = (1'h0); (forvar1264 < (2'h2)); forvar1264 = (forvar1264 + (1'h1)))
                    begin
                      reg1265 <= $unsigned($signed($signed(reg1283[(2'h3):(2'h2)])));
                      reg1266 <= (8'hb6);
                      reg1267 <= ($signed($unsigned($unsigned(reg1256))) ?
                          forvar1257[(1'h0):(1'h0)] : (wire1243 <= reg1263));
                      reg1268 <= (reg1283 ?
                          forvar1266 : {{(forvar1275 - reg1272)}});
                    end
                  for (forvar1269 = (1'h0); (forvar1269 < (2'h2)); forvar1269 = (forvar1269 + (1'h1)))
                    begin
                      reg1270 <= ($unsigned((+(reg1277 >= reg1264))) ?
                          reg1251[(4'hd):(4'hb)] : ($signed($signed((8'hb3))) < reg1262[(4'h8):(3'h4)]));
                      reg1271 <= (^(&(reg1259[(3'h5):(2'h2)] ~^ (!reg1277))));
                    end
                end
              for (forvar1272 = (1'h0); (forvar1272 < (2'h2)); forvar1272 = (forvar1272 + (1'h1)))
                begin
                  reg1273 <= ((8'hba) >>> forvar1255[(1'h1):(1'h0)]);
                  if ($signed($signed(reg1257[(1'h0):(1'h0)])))
                    begin
                      reg1274 <= $signed(reg1263);
                    end
                  else
                    begin
                      reg1274 <= $unsigned($signed($signed(reg1252[(2'h2):(1'h1)])));
                      reg1275 <= $unsigned($signed(reg1261[(3'h7):(3'h4)]));
                      reg1276 <= reg1254[(3'h4):(1'h1)];
                      reg1277 <= ($unsigned({{reg1266}}) ?
                          (!forvar1257[(2'h2):(2'h2)]) : (~^reg1262[(4'h8):(3'h5)]));
                    end
                  for (forvar1278 = (1'h0); (forvar1278 < (2'h2)); forvar1278 = (forvar1278 + (1'h1)))
                    begin
                      reg1279 <= $unsigned(($unsigned({reg1272}) ?
                          $unsigned((~&reg1251)) : reg1249));
                      reg1280 <= forvar1266[(4'h9):(3'h4)];
                      reg1281 <= ($signed($unsigned($signed(reg1263))) ?
                          ((8'hb9) && (~&(~reg1276))) : (^reg1269));
                    end
                  for (forvar1282 = (1'h0); (forvar1282 < (2'h2)); forvar1282 = (forvar1282 + (1'h1)))
                    begin
                      reg1283 <= {{{forvar1255[(2'h2):(1'h1)]}}};
                      reg1284 <= ((~|(reg1247[(1'h1):(1'h0)] ?
                          ((8'hb3) * reg1279) : reg1281)) >>> $signed(($signed(reg1283) << $signed(reg1256))));
                      reg1285 <= (&($unsigned((8'h9c)) ?
                          forvar1269 : forvar1252));
                      reg1286 <= (&(forvar1266 ?
                          {reg1279[(3'h5):(2'h3)]} : (~(reg1256 << (8'ha0)))));
                    end
                end
            end
          else
            begin
              for (forvar1248 = (1'h0); (forvar1248 < (1'h1)); forvar1248 = (forvar1248 + (1'h1)))
                begin
                  if (((^(+$signed(reg1260))) ?
                      ((reg1260 ?
                          $unsigned(reg1249) : (reg1278 ?
                              reg1277 : reg1252)) != $signed((reg1278 || reg1271))) : forvar1266[(4'ha):(3'h6)]))
                    begin
                      reg1249 <= (8'h9c);
                      reg1250 <= (reg1264[(1'h0):(1'h0)] ?
                          reg1262 : $unsigned(reg1268[(1'h1):(1'h0)]));
                      reg1251 <= (~|(^(-{reg1269})));
                    end
                  else
                    begin
                      reg1249 <= $signed($unsigned((((8'haf) ?
                              forvar1260 : reg1256) ?
                          $signed((8'hae)) : (reg1286 ?
                              forvar1266 : reg1249))));
                      reg1250 <= (~&$signed((~^(~&reg1260))));
                      reg1251 <= forvar1252[(2'h3):(2'h2)];
                      reg1252 <= forvar1249;
                    end
                  reg1253 <= wire1246[(1'h0):(1'h0)];
                end
              for (forvar1254 = (1'h0); (forvar1254 < (1'h1)); forvar1254 = (forvar1254 + (1'h1)))
                begin
                  for (forvar1255 = (1'h0); (forvar1255 < (2'h3)); forvar1255 = (forvar1255 + (1'h1)))
                    begin
                      reg1256 <= (~^reg1264[(2'h3):(2'h2)]);
                      reg1257 <= ($unsigned(({(8'hb8)} >= (+forvar1249))) ?
                          ($unsigned((reg1252 ?
                              forvar1260 : reg1270)) & forvar1249[(3'h6):(3'h6)]) : forvar1255[(2'h2):(1'h0)]);
                      reg1258 <= ($unsigned((!(reg1280 ? wire1245 : reg1256))) ?
                          wire1244[(3'h6):(2'h2)] : reg1252);
                    end
                  for (forvar1259 = (1'h0); (forvar1259 < (2'h3)); forvar1259 = (forvar1259 + (1'h1)))
                    begin
                      reg1260 <= forvar1271[(3'h5):(2'h3)];
                      reg1261 <= {$signed($signed((+reg1276)))};
                      reg1262 <= reg1263;
                      reg1263 <= {forvar1252[(3'h5):(1'h1)]};
                    end
                end
              if (reg1261)
                begin
                  for (forvar1264 = (1'h0); (forvar1264 < (2'h2)); forvar1264 = (forvar1264 + (1'h1)))
                    begin
                      reg1265 <= reg1267[(2'h3):(1'h1)];
                      reg1266 <= wire1246[(1'h1):(1'h0)];
                      reg1267 <= $signed($signed((8'hac)));
                      reg1268 <= {$signed((~|(~forvar1257)))};
                    end
                  for (forvar1269 = (1'h0); (forvar1269 < (1'h1)); forvar1269 = (forvar1269 + (1'h1)))
                    begin
                      reg1270 <= (-$unsigned($unsigned((reg1255 ?
                          forvar1260 : forvar1253))));
                      reg1271 <= ({forvar1266[(3'h4):(2'h2)]} << reg1268[(3'h5):(1'h0)]);
                    end
                  reg1272 <= ($unsigned($unsigned($signed((8'ha1)))) || {reg1255});
                  if ((8'hab))
                    begin
                      reg1273 <= ((-$unsigned((reg1282 ?
                              forvar1269 : reg1256))) ?
                          $signed(((~&forvar1275) ?
                              (forvar1259 ?
                                  forvar1255 : reg1275) : reg1268[(1'h0):(1'h0)])) : forvar1254[(1'h1):(1'h0)]);
                      reg1274 <= (^($unsigned({(8'hb5)}) && $signed($signed(reg1270))));
                      reg1275 <= ((~^forvar1278) ? forvar1248 : forvar1275);
                    end
                  else
                    begin
                      reg1273 <= reg1271[(4'he):(4'h8)];
                      reg1274 <= $unsigned({reg1267});
                    end
                end
              else
                begin
                  if (({reg1255[(1'h0):(1'h0)]} ~^ {$signed($signed(forvar1275))}))
                    begin
                      reg1264 <= $signed(reg1255);
                    end
                  else
                    begin
                      reg1264 <= (reg1269[(3'h4):(3'h4)] < ((forvar1275 ?
                              reg1278[(2'h3):(2'h2)] : reg1274[(2'h3):(2'h2)]) ?
                          reg1285[(3'h6):(1'h0)] : $unsigned(reg1283[(3'h7):(2'h2)])));
                      reg1265 <= ($signed((reg1249[(2'h3):(2'h2)] | (+reg1286))) <= ($signed(forvar1269[(4'h8):(2'h2)]) > reg1278));
                      reg1266 <= reg1276;
                      reg1267 <= $signed(reg1283);
                    end
                  for (forvar1268 = (1'h0); (forvar1268 < (2'h2)); forvar1268 = (forvar1268 + (1'h1)))
                    begin
                      reg1269 <= {{(+(^~wire1245))}};
                      reg1270 <= reg1261;
                      reg1271 <= (((8'ha5) ?
                              reg1266 : $unsigned($unsigned((8'ha5)))) ?
                          $unsigned($signed((reg1283 ?
                              forvar1264 : reg1272))) : $unsigned(($unsigned((8'hb0)) >>> {(8'ha3)})));
                      reg1272 <= $unsigned(((reg1284 ? forvar1260 : reg1251) ?
                          (^~((8'ha9) == (8'hb5))) : (((8'h9e) & reg1247) >>> reg1260[(4'h8):(2'h2)])));
                    end
                end
            end
          if ($signed(reg1286))
            begin
              for (forvar1287 = (1'h0); (forvar1287 < (1'h0)); forvar1287 = (forvar1287 + (1'h1)))
                begin
                  if ({((8'hb4) >> (+{forvar1253}))})
                    begin
                      reg1288 <= (~$unsigned($signed($unsigned(reg1279))));
                    end
                  else
                    begin
                      reg1288 <= ((&(&(!reg1263))) ?
                          $unsigned((~|(reg1249 ?
                              (8'ha0) : (8'ha5)))) : $unsigned(((reg1259 ?
                                  forvar1287 : reg1285) ?
                              reg1247 : reg1257[(2'h2):(1'h0)])));
                      reg1289 <= (~^reg1271);
                    end
                  if (($signed(forvar1260) ?
                      ({reg1263} ?
                          reg1253 : (~&$signed(forvar1249))) : (8'h9c)))
                    begin
                      reg1290 <= $unsigned(reg1286);
                      reg1291 <= reg1247;
                      reg1292 <= $signed($unsigned(reg1288));
                    end
                  else
                    begin
                      reg1290 <= (-(reg1247[(2'h3):(1'h0)] + (~^forvar1248[(2'h2):(1'h1)])));
                    end
                end
              for (forvar1293 = (1'h0); (forvar1293 < (1'h1)); forvar1293 = (forvar1293 + (1'h1)))
                begin
                  reg1294 <= (($unsigned({forvar1260}) | reg1274[(4'h8):(3'h5)]) ?
                      $signed((-(reg1252 ?
                          forvar1252 : (8'hb3)))) : (!$unsigned(wire1243)));
                  if ($signed(reg1274[(3'h5):(3'h4)]))
                    begin
                      reg1295 <= forvar1253[(2'h2):(1'h0)];
                      reg1296 <= reg1285;
                    end
                  else
                    begin
                      reg1295 <= forvar1249[(4'ha):(3'h7)];
                      reg1296 <= (~|((forvar1254 >> (~^reg1266)) >>> ((forvar1275 ?
                          reg1285 : reg1261) ^ ((8'h9d) ?
                          forvar1257 : reg1254))));
                      reg1297 <= $unsigned({(forvar1260[(3'h5):(2'h3)] ?
                              (reg1280 > reg1276) : forvar1269[(2'h2):(1'h1)])});
                      reg1298 <= (8'ha7);
                    end
                  for (forvar1299 = (1'h0); (forvar1299 < (2'h2)); forvar1299 = (forvar1299 + (1'h1)))
                    begin
                      reg1300 <= (|(reg1282 ?
                          (~(^~forvar1264)) : (~^(^~(8'hac)))));
                      reg1301 <= ((~|{$signed(reg1295)}) ^~ (reg1288 ?
                          ((forvar1257 <<< forvar1287) ?
                              forvar1253[(2'h3):(2'h2)] : reg1264[(1'h0):(1'h0)]) : ((^forvar1275) ?
                              {reg1249} : (reg1263 ?
                                  forvar1254 : forvar1260))));
                    end
                  reg1302 <= ($unsigned(reg1255) & ($signed($unsigned((8'ha0))) ?
                      $signed($signed(forvar1257)) : (~&reg1253)));
                end
              for (forvar1303 = (1'h0); (forvar1303 < (1'h1)); forvar1303 = (forvar1303 + (1'h1)))
                begin
                  if ((forvar1303[(3'h5):(2'h2)] || reg1284[(3'h4):(2'h2)]))
                    begin
                      reg1304 <= ((8'ha8) <= $unsigned($unsigned((~&forvar1255))));
                      reg1305 <= $unsigned(($unsigned({reg1264}) != {reg1271}));
                      reg1306 <= $unsigned((8'hba));
                    end
                  else
                    begin
                      reg1304 <= ({(^$unsigned(forvar1299))} && reg1296);
                      reg1305 <= ($unsigned(((reg1302 ? (8'ha5) : forvar1271) ?
                              forvar1270 : $unsigned(reg1273))) ?
                          $unsigned(reg1257) : (+((~^reg1300) >> {reg1263})));
                      reg1306 <= (8'h9e);
                    end
                end
            end
          else
            begin
              if ((~(^reg1295[(1'h0):(1'h0)])))
                begin
                  if ($unsigned(forvar1253[(1'h0):(1'h0)]))
                    begin
                      reg1287 <= (^~reg1257);
                      reg1288 <= (forvar1268[(3'h4):(3'h4)] >>> {(|(reg1287 || (8'ha9)))});
                      reg1289 <= $signed((-(^$unsigned(reg1285))));
                      reg1290 <= reg1264;
                    end
                  else
                    begin
                      reg1287 <= ((~|reg1298[(2'h3):(1'h1)]) ^~ $signed(reg1253));
                      reg1288 <= forvar1287[(3'h7):(1'h0)];
                      reg1289 <= {$signed((reg1262[(4'h8):(3'h7)] ^ reg1266[(1'h0):(1'h0)]))};
                      reg1290 <= $unsigned($signed(({(8'hb7)} * (reg1264 ?
                          (8'ha7) : forvar1264))));
                    end
                  if ($unsigned((reg1282 & $unsigned($signed(reg1284)))))
                    begin
                      reg1291 <= {$signed($signed($signed(reg1267)))};
                      reg1292 <= $unsigned((&({forvar1264} ^ (+reg1276))));
                      reg1293 <= reg1265;
                    end
                  else
                    begin
                      reg1291 <= reg1260;
                      reg1292 <= reg1270[(3'h4):(3'h4)];
                      reg1293 <= ($signed((&reg1271)) || ($signed(reg1266[(2'h2):(1'h1)]) ?
                          {reg1290} : reg1277));
                      reg1294 <= $signed((&$unsigned(forvar1266)));
                    end
                end
              else
                begin
                  for (forvar1287 = (1'h0); (forvar1287 < (2'h3)); forvar1287 = (forvar1287 + (1'h1)))
                    begin
                      reg1288 <= $unsigned($unsigned(forvar1257[(2'h3):(2'h2)]));
                      reg1289 <= reg1270[(1'h1):(1'h0)];
                      reg1290 <= ((~^reg1257[(3'h7):(3'h4)]) & (^((reg1271 << reg1288) ?
                          (forvar1278 && reg1295) : $unsigned(reg1253))));
                      reg1291 <= reg1287;
                    end
                  if (((!(^~$signed(reg1255))) ?
                      ((reg1249[(1'h1):(1'h0)] >>> (^~reg1283)) ^~ reg1259) : reg1259[(4'ha):(2'h2)]))
                    begin
                      reg1292 <= (forvar1299[(1'h1):(1'h0)] * ({(forvar1260 ?
                                  reg1277 : reg1265)} ?
                          $signed($signed(reg1253)) : $signed((reg1258 || forvar1253))));
                      reg1293 <= reg1267[(2'h3):(1'h0)];
                      reg1294 <= $signed((8'hb2));
                      reg1295 <= forvar1253[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg1292 <= (reg1280 << (((^~reg1252) ?
                              (reg1261 ^ reg1306) : (&(8'hac))) ?
                          $unsigned(forvar1254[(1'h1):(1'h0)]) : {$signed(forvar1254)}));
                      reg1293 <= $signed((reg1247[(2'h3):(1'h0)] ?
                          (^~(reg1273 ? reg1252 : (8'h9e))) : forvar1266));
                    end
                end
              if ((reg1274 ? reg1272[(1'h0):(1'h0)] : reg1271[(4'ha):(4'h8)]))
                begin
                  if ((reg1264[(3'h4):(1'h1)] ?
                      forvar1287 : (reg1254 ?
                          ((reg1263 ?
                              reg1292 : forvar1303) & reg1256[(4'h8):(2'h2)]) : (8'hb3))))
                    begin
                      reg1296 <= (+($unsigned(reg1298[(3'h4):(1'h0)]) && ($unsigned((8'ha3)) ?
                          (~^reg1278) : $unsigned(reg1278))));
                      reg1297 <= reg1298;
                      reg1298 <= ($signed({$signed((8'hb0))}) ?
                          $unsigned(forvar1299) : $signed((^(&(8'ha5)))));
                    end
                  else
                    begin
                      reg1296 <= $signed(reg1256);
                      reg1297 <= ($signed($unsigned(reg1304[(3'h6):(2'h3)])) < forvar1272[(3'h6):(1'h0)]);
                      reg1298 <= $signed(forvar1249[(3'h5):(2'h3)]);
                    end
                  for (forvar1299 = (1'h0); (forvar1299 < (2'h2)); forvar1299 = (forvar1299 + (1'h1)))
                    begin
                      reg1300 <= $signed($unsigned((~(reg1291 ?
                          reg1263 : forvar1287))));
                      reg1301 <= $signed(($signed(reg1301) < (reg1250[(4'hb):(3'h7)] ?
                          wire1243[(3'h4):(1'h1)] : (forvar1253 >> reg1288))));
                    end
                  if ($signed((reg1301[(2'h2):(2'h2)] ^ ({reg1305} ~^ (~&(8'haa))))))
                    begin
                      reg1302 <= $unsigned($unsigned({(reg1256 ?
                              reg1283 : wire1243)}));
                      reg1303 <= $unsigned(((reg1267[(1'h0):(1'h0)] ?
                              (~|(8'ha3)) : $signed(reg1257)) ?
                          $signed((reg1265 - reg1297)) : $signed({reg1249})));
                      reg1304 <= $unsigned(($unsigned(reg1257[(2'h2):(1'h0)]) ?
                          {$signed(forvar1269)} : (~^$unsigned(reg1286))));
                      reg1305 <= $signed((|(((8'ha1) ? reg1252 : reg1281) ?
                          $signed(forvar1268) : $signed(reg1252))));
                    end
                  else
                    begin
                      reg1302 <= forvar1268;
                      reg1303 <= ({{forvar1249}} != (!(&reg1269[(3'h6):(3'h6)])));
                    end
                  for (forvar1306 = (1'h0); (forvar1306 < (2'h2)); forvar1306 = (forvar1306 + (1'h1)))
                    begin
                      reg1307 <= (forvar1270 > forvar1303);
                      reg1308 <= forvar1253[(3'h6):(3'h6)];
                      reg1309 <= reg1289[(4'h8):(3'h5)];
                      reg1310 <= (!forvar1259[(3'h6):(2'h3)]);
                    end
                end
              else
                begin
                  if ($signed(({(reg1247 ?
                          wire1245 : reg1300)} >= ((!reg1278) ^ (forvar1253 ?
                      reg1263 : reg1274)))))
                    begin
                      reg1296 <= reg1292[(2'h3):(1'h1)];
                      reg1297 <= $unsigned($unsigned(((-forvar1303) ~^ $unsigned(forvar1264))));
                    end
                  else
                    begin
                      reg1296 <= $signed($signed({reg1296[(3'h6):(2'h2)]}));
                      reg1297 <= $signed(reg1265);
                      reg1298 <= (reg1276 ?
                          $unsigned($unsigned({(8'hb9)})) : (((reg1289 >> reg1272) >> $unsigned(forvar1264)) <= reg1307));
                      reg1299 <= $signed(reg1260[(4'hd):(4'hb)]);
                    end
                  if (wire1244[(3'h7):(3'h6)])
                    begin
                      reg1300 <= forvar1248;
                      reg1301 <= {forvar1266};
                    end
                  else
                    begin
                      reg1300 <= $unsigned(wire1244[(3'h5):(2'h2)]);
                      reg1301 <= $signed($unsigned(wire1243[(1'h0):(1'h0)]));
                      reg1302 <= {reg1249};
                      reg1303 <= $unsigned((forvar1259[(2'h3):(2'h3)] ?
                          $signed(reg1288[(2'h3):(2'h3)]) : (forvar1269[(3'h7):(1'h0)] ?
                              reg1253[(1'h1):(1'h0)] : (~forvar1282))));
                    end
                end
              for (forvar1311 = (1'h0); (forvar1311 < (1'h0)); forvar1311 = (forvar1311 + (1'h1)))
                begin
                  if ($unsigned(reg1295))
                    begin
                      reg1312 <= ((+(-forvar1293[(2'h2):(2'h2)])) ~^ forvar1259[(1'h0):(1'h0)]);
                      reg1313 <= reg1285[(4'ha):(2'h3)];
                      reg1314 <= ((~|($signed(reg1299) >= (reg1257 <= forvar1249))) ?
                          reg1256 : (^(~{reg1259})));
                      reg1315 <= ((reg1287 || $signed((forvar1259 >> reg1280))) - ((forvar1303 ~^ $unsigned((8'hb9))) ?
                          reg1249[(1'h0):(1'h0)] : $unsigned({forvar1275})));
                    end
                  else
                    begin
                      reg1312 <= $unsigned(((^~$signed(forvar1253)) ?
                          $unsigned($signed(forvar1299)) : (((8'hb4) ?
                              forvar1257 : reg1266) >>> forvar1270)));
                      reg1313 <= ((($signed(forvar1260) ?
                              reg1264[(1'h0):(1'h0)] : (|forvar1268)) ?
                          reg1266[(1'h0):(1'h0)] : $unsigned($unsigned(reg1271))) == $signed(($signed(reg1257) ?
                          (reg1314 ?
                              reg1265 : reg1272) : $signed(forvar1278))));
                    end
                  for (forvar1316 = (1'h0); (forvar1316 < (2'h3)); forvar1316 = (forvar1316 + (1'h1)))
                    begin
                      reg1317 <= ((($unsigned((8'hb2)) | reg1282) ?
                          $unsigned($signed(wire1245)) : reg1293[(3'h5):(3'h4)]) == ($signed($signed(reg1252)) && $unsigned((reg1307 ?
                          (8'h9f) : reg1271))));
                    end
                  for (forvar1318 = (1'h0); (forvar1318 < (2'h3)); forvar1318 = (forvar1318 + (1'h1)))
                    begin
                      reg1319 <= forvar1255;
                      reg1320 <= forvar1270;
                      reg1321 <= (~forvar1259[(3'h6):(3'h5)]);
                      reg1322 <= $unsigned(({$signed(reg1296)} * forvar1255[(2'h3):(2'h3)]));
                    end
                  reg1323 <= reg1312;
                end
            end
          reg1324 <= (+((&{(8'ha5)}) ?
              $signed((reg1284 ?
                  reg1260 : reg1273)) : forvar1259[(3'h6):(2'h2)]));
          if (($unsigned($unsigned((^~reg1265))) >> $unsigned(((reg1282 >> reg1303) && reg1262))))
            begin
              if ((((~forvar1268[(2'h2):(1'h0)]) <= {$signed(reg1277)}) ^ (8'h9d)))
                begin
                  if (reg1307)
                    begin
                      reg1325 <= {reg1258};
                      reg1326 <= reg1272[(2'h2):(2'h2)];
                      reg1327 <= ($unsigned(forvar1278) - ($signed(reg1284[(3'h5):(3'h5)]) ?
                          reg1306[(1'h1):(1'h1)] : $unsigned(forvar1249[(4'h8):(1'h1)])));
                    end
                  else
                    begin
                      reg1325 <= (|{(reg1314 ? reg1296 : $signed(reg1319))});
                      reg1326 <= (reg1287[(2'h2):(1'h1)] * (|$signed($signed(reg1258))));
                      reg1327 <= (8'ha4);
                    end
                  for (forvar1328 = (1'h0); (forvar1328 < (1'h1)); forvar1328 = (forvar1328 + (1'h1)))
                    begin
                      reg1329 <= reg1268;
                      reg1330 <= {reg1277[(1'h1):(1'h0)]};
                    end
                end
              else
                begin
                  if ((8'ha3))
                    begin
                      reg1325 <= $unsigned(($unsigned((reg1285 ?
                              reg1266 : forvar1254)) ?
                          (~&$unsigned((8'ha7))) : forvar1272));
                    end
                  else
                    begin
                      reg1325 <= $signed(($unsigned((reg1309 ^~ reg1276)) ?
                          $unsigned($signed(forvar1253)) : (^$signed(wire1246))));
                    end
                  reg1326 <= (((&((8'hb3) ? forvar1311 : reg1272)) ?
                          (~|{reg1288}) : reg1269[(3'h5):(1'h0)]) ?
                      {reg1252} : (forvar1293 ~^ reg1258[(4'h9):(3'h7)]));
                  reg1327 <= ($signed(reg1325) ?
                      reg1260 : $unsigned($unsigned({reg1310})));
                  if (($signed(reg1275[(1'h1):(1'h0)]) != (^(~|$signed(reg1307)))))
                    begin
                      reg1328 <= $unsigned(forvar1318[(2'h2):(1'h1)]);
                      reg1329 <= ($unsigned((~^$signed((8'hac)))) ?
                          {(~&(reg1261 == reg1285))} : (((forvar1272 >>> reg1329) <= (forvar1255 ?
                                  wire1245 : reg1310)) ?
                              $unsigned($unsigned(reg1271)) : {reg1273[(3'h4):(3'h4)]}));
                    end
                  else
                    begin
                      reg1328 <= ($signed(((reg1290 ? (8'hb1) : reg1297) ?
                              (&reg1309) : $signed(reg1282))) ?
                          (&reg1260) : ((!forvar1306) ?
                              $signed(reg1273[(3'h7):(3'h6)]) : ($unsigned(forvar1287) >> (reg1307 != reg1253))));
                      reg1329 <= ($signed({(reg1315 ?
                              reg1310 : reg1315)}) && $signed(((reg1280 ^ reg1280) <<< $signed(reg1330))));
                      reg1330 <= {(-($unsigned(reg1296) && wire1246[(2'h2):(1'h1)]))};
                    end
                end
              for (forvar1331 = (1'h0); (forvar1331 < (1'h1)); forvar1331 = (forvar1331 + (1'h1)))
                begin
                  if ((forvar1318 <= $signed(((~^reg1261) <<< $signed(forvar1306)))))
                    begin
                      reg1332 <= $unsigned($signed({{reg1271}}));
                      reg1333 <= reg1266;
                      reg1334 <= reg1283;
                      reg1335 <= {(8'ha5)};
                    end
                  else
                    begin
                      reg1332 <= {(^~reg1276[(2'h2):(1'h1)])};
                    end
                  reg1336 <= (8'hba);
                  if (reg1317)
                    begin
                      reg1337 <= (reg1304 ?
                          reg1261 : (((reg1313 ?
                                  reg1313 : reg1270) >>> (^reg1256)) ?
                              ({(8'ha4)} ?
                                  (reg1336 | forvar1248) : {reg1289}) : forvar1328));
                      reg1338 <= ((8'hb0) >> {$signed((8'ha5))});
                    end
                  else
                    begin
                      reg1337 <= reg1324;
                      reg1338 <= (~(($signed(forvar1311) ?
                          (^~reg1305) : reg1292[(1'h0):(1'h0)]) >>> reg1283));
                      reg1339 <= (reg1285[(3'h4):(2'h2)] < reg1336);
                    end
                end
              if ({($unsigned($signed(reg1327)) < {reg1263[(3'h4):(3'h4)]})})
                begin
                  for (forvar1340 = (1'h0); (forvar1340 < (2'h2)); forvar1340 = (forvar1340 + (1'h1)))
                    begin
                      reg1341 <= (forvar1259[(2'h2):(1'h0)] > $signed((^~(reg1285 & reg1335))));
                      reg1342 <= forvar1340[(3'h5):(2'h3)];
                      reg1343 <= {(~&(forvar1306[(4'ha):(3'h4)] ?
                              $unsigned((8'hb3)) : forvar1306[(4'hd):(3'h4)]))};
                    end
                  for (forvar1344 = (1'h0); (forvar1344 < (1'h0)); forvar1344 = (forvar1344 + (1'h1)))
                    begin
                      reg1345 <= $unsigned((~&$signed($signed(forvar1269))));
                      reg1346 <= (((8'ha7) ?
                          reg1249 : ((reg1265 - reg1278) ?
                              $signed(reg1314) : (^forvar1248))) <<< forvar1306[(4'hd):(4'ha)]);
                      reg1347 <= $signed($unsigned(forvar1260[(2'h2):(1'h0)]));
                      reg1348 <= (reg1317[(4'hd):(4'hd)] ?
                          {reg1260} : $unsigned({reg1313[(2'h2):(1'h0)]}));
                    end
                  for (forvar1349 = (1'h0); (forvar1349 < (1'h0)); forvar1349 = (forvar1349 + (1'h1)))
                    begin
                      reg1350 <= forvar1344[(2'h2):(2'h2)];
                    end
                  if (forvar1287[(2'h2):(1'h1)])
                    begin
                      reg1351 <= {(($unsigned((8'ha7)) ?
                              (reg1275 ?
                                  forvar1316 : reg1330) : $signed(reg1277)) <<< reg1325[(4'h9):(1'h0)])};
                      reg1352 <= (~((^~reg1272) ?
                          reg1290 : $unsigned((+reg1263))));
                    end
                  else
                    begin
                      reg1351 <= (^~$unsigned((8'hb1)));
                    end
                end
              else
                begin
                  for (forvar1340 = (1'h0); (forvar1340 < (1'h1)); forvar1340 = (forvar1340 + (1'h1)))
                    begin
                      reg1341 <= ((^$signed((reg1332 | reg1278))) == ($signed($unsigned(forvar1249)) ?
                          reg1277[(1'h0):(1'h0)] : {{reg1276}}));
                      reg1342 <= forvar1328;
                    end
                end
            end
          else
            begin
              for (forvar1325 = (1'h0); (forvar1325 < (1'h0)); forvar1325 = (forvar1325 + (1'h1)))
                begin
                  for (forvar1326 = (1'h0); (forvar1326 < (2'h3)); forvar1326 = (forvar1326 + (1'h1)))
                    begin
                      reg1327 <= $unsigned(((~(-forvar1316)) ?
                          (reg1343[(2'h3):(1'h0)] ?
                              (reg1333 & forvar1325) : {forvar1287}) : reg1257[(3'h5):(3'h4)]));
                    end
                  if ($signed(reg1348))
                    begin
                      reg1328 <= ((^~(+((8'ha8) ? forvar1255 : (8'hb7)))) ?
                          (forvar1270[(3'h4):(1'h1)] + forvar1306[(4'ha):(4'h9)]) : reg1269[(3'h7):(3'h6)]);
                      reg1329 <= reg1308[(4'hd):(4'h8)];
                    end
                  else
                    begin
                      reg1328 <= (reg1343 ?
                          ((~(!reg1303)) != (+reg1259)) : forvar1253);
                      reg1329 <= $signed((reg1314[(2'h2):(2'h2)] ^ forvar1325[(1'h0):(1'h0)]));
                      reg1330 <= ($unsigned($signed(reg1268[(3'h4):(2'h2)])) + reg1317[(3'h6):(3'h4)]);
                    end
                  reg1331 <= (^~$unsigned($signed((reg1293 ?
                      (8'ha3) : reg1272))));
                end
            end
        end
      reg1353 <= $unsigned(wire1243[(3'h6):(3'h4)]);
      reg1354 <= (((8'h9f) ?
          reg1294[(3'h7):(2'h3)] : reg1261[(2'h2):(2'h2)]) == (|(~|{wire1246})));
    end
  assign wire1355 = (~|(~^$unsigned(reg1320[(3'h7):(3'h5)])));
  always
    @(posedge clk) begin
      if (reg1266[(2'h2):(1'h1)])
        begin
          for (forvar1356 = (1'h0); (forvar1356 < (2'h3)); forvar1356 = (forvar1356 + (1'h1)))
            begin
              for (forvar1357 = (1'h0); (forvar1357 < (2'h3)); forvar1357 = (forvar1357 + (1'h1)))
                begin
                  for (forvar1358 = (1'h0); (forvar1358 < (2'h2)); forvar1358 = (forvar1358 + (1'h1)))
                    begin
                      reg1359 <= reg1286[(3'h5):(2'h2)];
                      reg1360 <= (reg1303[(3'h4):(3'h4)] ?
                          (((reg1335 ? (8'hb5) : reg1278) ?
                                  {(8'h9f)} : $unsigned(reg1276)) ?
                              reg1288 : ({(8'ha8)} || (reg1279 ?
                                  (8'ha5) : reg1317))) : wire1243[(4'ha):(3'h7)]);
                      reg1361 <= reg1325[(1'h1):(1'h1)];
                      reg1362 <= {$unsigned(($signed((8'hb6)) ?
                              $signed(reg1258) : $signed(reg1343)))};
                    end
                  for (forvar1363 = (1'h0); (forvar1363 < (2'h3)); forvar1363 = (forvar1363 + (1'h1)))
                    begin
                      reg1364 <= $signed(reg1283[(4'ha):(3'h7)]);
                      reg1365 <= reg1309[(3'h5):(2'h2)];
                    end
                  for (forvar1366 = (1'h0); (forvar1366 < (1'h0)); forvar1366 = (forvar1366 + (1'h1)))
                    begin
                      reg1367 <= reg1247[(2'h3):(1'h0)];
                      reg1368 <= reg1338[(3'h6):(2'h3)];
                    end
                end
              for (forvar1369 = (1'h0); (forvar1369 < (2'h3)); forvar1369 = (forvar1369 + (1'h1)))
                begin
                  if ((8'h9c))
                    begin
                      reg1370 <= $unsigned(reg1266);
                      reg1371 <= reg1330[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1370 <= reg1297[(3'h4):(1'h1)];
                      reg1371 <= reg1269[(2'h2):(2'h2)];
                    end
                end
              for (forvar1372 = (1'h0); (forvar1372 < (1'h0)); forvar1372 = (forvar1372 + (1'h1)))
                begin
                  for (forvar1373 = (1'h0); (forvar1373 < (2'h3)); forvar1373 = (forvar1373 + (1'h1)))
                    begin
                      reg1374 <= reg1303;
                      reg1375 <= $signed((-$unsigned(reg1285)));
                      reg1376 <= ((~^(reg1306 ?
                              reg1299[(4'hc):(4'hc)] : reg1317[(4'h8):(2'h2)])) ?
                          reg1254 : $signed(wire1243[(1'h0):(1'h0)]));
                    end
                end
            end
          if ((^{reg1293}))
            begin
              reg1377 <= reg1309[(4'h9):(2'h2)];
            end
          else
            begin
              if (reg1266)
                begin
                  reg1377 <= $unsigned($unsigned((reg1345[(1'h1):(1'h1)] != {(8'ha4)})));
                  reg1378 <= $unsigned((~$unsigned(reg1255[(1'h0):(1'h0)])));
                  for (forvar1379 = (1'h0); (forvar1379 < (1'h0)); forvar1379 = (forvar1379 + (1'h1)))
                    begin
                      reg1380 <= reg1259[(3'h7):(2'h3)];
                      reg1381 <= reg1375;
                    end
                  if ($unsigned($signed(((reg1279 ?
                      reg1268 : reg1261) ^ (reg1276 ? reg1312 : reg1299)))))
                    begin
                      reg1382 <= reg1359;
                    end
                  else
                    begin
                      reg1382 <= (8'h9c);
                      reg1383 <= {reg1354};
                    end
                end
              else
                begin
                  for (forvar1377 = (1'h0); (forvar1377 < (2'h3)); forvar1377 = (forvar1377 + (1'h1)))
                    begin
                      reg1378 <= ($unsigned($unsigned(reg1352)) + wire1355[(1'h1):(1'h1)]);
                      reg1379 <= (+forvar1373[(3'h7):(3'h6)]);
                    end
                end
              if (forvar1373)
                begin
                  for (forvar1384 = (1'h0); (forvar1384 < (1'h0)); forvar1384 = (forvar1384 + (1'h1)))
                    begin
                      reg1385 <= $signed($signed(((+reg1321) >> $unsigned((8'h9f)))));
                      reg1386 <= $unsigned($unsigned(($unsigned(forvar1369) ?
                          (!reg1375) : (-reg1325))));
                      reg1387 <= reg1333;
                    end
                  for (forvar1388 = (1'h0); (forvar1388 < (1'h0)); forvar1388 = (forvar1388 + (1'h1)))
                    begin
                      reg1389 <= (reg1336[(3'h7):(3'h7)] > {(&reg1247)});
                      reg1390 <= {(reg1278 * (-(reg1362 ? reg1272 : reg1365)))};
                      reg1391 <= reg1301[(2'h3):(2'h2)];
                      reg1392 <= {(+(8'ha3))};
                    end
                  reg1393 <= forvar1373[(4'hb):(2'h3)];
                end
              else
                begin
                  if (($unsigned(($unsigned((8'hb2)) >= reg1380)) > reg1312))
                    begin
                      reg1384 <= {(reg1312 ~^ $unsigned((wire1355 ?
                              reg1392 : reg1264)))};
                      reg1385 <= $signed($signed({$unsigned(reg1341)}));
                      reg1386 <= $signed(reg1300);
                    end
                  else
                    begin
                      reg1384 <= ((($signed(reg1268) + reg1296) <<< $unsigned({reg1387})) << {$signed($signed(reg1371))});
                      reg1385 <= {forvar1369};
                      reg1386 <= $signed($unsigned((reg1324[(4'hb):(3'h7)] ?
                          reg1374[(2'h2):(2'h2)] : (~&reg1283))));
                    end
                end
            end
          reg1394 <= reg1277[(3'h4):(2'h2)];
          if ((8'h9c))
            begin
              if (((reg1273 - (|(^~reg1261))) ?
                  $signed(reg1281[(1'h0):(1'h0)]) : (&$signed((-reg1336)))))
                begin
                  for (forvar1395 = (1'h0); (forvar1395 < (1'h1)); forvar1395 = (forvar1395 + (1'h1)))
                    begin
                      reg1396 <= ($signed($signed((reg1345 ?
                              reg1323 : reg1251))) ?
                          $signed(($signed((8'hb2)) || $unsigned((8'haf)))) : {reg1321[(4'ha):(3'h7)]});
                      reg1397 <= $signed(reg1277[(3'h6):(3'h5)]);
                      reg1398 <= ((8'hb2) ?
                          forvar1357[(1'h0):(1'h0)] : ($signed($unsigned((8'ha2))) ?
                              (|((8'hb7) <<< (8'ha6))) : (reg1337 << reg1284[(1'h1):(1'h1)])));
                    end
                  for (forvar1399 = (1'h0); (forvar1399 < (1'h0)); forvar1399 = (forvar1399 + (1'h1)))
                    begin
                      reg1400 <= (8'haa);
                      reg1401 <= ($signed(forvar1363[(1'h0):(1'h0)]) ?
                          $signed(((reg1345 ?
                              (8'h9e) : reg1330) ~^ $signed(reg1387))) : reg1264[(1'h1):(1'h1)]);
                      reg1402 <= $signed((wire1355[(3'h6):(3'h4)] ?
                          reg1396 : reg1322[(1'h1):(1'h0)]));
                      reg1403 <= $signed($unsigned($unsigned(reg1264)));
                    end
                  for (forvar1404 = (1'h0); (forvar1404 < (2'h3)); forvar1404 = (forvar1404 + (1'h1)))
                    begin
                      reg1405 <= $signed((forvar1395 ~^ $signed(reg1337[(3'h4):(1'h1)])));
                      reg1406 <= ((&(+reg1308)) > $signed(reg1352[(3'h5):(3'h5)]));
                      reg1407 <= ({((reg1247 << reg1314) ~^ $unsigned(reg1376))} ^ $unsigned($unsigned((8'h9c))));
                    end
                end
              else
                begin
                  reg1395 <= {(-forvar1366[(2'h3):(1'h0)])};
                end
              reg1408 <= reg1385[(1'h1):(1'h1)];
            end
          else
            begin
              for (forvar1395 = (1'h0); (forvar1395 < (2'h3)); forvar1395 = (forvar1395 + (1'h1)))
                begin
                  if (reg1313)
                    begin
                      reg1396 <= ($unsigned(($unsigned(wire1246) ~^ $unsigned(reg1254))) < $unsigned(reg1379));
                    end
                  else
                    begin
                      reg1396 <= $signed($unsigned($unsigned((8'hb3))));
                      reg1397 <= {(~^$signed(((8'ha0) ?
                              wire1244 : forvar1358)))};
                    end
                end
              if (reg1320)
                begin
                  for (forvar1398 = (1'h0); (forvar1398 < (2'h3)); forvar1398 = (forvar1398 + (1'h1)))
                    begin
                      reg1399 <= reg1354;
                    end
                  reg1400 <= $signed(forvar1388[(1'h0):(1'h0)]);
                end
              else
                begin
                  reg1398 <= (8'hb7);
                  reg1399 <= reg1334[(3'h5):(2'h2)];
                end
              reg1401 <= {(((|reg1354) | {(8'ha0)}) ?
                      ({(8'ha1)} & reg1331[(2'h3):(1'h1)]) : reg1283[(4'hc):(4'hc)])};
              for (forvar1402 = (1'h0); (forvar1402 < (2'h2)); forvar1402 = (forvar1402 + (1'h1)))
                begin
                  for (forvar1403 = (1'h0); (forvar1403 < (1'h1)); forvar1403 = (forvar1403 + (1'h1)))
                    begin
                      reg1404 <= (-($signed((&(8'ha8))) ?
                          $unsigned((8'hb2)) : $unsigned(((8'hb6) ?
                              reg1266 : reg1345))));
                      reg1405 <= $signed(((((8'hb8) ? reg1305 : (8'ha3)) ?
                              $unsigned(reg1268) : (+reg1377)) ?
                          {{(8'ha1)}} : (reg1291 > (reg1262 ?
                              (8'ha4) : (8'hb7)))));
                      reg1406 <= ((^~{$unsigned(reg1352)}) >>> reg1250[(1'h0):(1'h0)]);
                      reg1407 <= (reg1375 ?
                          (&reg1329) : (((reg1259 ? reg1351 : reg1343) ?
                                  (~|reg1309) : reg1274) ?
                              $signed(reg1353) : $signed((-reg1247))));
                    end
                  reg1408 <= (8'hba);
                end
            end
        end
      else
        begin
          if (reg1330)
            begin
              if ($unsigned($unsigned((~|(^~reg1315)))))
                begin
                  for (forvar1356 = (1'h0); (forvar1356 < (1'h0)); forvar1356 = (forvar1356 + (1'h1)))
                    begin
                      reg1357 <= reg1375;
                    end
                  for (forvar1358 = (1'h0); (forvar1358 < (1'h1)); forvar1358 = (forvar1358 + (1'h1)))
                    begin
                      reg1359 <= ((^~$unsigned((8'hae))) >> (reg1361[(4'he):(1'h1)] ?
                          $signed(((8'hab) >> reg1291)) : $signed(reg1257[(4'hb):(3'h4)])));
                    end
                  for (forvar1360 = (1'h0); (forvar1360 < (2'h2)); forvar1360 = (forvar1360 + (1'h1)))
                    begin
                      reg1361 <= (~reg1361[(1'h1):(1'h1)]);
                    end
                  reg1362 <= (^~forvar1399[(2'h2):(1'h0)]);
                end
              else
                begin
                  if ($signed((reg1360 ?
                      {forvar1379} : ($signed(forvar1403) ?
                          ((8'hb9) - reg1315) : $signed(reg1330)))))
                    begin
                      reg1356 <= (forvar1384[(4'he):(3'h5)] ?
                          (($unsigned(reg1317) ?
                              reg1325[(3'h6):(3'h5)] : (reg1405 ?
                                  reg1379 : reg1251)) ^~ $unsigned({reg1333})) : ({$unsigned(reg1357)} ?
                              $signed(forvar1369) : reg1264));
                      reg1357 <= {$unsigned(reg1273[(3'h7):(1'h0)])};
                      reg1358 <= (~^{$unsigned(reg1402[(3'h7):(3'h4)])});
                      reg1359 <= (|reg1331[(3'h5):(3'h4)]);
                    end
                  else
                    begin
                      reg1356 <= (reg1406 ~^ (-reg1250));
                    end
                  if ({($unsigned((reg1264 >>> reg1293)) <= (reg1330[(2'h3):(2'h2)] ^~ $unsigned((8'ha5))))})
                    begin
                      reg1360 <= forvar1403[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1360 <= ($signed($unsigned((~&(8'hb7)))) - (~&(8'ha0)));
                    end
                end
            end
          else
            begin
              for (forvar1356 = (1'h0); (forvar1356 < (2'h2)); forvar1356 = (forvar1356 + (1'h1)))
                begin
                  reg1357 <= reg1350[(2'h2):(2'h2)];
                  for (forvar1358 = (1'h0); (forvar1358 < (2'h3)); forvar1358 = (forvar1358 + (1'h1)))
                    begin
                      reg1359 <= (reg1358 ?
                          $signed(reg1403[(3'h6):(3'h5)]) : ((((8'hb3) <<< reg1326) ?
                                  $unsigned(reg1408) : (reg1300 != (8'hb6))) ?
                              $signed($unsigned(reg1408)) : $signed((reg1315 <<< reg1288))));
                      reg1360 <= reg1402[(2'h2):(1'h1)];
                      reg1361 <= ($unsigned((~^$unsigned(reg1404))) >= reg1346);
                      reg1362 <= $unsigned((8'h9c));
                    end
                  for (forvar1363 = (1'h0); (forvar1363 < (2'h2)); forvar1363 = (forvar1363 + (1'h1)))
                    begin
                      reg1364 <= reg1298;
                      reg1365 <= forvar1398;
                      reg1366 <= $unsigned(reg1262[(4'hb):(1'h1)]);
                    end
                  for (forvar1367 = (1'h0); (forvar1367 < (2'h3)); forvar1367 = (forvar1367 + (1'h1)))
                    begin
                      reg1368 <= (($signed($signed(reg1395)) + reg1263) ?
                          (((forvar1367 ?
                              reg1371 : reg1362) + $signed(reg1271)) > ($unsigned(reg1382) ?
                              (reg1336 >> (8'ha6)) : (reg1247 >> reg1258))) : (((~reg1359) ?
                                  {reg1358} : (+reg1352)) ?
                              ($unsigned(reg1307) ?
                                  (reg1327 ?
                                      reg1280 : reg1337) : $unsigned(reg1305)) : (^~$signed((8'had)))));
                      reg1369 <= (((reg1353[(3'h6):(1'h1)] ?
                          $signed(reg1377) : (^(8'ha0))) & reg1345[(1'h1):(1'h1)]) << (((8'hab) == (wire1243 ?
                              reg1292 : reg1293)) ?
                          (~&(8'hab)) : {(reg1327 ? reg1287 : (8'hb1))}));
                    end
                end
              if (reg1326)
                begin
                  reg1370 <= ((((8'hb5) && (reg1342 * reg1257)) < $unsigned((|(8'ha4)))) ?
                      $unsigned((~|(reg1329 * (8'ha6)))) : ({(+reg1269)} >>> (8'haa)));
                  for (forvar1371 = (1'h0); (forvar1371 < (2'h3)); forvar1371 = (forvar1371 + (1'h1)))
                    begin
                      reg1372 <= reg1298;
                    end
                  if (reg1365)
                    begin
                      reg1373 <= ({$signed((reg1366 ?
                              reg1281 : reg1282))} ^ $unsigned((reg1268[(2'h2):(1'h1)] ?
                          {reg1353} : {reg1308})));
                    end
                  else
                    begin
                      reg1373 <= $unsigned((reg1259[(3'h6):(2'h3)] > $signed(reg1266[(1'h1):(1'h0)])));
                      reg1374 <= $unsigned($signed(reg1271[(3'h4):(3'h4)]));
                    end
                end
              else
                begin
                  for (forvar1370 = (1'h0); (forvar1370 < (1'h1)); forvar1370 = (forvar1370 + (1'h1)))
                    begin
                      reg1371 <= forvar1372;
                      reg1372 <= wire1244[(2'h3):(2'h3)];
                      reg1373 <= (reg1356 ?
                          reg1293 : ($signed((8'ha2)) >>> $signed(reg1301[(2'h3):(1'h1)])));
                      reg1374 <= (^~reg1301);
                    end
                  for (forvar1375 = (1'h0); (forvar1375 < (2'h2)); forvar1375 = (forvar1375 + (1'h1)))
                    begin
                      reg1376 <= ($unsigned($signed(reg1283[(3'h7):(2'h2)])) > (+$unsigned(forvar1402)));
                    end
                  reg1377 <= ({reg1315} && reg1348[(4'ha):(1'h1)]);
                end
            end
          for (forvar1378 = (1'h0); (forvar1378 < (2'h3)); forvar1378 = (forvar1378 + (1'h1)))
            begin
              for (forvar1379 = (1'h0); (forvar1379 < (2'h2)); forvar1379 = (forvar1379 + (1'h1)))
                begin
                  for (forvar1380 = (1'h0); (forvar1380 < (2'h3)); forvar1380 = (forvar1380 + (1'h1)))
                    begin
                      reg1381 <= {forvar1360};
                      reg1382 <= {reg1304};
                      reg1383 <= reg1345;
                    end
                  reg1384 <= ($unsigned(($unsigned(reg1314) ?
                          reg1287[(2'h2):(1'h0)] : reg1348)) ?
                      reg1343[(1'h0):(1'h0)] : (reg1303[(1'h0):(1'h0)] ?
                          forvar1371[(1'h1):(1'h1)] : $unsigned(reg1247[(2'h2):(1'h0)])));
                  reg1385 <= reg1288[(4'hc):(3'h6)];
                end
              for (forvar1386 = (1'h0); (forvar1386 < (1'h0)); forvar1386 = (forvar1386 + (1'h1)))
                begin
                  for (forvar1387 = (1'h0); (forvar1387 < (2'h3)); forvar1387 = (forvar1387 + (1'h1)))
                    begin
                      reg1388 <= forvar1378;
                      reg1389 <= reg1374;
                      reg1390 <= ({($signed(reg1273) != (reg1265 - reg1397))} ?
                          {$signed((reg1377 && reg1273))} : (((^(8'ha4)) ?
                              (8'h9c) : (reg1303 | reg1297)) && $unsigned(((8'ha8) >>> (8'ha8)))));
                    end
                end
            end
        end
    end
  assign wire1409 = {($signed(reg1252) ? reg1397[(4'hf):(4'he)] : reg1317)};
  assign wire1410 = {reg1395[(4'hb):(3'h7)]};
  module1411 #() modinst2587 (wire2586, clk, reg1360, reg1266, reg1267, reg1388);
  always
    @(posedge clk) begin
      for (forvar2588 = (1'h0); (forvar2588 < (2'h3)); forvar2588 = (forvar2588 + (1'h1)))
        begin
          for (forvar2589 = (1'h0); (forvar2589 < (2'h2)); forvar2589 = (forvar2589 + (1'h1)))
            begin
              if ($signed((+reg1332)))
                begin
                  if ((!$signed((~forvar2589[(3'h7):(3'h7)]))))
                    begin
                      reg2590 <= {($signed({reg1320}) ?
                              ((reg1336 && reg1341) ?
                                  reg1290[(4'hd):(2'h3)] : ((8'hae) <= reg1293)) : $signed($signed(wire1410)))};
                    end
                  else
                    begin
                      reg2590 <= $signed((8'h9d));
                      reg2591 <= ((reg1397 >> (&reg1303[(2'h2):(1'h0)])) ?
                          {(~^(~reg1378))} : $unsigned($unsigned(reg1336)));
                    end
                  for (forvar2592 = (1'h0); (forvar2592 < (2'h2)); forvar2592 = (forvar2592 + (1'h1)))
                    begin
                      reg2593 <= (~^(^~wire1243[(4'h9):(3'h4)]));
                    end
                  for (forvar2594 = (1'h0); (forvar2594 < (1'h0)); forvar2594 = (forvar2594 + (1'h1)))
                    begin
                      reg2595 <= reg1331[(1'h0):(1'h0)];
                    end
                  for (forvar2596 = (1'h0); (forvar2596 < (2'h2)); forvar2596 = (forvar2596 + (1'h1)))
                    begin
                      reg2597 <= $signed(reg1375);
                      reg2598 <= wire1244[(3'h4):(1'h1)];
                      reg2599 <= ((-($signed(reg1304) ?
                              (~reg2597) : (reg1302 ^ reg1404))) ?
                          forvar2596 : ($unsigned($unsigned(reg1346)) << ((reg1390 << (8'ha0)) == reg1250[(1'h1):(1'h0)])));
                      reg2600 <= ($signed($unsigned((reg2598 <= reg1277))) ?
                          $signed((((8'hb7) ~^ reg1385) ?
                              $unsigned(reg1325) : $signed(reg1394))) : (~{wire1246}));
                    end
                end
              else
                begin
                  for (forvar2590 = (1'h0); (forvar2590 < (2'h3)); forvar2590 = (forvar2590 + (1'h1)))
                    begin
                      reg2591 <= ($signed(reg1289[(4'hb):(1'h1)]) ?
                          reg1258[(1'h1):(1'h1)] : reg1375[(2'h2):(2'h2)]);
                      reg2592 <= $unsigned(((~|reg1282) ?
                          $unsigned((reg1406 ?
                              reg1255 : reg1303)) : $unsigned(((8'hae) ?
                              reg1400 : reg1390))));
                    end
                  for (forvar2593 = (1'h0); (forvar2593 < (2'h3)); forvar2593 = (forvar2593 + (1'h1)))
                    begin
                      reg2594 <= $signed(((~^$signed(reg1297)) - $unsigned({reg1370})));
                      reg2595 <= (forvar2596[(2'h2):(1'h1)] << forvar2593[(3'h7):(3'h7)]);
                    end
                  reg2596 <= ($unsigned($signed(reg1367[(2'h2):(1'h1)])) ?
                      ((+(^(8'hba))) ?
                          reg1366 : $signed($unsigned(reg1269))) : $signed(reg1256[(2'h3):(1'h0)]));
                end
              if ({($signed((^(8'h9e))) ?
                      (&(reg1327 > reg1356)) : ($unsigned(reg1327) ?
                          $signed(forvar2590) : (reg1403 ?
                              reg1259 : (8'ha9))))})
                begin
                  if ($signed({reg1395[(4'hb):(4'h9)]}))
                    begin
                      reg2601 <= (|$unsigned($unsigned((&reg1406))));
                      reg2602 <= (~^(~&((~^(8'ha9)) ?
                          (reg2597 <<< reg2598) : $unsigned((8'ha0)))));
                      reg2603 <= ((reg1304 ?
                          $unsigned((reg1368 ~^ reg1385)) : {(~^reg1283)}) && ($unsigned($signed(reg1297)) ?
                          reg1304 : (~^reg1299[(4'hc):(4'hb)])));
                      reg2604 <= reg1326;
                    end
                  else
                    begin
                      reg2601 <= $unsigned((($signed(wire1243) ?
                              (^reg1353) : (&reg1328)) ?
                          ((~reg1253) * reg2599) : (((8'hb3) >= reg1257) ?
                              reg1371[(1'h1):(1'h0)] : $unsigned(reg2602))));
                      reg2602 <= reg1348[(4'h8):(2'h3)];
                      reg2603 <= ((!reg1278) + $signed(reg1295));
                      reg2604 <= reg1375;
                    end
                  if (reg1293)
                    begin
                      reg2605 <= reg1290[(4'hb):(3'h6)];
                      reg2606 <= $unsigned(((~|reg1277) ?
                          ($unsigned(reg1350) ?
                              reg1370[(3'h4):(2'h3)] : (&(8'hac))) : $signed((~&reg1301))));
                      reg2607 <= (($unsigned((|reg1301)) ?
                          {(reg1306 ?
                                  wire1245 : reg1261)} : reg1393) - (~|{$signed(reg1275)}));
                    end
                  else
                    begin
                      reg2605 <= $unsigned($unsigned(({reg2594} ^ {(8'haf)})));
                      reg2606 <= reg2603;
                    end
                  for (forvar2608 = (1'h0); (forvar2608 < (1'h1)); forvar2608 = (forvar2608 + (1'h1)))
                    begin
                      reg2609 <= $unsigned($signed(((wire1409 < reg2591) & (8'hba))));
                      reg2610 <= reg1364;
                      reg2611 <= reg1276[(4'h8):(3'h5)];
                    end
                  reg2612 <= $signed($unsigned($signed($unsigned(reg1385))));
                end
              else
                begin
                  reg2601 <= (+reg1375[(2'h2):(2'h2)]);
                  for (forvar2602 = (1'h0); (forvar2602 < (2'h2)); forvar2602 = (forvar2602 + (1'h1)))
                    begin
                      reg2603 <= $unsigned(reg1314[(2'h2):(1'h0)]);
                    end
                end
            end
          if (reg2594[(1'h0):(1'h0)])
            begin
              for (forvar2613 = (1'h0); (forvar2613 < (2'h2)); forvar2613 = (forvar2613 + (1'h1)))
                begin
                  if ((~&($signed(reg1261[(4'hd):(4'h9)]) <= reg1365)))
                    begin
                      reg2614 <= $unsigned($unsigned({$unsigned(reg1290)}));
                      reg2615 <= reg1373[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg2614 <= (($unsigned((reg1307 ? reg1249 : reg1358)) ?
                              (8'hb2) : reg1366[(2'h3):(1'h1)]) ?
                          $signed(reg1398[(2'h2):(1'h0)]) : ((reg1306 ?
                                  $signed(reg1379) : reg1290[(3'h6):(1'h0)]) ?
                              reg1337 : (reg1348 <<< {reg1364})));
                      reg2615 <= (reg1405[(3'h5):(3'h5)] ?
                          $unsigned(reg1371[(1'h1):(1'h0)]) : ((reg1259[(3'h7):(3'h6)] < reg1347) ?
                              $signed(reg1272[(2'h2):(2'h2)]) : $signed(((8'haf) ?
                                  (8'ha3) : (8'hab)))));
                    end
                  for (forvar2616 = (1'h0); (forvar2616 < (2'h2)); forvar2616 = (forvar2616 + (1'h1)))
                    begin
                      reg2617 <= $signed($unsigned(reg1359[(3'h4):(3'h4)]));
                      reg2618 <= $unsigned((($signed(reg1371) ?
                          reg1397[(3'h5):(2'h3)] : {reg1288}) >> ((reg2595 ^~ wire1243) << $signed((8'haf)))));
                      reg2619 <= (-(8'hb6));
                    end
                  if (($signed(($unsigned(forvar2608) - reg1387)) ?
                      reg1250 : ((~&(reg1378 ?
                          reg1348 : reg1328)) <<< (^~(reg1293 + wire1409)))))
                    begin
                      reg2620 <= {{(^{forvar2596})}};
                      reg2621 <= reg1309[(4'hd):(1'h0)];
                      reg2622 <= {forvar2592[(1'h1):(1'h1)]};
                    end
                  else
                    begin
                      reg2620 <= {($unsigned($unsigned((8'ha3))) ~^ reg1342[(2'h2):(1'h1)])};
                      reg2621 <= $unsigned((reg2615 ?
                          (+$signed(reg2612)) : (reg1379[(4'hc):(4'h9)] ?
                              (forvar2593 ?
                                  reg1257 : (8'ha8)) : reg1343[(1'h0):(1'h0)])));
                      reg2622 <= $unsigned($unsigned(((reg1359 << reg1295) ?
                          {reg1372} : (reg1347 <<< reg1273))));
                      reg2623 <= reg1332[(1'h1):(1'h0)];
                    end
                  reg2624 <= reg2594;
                end
              reg2625 <= ($signed(reg1360) ?
                  $unsigned((|reg1396[(1'h1):(1'h1)])) : $unsigned({(-(8'ha7))}));
              for (forvar2626 = (1'h0); (forvar2626 < (1'h0)); forvar2626 = (forvar2626 + (1'h1)))
                begin
                  for (forvar2627 = (1'h0); (forvar2627 < (1'h0)); forvar2627 = (forvar2627 + (1'h1)))
                    begin
                      reg2628 <= (+{reg1367});
                    end
                end
              if ($unsigned(reg1295))
                begin
                  for (forvar2629 = (1'h0); (forvar2629 < (1'h0)); forvar2629 = (forvar2629 + (1'h1)))
                    begin
                      reg2630 <= ((!(reg1319[(1'h0):(1'h0)] ?
                              {reg1329} : {reg1249})) ?
                          forvar2589[(3'h5):(1'h1)] : $unsigned($unsigned(reg1276)));
                      reg2631 <= ((~|$unsigned(((8'hb2) ?
                              reg1362 : wire1355))) ?
                          reg1389[(3'h7):(1'h0)] : $signed(reg2593));
                      reg2632 <= $unsigned((reg1293 & ((reg1374 ?
                          reg2603 : reg2625) >> reg1308)));
                    end
                end
              else
                begin
                  for (forvar2629 = (1'h0); (forvar2629 < (2'h3)); forvar2629 = (forvar2629 + (1'h1)))
                    begin
                      reg2630 <= $unsigned($signed($signed(reg1335)));
                      reg2631 <= reg1322[(3'h6):(2'h3)];
                    end
                end
            end
          else
            begin
              for (forvar2613 = (1'h0); (forvar2613 < (1'h1)); forvar2613 = (forvar2613 + (1'h1)))
                begin
                  for (forvar2614 = (1'h0); (forvar2614 < (1'h0)); forvar2614 = (forvar2614 + (1'h1)))
                    begin
                      reg2615 <= ((^~({reg1352} || (reg2603 * reg1252))) <<< {(~reg2594[(3'h4):(1'h0)])});
                    end
                  if (({{reg1383[(3'h4):(2'h3)]}} <<< $signed($unsigned((reg1258 ^~ reg1297)))))
                    begin
                      reg2616 <= $unsigned($unsigned(reg1301[(1'h0):(1'h0)]));
                      reg2617 <= (reg1352 ?
                          $unsigned({((8'hb6) >= (8'had))}) : forvar2594);
                    end
                  else
                    begin
                      reg2616 <= $signed(reg1260);
                      reg2617 <= (!$signed((reg1269[(2'h2):(1'h1)] && $signed((8'hb9)))));
                      reg2618 <= (~^$signed(reg2617[(2'h2):(1'h0)]));
                    end
                end
            end
          reg2633 <= $signed($unsigned(reg1388));
          reg2634 <= reg1342;
        end
      for (forvar2635 = (1'h0); (forvar2635 < (1'h1)); forvar2635 = (forvar2635 + (1'h1)))
        begin
          reg2636 <= ((^~$signed(reg1347)) == $unsigned((-(reg1405 ?
              reg1268 : (8'hb8)))));
          reg2637 <= reg1297[(4'h8):(3'h4)];
        end
    end
  assign wire2638 = reg2619;
  always
    @(posedge clk) begin
      for (forvar2639 = (1'h0); (forvar2639 < (2'h3)); forvar2639 = (forvar2639 + (1'h1)))
        begin
          for (forvar2640 = (1'h0); (forvar2640 < (1'h0)); forvar2640 = (forvar2640 + (1'h1)))
            begin
              for (forvar2641 = (1'h0); (forvar2641 < (1'h0)); forvar2641 = (forvar2641 + (1'h1)))
                begin
                  for (forvar2642 = (1'h0); (forvar2642 < (2'h2)); forvar2642 = (forvar2642 + (1'h1)))
                    begin
                      reg2643 <= reg1406[(4'hb):(1'h1)];
                      reg2644 <= {$unsigned((~&$signed(reg1345)))};
                    end
                  for (forvar2645 = (1'h0); (forvar2645 < (1'h1)); forvar2645 = (forvar2645 + (1'h1)))
                    begin
                      reg2646 <= (reg2602 != reg1393[(2'h2):(1'h0)]);
                      reg2647 <= $signed(reg1255[(1'h1):(1'h1)]);
                      reg2648 <= reg1369;
                      reg2649 <= (($signed($signed(reg1387)) ?
                          (~(reg2634 ? (8'hb5) : reg1377)) : (((8'h9d) ?
                                  (8'hb2) : (8'hb9)) ?
                              (reg1391 > reg1308) : reg2590)) == (reg1269[(3'h6):(2'h2)] >> (+(reg1402 ?
                          (8'hac) : reg1362))));
                    end
                  if (((|(^~(reg1327 ? reg1382 : reg1312))) ?
                      ((reg1291[(2'h2):(1'h1)] ? (~|reg1264) : {reg1389}) ?
                          $signed(reg1376[(1'h1):(1'h1)]) : (|reg1343)) : $signed(($unsigned(reg1291) ?
                          (reg2647 ? reg1253 : wire1355) : (reg1283 ?
                              reg1367 : reg1408)))))
                    begin
                      reg2650 <= ((($signed(reg1334) || $signed(reg1274)) && reg2620[(3'h5):(3'h5)]) ^~ reg1326);
                    end
                  else
                    begin
                      reg2650 <= reg1341;
                      reg2651 <= $unsigned((^~reg1347[(3'h6):(3'h6)]));
                    end
                end
            end
          for (forvar2652 = (1'h0); (forvar2652 < (1'h1)); forvar2652 = (forvar2652 + (1'h1)))
            begin
              for (forvar2653 = (1'h0); (forvar2653 < (2'h2)); forvar2653 = (forvar2653 + (1'h1)))
                begin
                  for (forvar2654 = (1'h0); (forvar2654 < (1'h1)); forvar2654 = (forvar2654 + (1'h1)))
                    begin
                      reg2655 <= (($signed((reg1267 < reg1389)) >>> {$unsigned(reg1390)}) >>> (($signed(reg1359) ^~ $unsigned(reg1345)) <<< $unsigned((^reg1314))));
                      reg2656 <= $unsigned((+reg2597[(2'h2):(1'h1)]));
                      reg2657 <= (reg2656 ?
                          {{$unsigned((8'hb7))}} : (~&((^~forvar2639) + {reg2611})));
                      reg2658 <= reg1377[(3'h4):(3'h4)];
                    end
                  reg2659 <= (!($unsigned(reg1249) ?
                      {reg2602} : $signed(reg1257)));
                  reg2660 <= $unsigned(reg1312[(3'h6):(3'h4)]);
                end
              if ((reg1403 ^ reg1259[(3'h5):(1'h0)]))
                begin
                  for (forvar2661 = (1'h0); (forvar2661 < (2'h3)); forvar2661 = (forvar2661 + (1'h1)))
                    begin
                      reg2662 <= (-$signed(({reg2643} ?
                          $signed((8'haa)) : (^(8'hb7)))));
                      reg2663 <= $unsigned((&($unsigned(reg1259) ^ $unsigned(reg1269))));
                      reg2664 <= (reg1330 ?
                          $unsigned($unsigned((reg1309 >> reg2607))) : (+(reg2593[(3'h6):(3'h4)] ?
                              reg2647[(1'h0):(1'h0)] : $unsigned(reg2602))));
                      reg2665 <= {reg1335};
                    end
                  for (forvar2666 = (1'h0); (forvar2666 < (2'h2)); forvar2666 = (forvar2666 + (1'h1)))
                    begin
                      reg2667 <= reg2591[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  reg2661 <= (((wire1246[(2'h3):(1'h0)] ?
                          (8'h9c) : (reg2660 ?
                              reg1346 : (8'haf))) >> ($unsigned(reg1284) ?
                          $signed(reg2663) : reg1342)) ?
                      reg1310 : ((~&(reg1317 ?
                          reg2655 : reg2594)) <<< {$signed(reg1251)}));
                  reg2662 <= (^reg1376[(1'h0):(1'h0)]);
                  for (forvar2663 = (1'h0); (forvar2663 < (1'h1)); forvar2663 = (forvar2663 + (1'h1)))
                    begin
                      reg2664 <= (~|(^~$unsigned((reg1366 ?
                          reg2614 : reg1328))));
                    end
                  if ((~$unsigned($unsigned($signed(reg2590)))))
                    begin
                      reg2665 <= $signed((reg1399 >> (&(reg2649 <= reg2628))));
                      reg2666 <= reg1352[(1'h1):(1'h1)];
                      reg2667 <= reg1321[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg2665 <= reg1366;
                    end
                end
            end
          for (forvar2668 = (1'h0); (forvar2668 < (2'h2)); forvar2668 = (forvar2668 + (1'h1)))
            begin
              for (forvar2669 = (1'h0); (forvar2669 < (2'h3)); forvar2669 = (forvar2669 + (1'h1)))
                begin
                  if (reg1400[(4'hc):(2'h3)])
                    begin
                      reg2670 <= reg1303;
                      reg2671 <= reg2632;
                      reg2672 <= $signed(reg1387[(1'h1):(1'h1)]);
                      reg2673 <= ((({reg1327} ?
                          $signed(reg2633) : $signed(reg2593)) <<< reg1289) ^ reg1337);
                    end
                  else
                    begin
                      reg2670 <= reg1294[(4'ha):(2'h2)];
                      reg2671 <= $signed(($signed($unsigned(reg1333)) ?
                          reg1317 : (-(reg2665 ? reg1334 : reg1317))));
                      reg2672 <= reg1367;
                    end
                  if (reg2661[(1'h0):(1'h0)])
                    begin
                      reg2674 <= $signed((^~$unsigned($unsigned(reg1321))));
                      reg2675 <= reg2655[(3'h4):(2'h3)];
                      reg2676 <= ((~&$signed((8'ha5))) ~^ $unsigned({$unsigned(reg1404)}));
                      reg2677 <= $unsigned((((reg1308 ? reg1384 : reg1279) ?
                          (reg1390 <<< reg2599) : reg2598[(3'h4):(1'h1)]) && reg1326[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg2674 <= (~reg1339[(1'h1):(1'h1)]);
                      reg2675 <= reg1356;
                      reg2676 <= $signed({(reg1317 <<< $unsigned(reg1271))});
                    end
                  reg2678 <= reg1331[(2'h2):(1'h0)];
                  for (forvar2679 = (1'h0); (forvar2679 < (1'h0)); forvar2679 = (forvar2679 + (1'h1)))
                    begin
                      reg2680 <= $unsigned(($signed((wire1410 ?
                              (8'ha3) : wire1355)) ?
                          $signed((reg1345 <= reg1376)) : reg1299));
                    end
                end
              for (forvar2681 = (1'h0); (forvar2681 < (2'h2)); forvar2681 = (forvar2681 + (1'h1)))
                begin
                  if (($unsigned((reg2606 - reg1270)) && $unsigned((&wire1355[(2'h3):(1'h0)]))))
                    begin
                      reg2682 <= reg2620;
                      reg2683 <= ((~|$signed((forvar2639 && reg1293))) ?
                          (!{{(8'haa)}}) : $signed(reg1308[(3'h6):(1'h0)]));
                    end
                  else
                    begin
                      reg2682 <= $signed((((~reg1281) || reg2599) << (|reg1255[(3'h6):(2'h2)])));
                    end
                  for (forvar2684 = (1'h0); (forvar2684 < (1'h0)); forvar2684 = (forvar2684 + (1'h1)))
                    begin
                      reg2685 <= ({reg1406} ? reg1289[(3'h5):(1'h1)] : reg1301);
                      reg2686 <= reg1408;
                      reg2687 <= $signed(reg1304[(3'h5):(3'h4)]);
                    end
                end
              if ((8'hb3))
                begin
                  for (forvar2688 = (1'h0); (forvar2688 < (1'h0)); forvar2688 = (forvar2688 + (1'h1)))
                    begin
                      reg2689 <= ({((reg1249 ? forvar2681 : (8'hb0)) ?
                              (reg1386 ?
                                  reg1391 : (8'ha0)) : $unsigned(reg1283))} + ((&reg1322[(2'h2):(2'h2)]) - reg2593[(1'h0):(1'h0)]));
                      reg2690 <= ($signed(((reg1252 ? reg2619 : reg2599) ?
                              (reg1369 ?
                                  reg2670 : forvar2661) : $unsigned(reg2672))) ?
                          (|$signed(reg2597[(4'hb):(1'h0)])) : (($signed(reg1394) << (reg2591 ?
                                  reg1338 : reg1377)) ?
                              (8'had) : ({reg2673} << {reg2672})));
                      reg2691 <= reg1396;
                    end
                  for (forvar2692 = (1'h0); (forvar2692 < (2'h3)); forvar2692 = (forvar2692 + (1'h1)))
                    begin
                      reg2693 <= reg1377[(1'h1):(1'h0)];
                      reg2694 <= reg2643[(2'h2):(2'h2)];
                    end
                  reg2695 <= reg1270;
                end
              else
                begin
                  for (forvar2688 = (1'h0); (forvar2688 < (2'h2)); forvar2688 = (forvar2688 + (1'h1)))
                    begin
                      reg2689 <= (wire1410 <= (^~((reg2595 <<< (8'ha8)) ?
                          reg1263[(2'h3):(2'h2)] : ((8'hb9) ^~ reg1250))));
                    end
                end
              for (forvar2696 = (1'h0); (forvar2696 < (1'h0)); forvar2696 = (forvar2696 + (1'h1)))
                begin
                  for (forvar2697 = (1'h0); (forvar2697 < (2'h3)); forvar2697 = (forvar2697 + (1'h1)))
                    begin
                      reg2698 <= reg1400;
                      reg2699 <= wire1246[(2'h3):(2'h2)];
                    end
                  if ({$signed((~&(wire2586 ? reg2690 : reg2699)))})
                    begin
                      reg2700 <= reg1260;
                      reg2701 <= $signed((~^$unsigned(reg1301)));
                      reg2702 <= $unsigned(((-(reg1310 <= (8'ha8))) ?
                          (reg1386 | $unsigned((8'ha1))) : ({reg1270} ?
                              (~reg2611) : (^(8'hb7)))));
                    end
                  else
                    begin
                      reg2700 <= $unsigned(((~|reg1342[(3'h4):(3'h4)]) <= reg1247[(3'h6):(2'h2)]));
                      reg2701 <= $signed(reg2637[(2'h2):(1'h1)]);
                    end
                end
            end
        end
    end
  assign wire2703 = $signed(reg2601);
  assign wire2704 = reg1288;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1411  (y, clk, wire1412, wire1413, wire1414, wire1415);
  output wire [(32'h1ddd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire1412;
  input wire signed [(4'h9):(1'h0)] wire1413;
  input wire signed [(4'h8):(1'h0)] wire1414;
  input wire signed [(2'h2):(1'h0)] wire1415;
  wire signed [(3'h7):(1'h0)] wire2539;
  wire signed [(4'ha):(1'h0)] wire2331;
  wire signed [(4'ha):(1'h0)] wire2253;
  wire signed [(4'hd):(1'h0)] wire2252;
  wire signed [(3'h6):(1'h0)] wire2251;
  wire signed [(3'h6):(1'h0)] wire2250;
  wire [(2'h2):(1'h0)] wire2031;
  wire [(3'h6):(1'h0)] wire2030;
  wire [(2'h3):(1'h0)] wire2029;
  wire [(4'ha):(1'h0)] wire1416;
  wire signed [(3'h7):(1'h0)] wire2027;
  reg [(3'h6):(1'h0)] reg2540 = (1'h0);
  reg [(4'hf):(1'h0)] reg2584 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2580 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2577 = (1'h0);
  reg [(4'hf):(1'h0)] reg2585 = (1'h0);
  reg [(5'h10):(1'h0)] reg2583 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2582 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2581 = (1'h0);
  reg [(4'hb):(1'h0)] reg2578 = (1'h0);
  reg [(3'h4):(1'h0)] reg2576 = (1'h0);
  reg [(3'h6):(1'h0)] reg2575 = (1'h0);
  reg [(2'h2):(1'h0)] reg2574 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2573 = (1'h0);
  reg [(4'h9):(1'h0)] reg2572 = (1'h0);
  reg [(3'h7):(1'h0)] reg2571 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2570 = (1'h0);
  reg [(4'h9):(1'h0)] reg2569 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2568 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2567 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2566 = (1'h0);
  reg [(4'hd):(1'h0)] reg2565 = (1'h0);
  reg [(4'ha):(1'h0)] reg2564 = (1'h0);
  reg [(3'h6):(1'h0)] reg2563 = (1'h0);
  reg [(3'h6):(1'h0)] reg2562 = (1'h0);
  reg [(4'hb):(1'h0)] reg2561 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2560 = (1'h0);
  reg [(2'h3):(1'h0)] reg2558 = (1'h0);
  reg [(4'hc):(1'h0)] reg2557 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2555 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2554 = (1'h0);
  reg [(4'hb):(1'h0)] reg2553 = (1'h0);
  reg [(5'h10):(1'h0)] reg2552 = (1'h0);
  reg [(4'h9):(1'h0)] reg2551 = (1'h0);
  reg [(4'hb):(1'h0)] reg2549 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2548 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2547 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2546 = (1'h0);
  reg [(4'hb):(1'h0)] reg2544 = (1'h0);
  reg [(4'hc):(1'h0)] reg2541 = (1'h0);
  reg [(2'h2):(1'h0)] reg2538 = (1'h0);
  reg [(4'hb):(1'h0)] reg2537 = (1'h0);
  reg [(2'h3):(1'h0)] reg2536 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2534 = (1'h0);
  reg [(4'h8):(1'h0)] reg2533 = (1'h0);
  reg [(4'ha):(1'h0)] reg2532 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2531 = (1'h0);
  reg [(3'h5):(1'h0)] reg2520 = (1'h0);
  reg [(4'h8):(1'h0)] reg2529 = (1'h0);
  reg [(4'h8):(1'h0)] reg2528 = (1'h0);
  reg [(3'h4):(1'h0)] reg2527 = (1'h0);
  reg [(4'h8):(1'h0)] reg2526 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2525 = (1'h0);
  reg [(3'h5):(1'h0)] reg2524 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2523 = (1'h0);
  reg [(3'h4):(1'h0)] reg2522 = (1'h0);
  reg [(4'hf):(1'h0)] reg2521 = (1'h0);
  reg [(4'hd):(1'h0)] reg2517 = (1'h0);
  reg [(3'h6):(1'h0)] reg2516 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2515 = (1'h0);
  reg [(5'h10):(1'h0)] reg2514 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2512 = (1'h0);
  reg [(5'h10):(1'h0)] reg2511 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2510 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2509 = (1'h0);
  reg [(4'hf):(1'h0)] reg2508 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2507 = (1'h0);
  reg [(4'h8):(1'h0)] reg2506 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2505 = (1'h0);
  reg [(2'h3):(1'h0)] reg2504 = (1'h0);
  reg [(2'h2):(1'h0)] reg2503 = (1'h0);
  reg [(5'h10):(1'h0)] reg2502 = (1'h0);
  reg [(3'h4):(1'h0)] reg2501 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2500 = (1'h0);
  reg [(5'h10):(1'h0)] reg2499 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2498 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2496 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2495 = (1'h0);
  reg [(2'h2):(1'h0)] reg2494 = (1'h0);
  reg [(4'hf):(1'h0)] reg2493 = (1'h0);
  reg [(4'h9):(1'h0)] reg2491 = (1'h0);
  reg [(3'h5):(1'h0)] reg2487 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2486 = (1'h0);
  reg [(4'ha):(1'h0)] reg2485 = (1'h0);
  reg [(4'ha):(1'h0)] reg2483 = (1'h0);
  reg [(3'h7):(1'h0)] reg2482 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2481 = (1'h0);
  reg [(3'h4):(1'h0)] reg2480 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2479 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2478 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2477 = (1'h0);
  reg [(3'h4):(1'h0)] reg2476 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2475 = (1'h0);
  reg [(2'h2):(1'h0)] reg2473 = (1'h0);
  reg [(4'hd):(1'h0)] reg2471 = (1'h0);
  reg [(5'h10):(1'h0)] reg2470 = (1'h0);
  reg [(4'h9):(1'h0)] reg2469 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2468 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2465 = (1'h0);
  reg [(4'hd):(1'h0)] reg2467 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2466 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2464 = (1'h0);
  reg [(4'hf):(1'h0)] reg2463 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2462 = (1'h0);
  reg [(4'hd):(1'h0)] reg2460 = (1'h0);
  reg [(5'h10):(1'h0)] reg2459 = (1'h0);
  reg [(5'h10):(1'h0)] reg2458 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2457 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2453 = (1'h0);
  reg [(4'hf):(1'h0)] reg2451 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2450 = (1'h0);
  reg [(5'h10):(1'h0)] reg2449 = (1'h0);
  reg [(4'he):(1'h0)] reg2448 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2447 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2446 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2445 = (1'h0);
  reg [(3'h5):(1'h0)] reg2444 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2442 = (1'h0);
  reg [(4'he):(1'h0)] reg2440 = (1'h0);
  reg [(4'h8):(1'h0)] reg2439 = (1'h0);
  reg [(2'h2):(1'h0)] reg2438 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2437 = (1'h0);
  reg [(3'h7):(1'h0)] reg2433 = (1'h0);
  reg [(5'h10):(1'h0)] reg2418 = (1'h0);
  reg [(2'h3):(1'h0)] reg2404 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2399 = (1'h0);
  reg [(3'h4):(1'h0)] reg2398 = (1'h0);
  reg [(3'h7):(1'h0)] reg2386 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2385 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2364 = (1'h0);
  reg [(3'h7):(1'h0)] reg2361 = (1'h0);
  reg [(3'h6):(1'h0)] reg2356 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2355 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2341 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2340 = (1'h0);
  reg [(4'he):(1'h0)] reg2337 = (1'h0);
  reg [(4'he):(1'h0)] reg2432 = (1'h0);
  reg [(3'h7):(1'h0)] reg2431 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2429 = (1'h0);
  reg [(4'h9):(1'h0)] reg2428 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2427 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2425 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2424 = (1'h0);
  reg [(4'h9):(1'h0)] reg2423 = (1'h0);
  reg [(2'h2):(1'h0)] reg2422 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2421 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2420 = (1'h0);
  reg [(3'h6):(1'h0)] reg2417 = (1'h0);
  reg [(4'h8):(1'h0)] reg2416 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2415 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2414 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2413 = (1'h0);
  reg [(3'h5):(1'h0)] reg2407 = (1'h0);
  reg [(4'hd):(1'h0)] reg2412 = (1'h0);
  reg [(4'hd):(1'h0)] reg2411 = (1'h0);
  reg [(4'h8):(1'h0)] reg2410 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2409 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2408 = (1'h0);
  reg [(3'h4):(1'h0)] reg2406 = (1'h0);
  reg [(2'h3):(1'h0)] reg2405 = (1'h0);
  reg [(4'h8):(1'h0)] reg2403 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2402 = (1'h0);
  reg [(3'h7):(1'h0)] reg2401 = (1'h0);
  reg [(3'h7):(1'h0)] reg2400 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2397 = (1'h0);
  reg [(3'h5):(1'h0)] reg2396 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2395 = (1'h0);
  reg [(4'hf):(1'h0)] reg2393 = (1'h0);
  reg [(4'h9):(1'h0)] reg2392 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2391 = (1'h0);
  reg [(3'h4):(1'h0)] reg2390 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2389 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2388 = (1'h0);
  reg [(3'h5):(1'h0)] reg2387 = (1'h0);
  reg [(5'h10):(1'h0)] reg2384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2383 = (1'h0);
  reg [(2'h2):(1'h0)] reg2382 = (1'h0);
  reg [(4'ha):(1'h0)] reg2381 = (1'h0);
  reg [(4'h8):(1'h0)] reg2379 = (1'h0);
  reg [(3'h7):(1'h0)] reg2373 = (1'h0);
  reg [(4'ha):(1'h0)] reg2378 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2377 = (1'h0);
  reg [(5'h10):(1'h0)] reg2376 = (1'h0);
  reg [(4'hf):(1'h0)] reg2375 = (1'h0);
  reg [(3'h7):(1'h0)] reg2374 = (1'h0);
  reg [(3'h7):(1'h0)] reg2372 = (1'h0);
  reg [(3'h4):(1'h0)] reg2371 = (1'h0);
  reg [(4'hb):(1'h0)] reg2370 = (1'h0);
  reg [(4'hd):(1'h0)] reg2369 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2368 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2367 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2366 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2365 = (1'h0);
  reg [(3'h4):(1'h0)] reg2363 = (1'h0);
  reg [(4'hd):(1'h0)] reg2362 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2360 = (1'h0);
  reg [(4'hd):(1'h0)] reg2359 = (1'h0);
  reg [(2'h3):(1'h0)] reg2358 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2357 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2354 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2353 = (1'h0);
  reg [(3'h5):(1'h0)] reg2352 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2351 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2350 = (1'h0);
  reg [(3'h6):(1'h0)] reg2349 = (1'h0);
  reg [(5'h10):(1'h0)] reg2348 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2347 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2346 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2345 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2344 = (1'h0);
  reg [(4'hd):(1'h0)] reg2343 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2342 = (1'h0);
  reg [(3'h4):(1'h0)] reg2339 = (1'h0);
  reg [(3'h4):(1'h0)] reg2338 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2336 = (1'h0);
  reg [(3'h5):(1'h0)] reg2335 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2334 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2333 = (1'h0);
  reg [(5'h10):(1'h0)] reg2330 = (1'h0);
  reg [(2'h2):(1'h0)] reg2329 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2328 = (1'h0);
  reg [(4'h9):(1'h0)] reg2327 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2326 = (1'h0);
  reg [(4'h9):(1'h0)] reg2325 = (1'h0);
  reg [(4'hc):(1'h0)] reg2324 = (1'h0);
  reg [(3'h4):(1'h0)] reg2323 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2322 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2320 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2319 = (1'h0);
  reg [(2'h2):(1'h0)] reg2318 = (1'h0);
  reg [(4'h9):(1'h0)] reg2317 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2316 = (1'h0);
  reg [(4'hf):(1'h0)] reg2315 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2314 = (1'h0);
  reg [(5'h10):(1'h0)] reg2312 = (1'h0);
  reg [(3'h5):(1'h0)] reg2313 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2311 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2309 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2308 = (1'h0);
  reg [(4'hb):(1'h0)] reg2307 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2306 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2305 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2304 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2303 = (1'h0);
  reg [(4'ha):(1'h0)] reg2302 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2301 = (1'h0);
  reg [(3'h6):(1'h0)] reg2298 = (1'h0);
  reg [(3'h4):(1'h0)] reg2297 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2296 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2295 = (1'h0);
  reg [(3'h6):(1'h0)] reg2293 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2292 = (1'h0);
  reg [(4'hd):(1'h0)] reg2291 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2290 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2289 = (1'h0);
  reg [(4'h9):(1'h0)] reg2288 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2287 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2286 = (1'h0);
  reg [(4'hc):(1'h0)] reg2285 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2270 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2283 = (1'h0);
  reg [(3'h6):(1'h0)] reg2282 = (1'h0);
  reg [(3'h5):(1'h0)] reg2281 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2280 = (1'h0);
  reg [(3'h5):(1'h0)] reg2279 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2278 = (1'h0);
  reg [(4'hd):(1'h0)] reg2277 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2276 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2275 = (1'h0);
  reg [(5'h10):(1'h0)] reg2274 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2273 = (1'h0);
  reg [(3'h7):(1'h0)] reg2272 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2271 = (1'h0);
  reg [(3'h6):(1'h0)] reg2269 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2268 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2263 = (1'h0);
  reg [(3'h6):(1'h0)] reg2260 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2267 = (1'h0);
  reg [(4'hd):(1'h0)] reg2266 = (1'h0);
  reg [(5'h10):(1'h0)] reg2265 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2264 = (1'h0);
  reg [(4'hf):(1'h0)] reg2262 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2261 = (1'h0);
  reg [(4'he):(1'h0)] reg2259 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2258 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2257 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2256 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2255 = (1'h0);
  reg [(4'hb):(1'h0)] reg2254 = (1'h0);
  reg [(4'h9):(1'h0)] reg2245 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2249 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2248 = (1'h0);
  reg [(2'h3):(1'h0)] reg2247 = (1'h0);
  reg [(2'h3):(1'h0)] reg2246 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2244 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2242 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2241 = (1'h0);
  reg [(3'h6):(1'h0)] reg2240 = (1'h0);
  reg [(2'h2):(1'h0)] reg2238 = (1'h0);
  reg [(2'h3):(1'h0)] reg2235 = (1'h0);
  reg [(3'h6):(1'h0)] reg2234 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2233 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2232 = (1'h0);
  reg [(4'hd):(1'h0)] reg2231 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2230 = (1'h0);
  reg [(4'hc):(1'h0)] reg2228 = (1'h0);
  reg [(4'h8):(1'h0)] reg2227 = (1'h0);
  reg [(2'h3):(1'h0)] reg2226 = (1'h0);
  reg [(4'h9):(1'h0)] reg2225 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2223 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2209 = (1'h0);
  reg [(3'h5):(1'h0)] reg2222 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2221 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2220 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2219 = (1'h0);
  reg [(4'he):(1'h0)] reg2218 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2216 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2215 = (1'h0);
  reg [(4'hc):(1'h0)] reg2203 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2198 = (1'h0);
  reg [(4'h8):(1'h0)] reg2196 = (1'h0);
  reg [(3'h7):(1'h0)] reg2214 = (1'h0);
  reg [(2'h3):(1'h0)] reg2213 = (1'h0);
  reg [(5'h10):(1'h0)] reg2212 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2211 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2210 = (1'h0);
  reg [(4'ha):(1'h0)] reg2208 = (1'h0);
  reg [(5'h10):(1'h0)] reg2207 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2206 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2205 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2204 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2202 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2201 = (1'h0);
  reg [(4'hb):(1'h0)] reg2200 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2199 = (1'h0);
  reg [(4'hb):(1'h0)] reg2197 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2194 = (1'h0);
  reg [(2'h3):(1'h0)] reg2193 = (1'h0);
  reg [(5'h10):(1'h0)] reg2191 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2190 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2189 = (1'h0);
  reg [(4'ha):(1'h0)] reg2188 = (1'h0);
  reg [(4'h8):(1'h0)] reg2187 = (1'h0);
  reg [(3'h6):(1'h0)] reg2186 = (1'h0);
  reg [(2'h2):(1'h0)] reg2183 = (1'h0);
  reg [(2'h2):(1'h0)] reg2179 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2185 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2184 = (1'h0);
  reg [(3'h7):(1'h0)] reg2182 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2181 = (1'h0);
  reg [(4'he):(1'h0)] reg2180 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2178 = (1'h0);
  reg [(3'h4):(1'h0)] reg2177 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2176 = (1'h0);
  reg [(4'hf):(1'h0)] reg2175 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2172 = (1'h0);
  reg [(4'hd):(1'h0)] reg2170 = (1'h0);
  reg [(4'ha):(1'h0)] reg2169 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2168 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2165 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2164 = (1'h0);
  reg [(4'ha):(1'h0)] reg2163 = (1'h0);
  reg [(4'ha):(1'h0)] reg2162 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2160 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2159 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2154 = (1'h0);
  reg [(3'h5):(1'h0)] reg2158 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2157 = (1'h0);
  reg [(4'he):(1'h0)] reg2156 = (1'h0);
  reg [(4'hf):(1'h0)] reg2155 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2153 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2151 = (1'h0);
  reg [(3'h6):(1'h0)] reg2150 = (1'h0);
  reg [(2'h3):(1'h0)] reg2147 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2131 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2127 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2124 = (1'h0);
  reg [(3'h7):(1'h0)] reg2149 = (1'h0);
  reg [(2'h2):(1'h0)] reg2148 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2146 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2145 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2144 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2143 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2142 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2141 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2134 = (1'h0);
  reg [(4'hb):(1'h0)] reg2139 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2138 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2137 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2136 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2135 = (1'h0);
  reg [(4'hf):(1'h0)] reg2133 = (1'h0);
  reg [(5'h10):(1'h0)] reg2120 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2132 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2130 = (1'h0);
  reg [(2'h3):(1'h0)] reg2129 = (1'h0);
  reg [(4'h9):(1'h0)] reg2128 = (1'h0);
  reg [(2'h3):(1'h0)] reg2126 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2125 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2123 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2122 = (1'h0);
  reg [(3'h4):(1'h0)] reg2121 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2118 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2117 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2116 = (1'h0);
  reg [(3'h7):(1'h0)] reg2115 = (1'h0);
  reg [(4'ha):(1'h0)] reg2113 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2112 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2111 = (1'h0);
  reg [(4'h8):(1'h0)] reg2110 = (1'h0);
  reg [(4'h9):(1'h0)] reg2108 = (1'h0);
  reg [(3'h4):(1'h0)] reg2107 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2106 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2097 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2095 = (1'h0);
  reg [(4'he):(1'h0)] reg2087 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2086 = (1'h0);
  reg [(3'h7):(1'h0)] reg2105 = (1'h0);
  reg [(4'hd):(1'h0)] reg2104 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2103 = (1'h0);
  reg [(2'h3):(1'h0)] reg2102 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2100 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2099 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2098 = (1'h0);
  reg [(4'he):(1'h0)] reg2094 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2093 = (1'h0);
  reg [(5'h10):(1'h0)] reg2092 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2090 = (1'h0);
  reg [(4'hc):(1'h0)] reg2089 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2088 = (1'h0);
  reg [(4'hd):(1'h0)] reg2085 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2084 = (1'h0);
  reg [(5'h10):(1'h0)] reg2069 = (1'h0);
  reg [(2'h3):(1'h0)] reg2072 = (1'h0);
  reg [(4'ha):(1'h0)] reg2083 = (1'h0);
  reg [(3'h5):(1'h0)] reg2082 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2081 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2080 = (1'h0);
  reg [(2'h3):(1'h0)] reg2079 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2078 = (1'h0);
  reg [(3'h5):(1'h0)] reg2077 = (1'h0);
  reg [(4'he):(1'h0)] reg2076 = (1'h0);
  reg [(5'h10):(1'h0)] reg2075 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2074 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2073 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2071 = (1'h0);
  reg [(4'hb):(1'h0)] reg2070 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2068 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2067 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2056 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2062 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2055 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2054 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2049 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2036 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2035 = (1'h0);
  reg [(4'h8):(1'h0)] reg2066 = (1'h0);
  reg [(4'hf):(1'h0)] reg2065 = (1'h0);
  reg [(2'h3):(1'h0)] reg2064 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2063 = (1'h0);
  reg [(3'h5):(1'h0)] reg2061 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2060 = (1'h0);
  reg [(2'h2):(1'h0)] reg2059 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2058 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2057 = (1'h0);
  reg [(5'h10):(1'h0)] reg2053 = (1'h0);
  reg [(4'hc):(1'h0)] reg2052 = (1'h0);
  reg [(3'h6):(1'h0)] reg2051 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2050 = (1'h0);
  reg [(3'h7):(1'h0)] reg2048 = (1'h0);
  reg [(4'hd):(1'h0)] reg2047 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2046 = (1'h0);
  reg [(2'h3):(1'h0)] reg2045 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2043 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2042 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2041 = (1'h0);
  reg [(4'hd):(1'h0)] reg2040 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2039 = (1'h0);
  reg [(4'ha):(1'h0)] reg2038 = (1'h0);
  reg [(2'h3):(1'h0)] reg2037 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2033 = (1'h0);
  reg [(4'he):(1'h0)] reg1497 = (1'h0);
  reg [(4'he):(1'h0)] reg1494 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1483 = (1'h0);
  reg [(3'h5):(1'h0)] reg1533 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1539 = (1'h0);
  reg [(4'h9):(1'h0)] reg1538 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1537 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1536 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1535 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1534 = (1'h0);
  reg [(4'he):(1'h0)] reg1532 = (1'h0);
  reg [(4'hd):(1'h0)] reg1531 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1530 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1529 = (1'h0);
  reg [(5'h10):(1'h0)] reg1527 = (1'h0);
  reg [(3'h4):(1'h0)] reg1526 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1525 = (1'h0);
  reg [(3'h7):(1'h0)] reg1524 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1522 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1521 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1520 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1519 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1517 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1516 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1514 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1515 = (1'h0);
  reg [(4'h8):(1'h0)] reg1513 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1512 = (1'h0);
  reg [(3'h7):(1'h0)] reg1511 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1484 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1509 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1508 = (1'h0);
  reg [(4'ha):(1'h0)] reg1507 = (1'h0);
  reg [(4'ha):(1'h0)] reg1506 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1505 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1504 = (1'h0);
  reg [(2'h3):(1'h0)] reg1503 = (1'h0);
  reg [(4'he):(1'h0)] reg1502 = (1'h0);
  reg [(4'hf):(1'h0)] reg1501 = (1'h0);
  reg [(3'h5):(1'h0)] reg1500 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1499 = (1'h0);
  reg [(3'h5):(1'h0)] reg1498 = (1'h0);
  reg [(3'h6):(1'h0)] reg1496 = (1'h0);
  reg [(3'h4):(1'h0)] reg1495 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1493 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1492 = (1'h0);
  reg [(3'h5):(1'h0)] reg1491 = (1'h0);
  reg [(3'h7):(1'h0)] reg1490 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1489 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1488 = (1'h0);
  reg [(4'ha):(1'h0)] reg1487 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1486 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1485 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1482 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1481 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1480 = (1'h0);
  reg [(3'h5):(1'h0)] reg1479 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1478 = (1'h0);
  reg [(4'hd):(1'h0)] reg1477 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1476 = (1'h0);
  reg [(2'h3):(1'h0)] reg1475 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1473 = (1'h0);
  reg [(4'h8):(1'h0)] reg1472 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1471 = (1'h0);
  reg [(4'hc):(1'h0)] reg1469 = (1'h0);
  reg [(3'h4):(1'h0)] reg1468 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1467 = (1'h0);
  reg [(3'h4):(1'h0)] reg1465 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1464 = (1'h0);
  reg [(3'h5):(1'h0)] reg1463 = (1'h0);
  reg [(3'h4):(1'h0)] reg1462 = (1'h0);
  reg [(4'hd):(1'h0)] reg1461 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1460 = (1'h0);
  reg [(3'h6):(1'h0)] reg1459 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1458 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1457 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1456 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1455 = (1'h0);
  reg [(2'h3):(1'h0)] reg1454 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1453 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1452 = (1'h0);
  reg [(3'h4):(1'h0)] reg1449 = (1'h0);
  reg [(2'h3):(1'h0)] reg1447 = (1'h0);
  reg [(4'h8):(1'h0)] reg1451 = (1'h0);
  reg [(3'h4):(1'h0)] reg1450 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1448 = (1'h0);
  reg [(3'h6):(1'h0)] reg1440 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1446 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1445 = (1'h0);
  reg [(4'h9):(1'h0)] reg1444 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1443 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1442 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1441 = (1'h0);
  reg [(4'h9):(1'h0)] reg1438 = (1'h0);
  reg [(4'hf):(1'h0)] reg1437 = (1'h0);
  reg [(4'hf):(1'h0)] reg1436 = (1'h0);
  reg [(4'hc):(1'h0)] reg1435 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1423 = (1'h0);
  reg [(4'h8):(1'h0)] reg1434 = (1'h0);
  reg [(3'h5):(1'h0)] reg1433 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1432 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1431 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1430 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1429 = (1'h0);
  reg [(3'h4):(1'h0)] reg1428 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1427 = (1'h0);
  reg [(4'hc):(1'h0)] reg1426 = (1'h0);
  reg [(3'h6):(1'h0)] reg1425 = (1'h0);
  reg [(2'h3):(1'h0)] reg1424 = (1'h0);
  reg [(3'h6):(1'h0)] reg1422 = (1'h0);
  reg [(3'h5):(1'h0)] reg1421 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1420 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1419 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1418 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1417 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2576 = (1'h0);
  reg [(4'he):(1'h0)] forvar2571 = (1'h0);
  reg [(4'he):(1'h0)] forvar2565 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2584 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2580 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2579 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2577 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2567 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2564 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2559 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2556 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2550 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2545 = (1'h0);
  reg [(4'he):(1'h0)] forvar2543 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2542 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2540 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2535 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2530 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2525 = (1'h0);
  reg [(4'he):(1'h0)] forvar2520 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2519 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2518 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2506 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2502 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2513 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2497 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2492 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2490 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2489 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2488 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2484 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2477 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2474 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2472 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2464 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2465 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2461 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2456 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2455 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2454 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2452 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2443 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2441 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2436 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2435 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2434 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2414 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2410 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2409 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2403 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2401 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2391 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2390 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2350 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2384 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2378 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2368 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2360 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2362 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2358 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2339 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2336 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2430 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2426 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2419 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2418 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2407 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2404 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2399 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2398 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2394 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2386 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2385 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2380 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2375 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2371 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2373 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2364 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2361 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2356 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2355 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2349 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2346 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2341 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2340 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2337 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2333 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2332 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2321 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2311 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2312 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2310 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2300 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2299 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2294 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2284 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2280 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2274 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2261 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2265 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2256 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2257 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2259 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2277 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2275 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2271 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2270 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2266 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2264 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2263 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2260 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2246 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2245 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2243 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2239 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2237 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2236 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2229 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2224 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2217 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2214 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2204 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2201 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2199 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2197 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2209 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2203 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2198 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2196 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2195 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2189 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2181 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2178 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2192 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2184 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2183 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2179 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2174 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2173 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2171 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2167 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2166 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2161 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2156 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2154 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2152 = (1'h0);
  reg [(4'he):(1'h0)] forvar2143 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2141 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2137 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2118 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2147 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2140 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2134 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2121 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2131 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2127 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2124 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2120 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2119 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2114 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2109 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2105 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2103 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2093 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2090 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2085 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2082 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2077 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2101 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2097 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2096 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2095 = (1'h0);
  reg [(4'he):(1'h0)] forvar2091 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2087 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2086 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2081 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2078 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2075 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2070 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2076 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2072 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2069 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2064 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2051 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2061 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2052 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2048 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2040 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2039 = (1'h0);
  reg [(4'he):(1'h0)] forvar2033 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2062 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2056 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2055 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2054 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2049 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2044 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2036 = (1'h0);
  reg [(4'he):(1'h0)] forvar2035 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2034 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2032 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1502 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1501 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1498 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1495 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1486 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1482 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1536 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1534 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1533 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1528 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1523 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1518 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1515 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1514 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1510 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1497 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1490 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1494 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1484 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1483 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1474 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1470 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1466 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1456 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1450 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1445 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1448 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1449 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1447 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1440 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1439 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1432 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1427 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1430 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1429 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1424 = (1'h0);
  reg [(4'he):(1'h0)] forvar1418 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1423 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1417 = (1'h0);
  assign y = {wire2539,
                 wire2331,
                 wire2253,
                 wire2252,
                 wire2251,
                 wire2250,
                 wire2031,
                 wire2030,
                 wire2029,
                 wire1416,
                 wire2027,
                 reg2540,
                 reg2584,
                 reg2580,
                 reg2577,
                 reg2585,
                 reg2583,
                 reg2582,
                 reg2581,
                 reg2578,
                 reg2576,
                 reg2575,
                 reg2574,
                 reg2573,
                 reg2572,
                 reg2571,
                 reg2570,
                 reg2569,
                 reg2568,
                 reg2567,
                 reg2566,
                 reg2565,
                 reg2564,
                 reg2563,
                 reg2562,
                 reg2561,
                 reg2560,
                 reg2558,
                 reg2557,
                 reg2555,
                 reg2554,
                 reg2553,
                 reg2552,
                 reg2551,
                 reg2549,
                 reg2548,
                 reg2547,
                 reg2546,
                 reg2544,
                 reg2541,
                 reg2538,
                 reg2537,
                 reg2536,
                 reg2534,
                 reg2533,
                 reg2532,
                 reg2531,
                 reg2520,
                 reg2529,
                 reg2528,
                 reg2527,
                 reg2526,
                 reg2525,
                 reg2524,
                 reg2523,
                 reg2522,
                 reg2521,
                 reg2517,
                 reg2516,
                 reg2515,
                 reg2514,
                 reg2512,
                 reg2511,
                 reg2510,
                 reg2509,
                 reg2508,
                 reg2507,
                 reg2506,
                 reg2505,
                 reg2504,
                 reg2503,
                 reg2502,
                 reg2501,
                 reg2500,
                 reg2499,
                 reg2498,
                 reg2496,
                 reg2495,
                 reg2494,
                 reg2493,
                 reg2491,
                 reg2487,
                 reg2486,
                 reg2485,
                 reg2483,
                 reg2482,
                 reg2481,
                 reg2480,
                 reg2479,
                 reg2478,
                 reg2477,
                 reg2476,
                 reg2475,
                 reg2473,
                 reg2471,
                 reg2470,
                 reg2469,
                 reg2468,
                 reg2465,
                 reg2467,
                 reg2466,
                 reg2464,
                 reg2463,
                 reg2462,
                 reg2460,
                 reg2459,
                 reg2458,
                 reg2457,
                 reg2453,
                 reg2451,
                 reg2450,
                 reg2449,
                 reg2448,
                 reg2447,
                 reg2446,
                 reg2445,
                 reg2444,
                 reg2442,
                 reg2440,
                 reg2439,
                 reg2438,
                 reg2437,
                 reg2433,
                 reg2418,
                 reg2404,
                 reg2399,
                 reg2398,
                 reg2386,
                 reg2385,
                 reg2364,
                 reg2361,
                 reg2356,
                 reg2355,
                 reg2341,
                 reg2340,
                 reg2337,
                 reg2432,
                 reg2431,
                 reg2429,
                 reg2428,
                 reg2427,
                 reg2425,
                 reg2424,
                 reg2423,
                 reg2422,
                 reg2421,
                 reg2420,
                 reg2417,
                 reg2416,
                 reg2415,
                 reg2414,
                 reg2413,
                 reg2407,
                 reg2412,
                 reg2411,
                 reg2410,
                 reg2409,
                 reg2408,
                 reg2406,
                 reg2405,
                 reg2403,
                 reg2402,
                 reg2401,
                 reg2400,
                 reg2397,
                 reg2396,
                 reg2395,
                 reg2393,
                 reg2392,
                 reg2391,
                 reg2390,
                 reg2389,
                 reg2388,
                 reg2387,
                 reg2384,
                 reg2383,
                 reg2382,
                 reg2381,
                 reg2379,
                 reg2373,
                 reg2378,
                 reg2377,
                 reg2376,
                 reg2375,
                 reg2374,
                 reg2372,
                 reg2371,
                 reg2370,
                 reg2369,
                 reg2368,
                 reg2367,
                 reg2366,
                 reg2365,
                 reg2363,
                 reg2362,
                 reg2360,
                 reg2359,
                 reg2358,
                 reg2357,
                 reg2354,
                 reg2353,
                 reg2352,
                 reg2351,
                 reg2350,
                 reg2349,
                 reg2348,
                 reg2347,
                 reg2346,
                 reg2345,
                 reg2344,
                 reg2343,
                 reg2342,
                 reg2339,
                 reg2338,
                 reg2336,
                 reg2335,
                 reg2334,
                 reg2333,
                 reg2330,
                 reg2329,
                 reg2328,
                 reg2327,
                 reg2326,
                 reg2325,
                 reg2324,
                 reg2323,
                 reg2322,
                 reg2320,
                 reg2319,
                 reg2318,
                 reg2317,
                 reg2316,
                 reg2315,
                 reg2314,
                 reg2312,
                 reg2313,
                 reg2311,
                 reg2309,
                 reg2308,
                 reg2307,
                 reg2306,
                 reg2305,
                 reg2304,
                 reg2303,
                 reg2302,
                 reg2301,
                 reg2298,
                 reg2297,
                 reg2296,
                 reg2295,
                 reg2293,
                 reg2292,
                 reg2291,
                 reg2290,
                 reg2289,
                 reg2288,
                 reg2287,
                 reg2286,
                 reg2285,
                 reg2270,
                 reg2283,
                 reg2282,
                 reg2281,
                 reg2280,
                 reg2279,
                 reg2278,
                 reg2277,
                 reg2276,
                 reg2275,
                 reg2274,
                 reg2273,
                 reg2272,
                 reg2271,
                 reg2269,
                 reg2268,
                 reg2263,
                 reg2260,
                 reg2267,
                 reg2266,
                 reg2265,
                 reg2264,
                 reg2262,
                 reg2261,
                 reg2259,
                 reg2258,
                 reg2257,
                 reg2256,
                 reg2255,
                 reg2254,
                 reg2245,
                 reg2249,
                 reg2248,
                 reg2247,
                 reg2246,
                 reg2244,
                 reg2242,
                 reg2241,
                 reg2240,
                 reg2238,
                 reg2235,
                 reg2234,
                 reg2233,
                 reg2232,
                 reg2231,
                 reg2230,
                 reg2228,
                 reg2227,
                 reg2226,
                 reg2225,
                 reg2223,
                 reg2209,
                 reg2222,
                 reg2221,
                 reg2220,
                 reg2219,
                 reg2218,
                 reg2216,
                 reg2215,
                 reg2203,
                 reg2198,
                 reg2196,
                 reg2214,
                 reg2213,
                 reg2212,
                 reg2211,
                 reg2210,
                 reg2208,
                 reg2207,
                 reg2206,
                 reg2205,
                 reg2204,
                 reg2202,
                 reg2201,
                 reg2200,
                 reg2199,
                 reg2197,
                 reg2194,
                 reg2193,
                 reg2191,
                 reg2190,
                 reg2189,
                 reg2188,
                 reg2187,
                 reg2186,
                 reg2183,
                 reg2179,
                 reg2185,
                 reg2184,
                 reg2182,
                 reg2181,
                 reg2180,
                 reg2178,
                 reg2177,
                 reg2176,
                 reg2175,
                 reg2172,
                 reg2170,
                 reg2169,
                 reg2168,
                 reg2165,
                 reg2164,
                 reg2163,
                 reg2162,
                 reg2160,
                 reg2159,
                 reg2154,
                 reg2158,
                 reg2157,
                 reg2156,
                 reg2155,
                 reg2153,
                 reg2151,
                 reg2150,
                 reg2147,
                 reg2131,
                 reg2127,
                 reg2124,
                 reg2149,
                 reg2148,
                 reg2146,
                 reg2145,
                 reg2144,
                 reg2143,
                 reg2142,
                 reg2141,
                 reg2134,
                 reg2139,
                 reg2138,
                 reg2137,
                 reg2136,
                 reg2135,
                 reg2133,
                 reg2120,
                 reg2132,
                 reg2130,
                 reg2129,
                 reg2128,
                 reg2126,
                 reg2125,
                 reg2123,
                 reg2122,
                 reg2121,
                 reg2118,
                 reg2117,
                 reg2116,
                 reg2115,
                 reg2113,
                 reg2112,
                 reg2111,
                 reg2110,
                 reg2108,
                 reg2107,
                 reg2106,
                 reg2097,
                 reg2095,
                 reg2087,
                 reg2086,
                 reg2105,
                 reg2104,
                 reg2103,
                 reg2102,
                 reg2100,
                 reg2099,
                 reg2098,
                 reg2094,
                 reg2093,
                 reg2092,
                 reg2090,
                 reg2089,
                 reg2088,
                 reg2085,
                 reg2084,
                 reg2069,
                 reg2072,
                 reg2083,
                 reg2082,
                 reg2081,
                 reg2080,
                 reg2079,
                 reg2078,
                 reg2077,
                 reg2076,
                 reg2075,
                 reg2074,
                 reg2073,
                 reg2071,
                 reg2070,
                 reg2068,
                 reg2067,
                 reg2056,
                 reg2062,
                 reg2055,
                 reg2054,
                 reg2049,
                 reg2036,
                 reg2035,
                 reg2066,
                 reg2065,
                 reg2064,
                 reg2063,
                 reg2061,
                 reg2060,
                 reg2059,
                 reg2058,
                 reg2057,
                 reg2053,
                 reg2052,
                 reg2051,
                 reg2050,
                 reg2048,
                 reg2047,
                 reg2046,
                 reg2045,
                 reg2043,
                 reg2042,
                 reg2041,
                 reg2040,
                 reg2039,
                 reg2038,
                 reg2037,
                 reg2033,
                 reg1497,
                 reg1494,
                 reg1483,
                 reg1533,
                 reg1539,
                 reg1538,
                 reg1537,
                 reg1536,
                 reg1535,
                 reg1534,
                 reg1532,
                 reg1531,
                 reg1530,
                 reg1529,
                 reg1527,
                 reg1526,
                 reg1525,
                 reg1524,
                 reg1522,
                 reg1521,
                 reg1520,
                 reg1519,
                 reg1517,
                 reg1516,
                 reg1514,
                 reg1515,
                 reg1513,
                 reg1512,
                 reg1511,
                 reg1484,
                 reg1509,
                 reg1508,
                 reg1507,
                 reg1506,
                 reg1505,
                 reg1504,
                 reg1503,
                 reg1502,
                 reg1501,
                 reg1500,
                 reg1499,
                 reg1498,
                 reg1496,
                 reg1495,
                 reg1493,
                 reg1492,
                 reg1491,
                 reg1490,
                 reg1489,
                 reg1488,
                 reg1487,
                 reg1486,
                 reg1485,
                 reg1482,
                 reg1481,
                 reg1480,
                 reg1479,
                 reg1478,
                 reg1477,
                 reg1476,
                 reg1475,
                 reg1473,
                 reg1472,
                 reg1471,
                 reg1469,
                 reg1468,
                 reg1467,
                 reg1465,
                 reg1464,
                 reg1463,
                 reg1462,
                 reg1461,
                 reg1460,
                 reg1459,
                 reg1458,
                 reg1457,
                 reg1456,
                 reg1455,
                 reg1454,
                 reg1453,
                 reg1452,
                 reg1449,
                 reg1447,
                 reg1451,
                 reg1450,
                 reg1448,
                 reg1440,
                 reg1446,
                 reg1445,
                 reg1444,
                 reg1443,
                 reg1442,
                 reg1441,
                 reg1438,
                 reg1437,
                 reg1436,
                 reg1435,
                 reg1423,
                 reg1434,
                 reg1433,
                 reg1432,
                 reg1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1427,
                 reg1426,
                 reg1425,
                 reg1424,
                 reg1422,
                 reg1421,
                 reg1420,
                 reg1419,
                 reg1418,
                 reg1417,
                 forvar2576,
                 forvar2571,
                 forvar2565,
                 forvar2584,
                 forvar2580,
                 forvar2579,
                 forvar2577,
                 forvar2567,
                 forvar2564,
                 forvar2559,
                 forvar2556,
                 forvar2550,
                 forvar2545,
                 forvar2543,
                 forvar2542,
                 forvar2540,
                 forvar2535,
                 forvar2530,
                 forvar2525,
                 forvar2520,
                 forvar2519,
                 forvar2518,
                 forvar2506,
                 forvar2502,
                 forvar2513,
                 forvar2497,
                 forvar2492,
                 forvar2490,
                 forvar2489,
                 forvar2488,
                 forvar2484,
                 forvar2477,
                 forvar2474,
                 forvar2472,
                 forvar2464,
                 forvar2465,
                 forvar2461,
                 forvar2456,
                 forvar2455,
                 forvar2454,
                 forvar2452,
                 forvar2443,
                 forvar2441,
                 forvar2436,
                 forvar2435,
                 forvar2434,
                 forvar2414,
                 forvar2410,
                 forvar2409,
                 forvar2403,
                 forvar2401,
                 forvar2391,
                 forvar2390,
                 forvar2350,
                 forvar2384,
                 forvar2378,
                 forvar2368,
                 forvar2360,
                 forvar2362,
                 forvar2358,
                 forvar2339,
                 forvar2336,
                 forvar2430,
                 forvar2426,
                 forvar2419,
                 forvar2418,
                 forvar2407,
                 forvar2404,
                 forvar2399,
                 forvar2398,
                 forvar2394,
                 forvar2386,
                 forvar2385,
                 forvar2380,
                 forvar2375,
                 forvar2371,
                 forvar2373,
                 forvar2364,
                 forvar2361,
                 forvar2356,
                 forvar2355,
                 forvar2349,
                 forvar2346,
                 forvar2341,
                 forvar2340,
                 forvar2337,
                 forvar2333,
                 forvar2332,
                 forvar2321,
                 forvar2311,
                 forvar2312,
                 forvar2310,
                 forvar2300,
                 forvar2299,
                 forvar2294,
                 forvar2284,
                 forvar2280,
                 forvar2274,
                 forvar2261,
                 forvar2265,
                 forvar2256,
                 forvar2257,
                 forvar2259,
                 forvar2277,
                 forvar2275,
                 forvar2271,
                 forvar2270,
                 forvar2266,
                 forvar2264,
                 forvar2263,
                 forvar2260,
                 forvar2246,
                 forvar2245,
                 forvar2243,
                 forvar2239,
                 forvar2237,
                 forvar2236,
                 forvar2229,
                 forvar2224,
                 forvar2217,
                 forvar2214,
                 forvar2204,
                 forvar2201,
                 forvar2199,
                 forvar2197,
                 forvar2209,
                 forvar2203,
                 forvar2198,
                 forvar2196,
                 forvar2195,
                 forvar2189,
                 forvar2181,
                 forvar2178,
                 forvar2192,
                 forvar2184,
                 forvar2183,
                 forvar2179,
                 forvar2174,
                 forvar2173,
                 forvar2171,
                 forvar2167,
                 forvar2166,
                 forvar2161,
                 forvar2156,
                 forvar2154,
                 forvar2152,
                 forvar2143,
                 forvar2141,
                 forvar2137,
                 forvar2118,
                 forvar2147,
                 forvar2140,
                 forvar2134,
                 forvar2121,
                 forvar2131,
                 forvar2127,
                 forvar2124,
                 forvar2120,
                 forvar2119,
                 forvar2114,
                 forvar2109,
                 forvar2105,
                 forvar2103,
                 forvar2093,
                 forvar2090,
                 forvar2085,
                 forvar2082,
                 forvar2077,
                 forvar2101,
                 forvar2097,
                 forvar2096,
                 forvar2095,
                 forvar2091,
                 forvar2087,
                 forvar2086,
                 forvar2081,
                 forvar2078,
                 forvar2075,
                 forvar2070,
                 forvar2076,
                 forvar2072,
                 forvar2069,
                 forvar2064,
                 forvar2051,
                 forvar2061,
                 forvar2052,
                 forvar2048,
                 forvar2040,
                 forvar2039,
                 forvar2033,
                 forvar2062,
                 forvar2056,
                 forvar2055,
                 forvar2054,
                 forvar2049,
                 forvar2044,
                 forvar2036,
                 forvar2035,
                 forvar2034,
                 forvar2032,
                 forvar1502,
                 forvar1501,
                 forvar1498,
                 forvar1495,
                 forvar1486,
                 forvar1482,
                 forvar1536,
                 forvar1534,
                 forvar1533,
                 forvar1528,
                 forvar1523,
                 forvar1518,
                 forvar1515,
                 forvar1514,
                 forvar1510,
                 forvar1497,
                 forvar1490,
                 forvar1494,
                 forvar1484,
                 forvar1483,
                 forvar1474,
                 forvar1470,
                 forvar1466,
                 forvar1456,
                 forvar1450,
                 forvar1445,
                 forvar1448,
                 forvar1449,
                 forvar1447,
                 forvar1440,
                 forvar1439,
                 forvar1432,
                 forvar1427,
                 forvar1430,
                 forvar1429,
                 forvar1424,
                 forvar1418,
                 forvar1423,
                 forvar1417,
                 (1'h0)};
  assign wire1416 = $signed(((wire1413 & wire1414[(3'h6):(3'h6)]) <= $unsigned({wire1412})));
  always
    @(posedge clk) begin
      if (wire1414)
        begin
          if ($signed((^~(!$signed((8'hb8))))))
            begin
              reg1417 <= {(+(&$unsigned(wire1413)))};
              reg1418 <= $signed(wire1412[(3'h4):(1'h0)]);
            end
          else
            begin
              for (forvar1417 = (1'h0); (forvar1417 < (2'h2)); forvar1417 = (forvar1417 + (1'h1)))
                begin
                  if (wire1416)
                    begin
                      reg1418 <= ($signed(wire1414) ?
                          reg1418[(1'h1):(1'h0)] : reg1417[(1'h0):(1'h0)]);
                      reg1419 <= $unsigned(reg1417);
                      reg1420 <= wire1415[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1418 <= wire1413;
                    end
                  reg1421 <= (!wire1413);
                end
              reg1422 <= (|($signed(reg1418[(1'h0):(1'h0)]) * (wire1415 > (wire1414 ?
                  reg1419 : reg1417))));
              for (forvar1423 = (1'h0); (forvar1423 < (1'h1)); forvar1423 = (forvar1423 + (1'h1)))
                begin
                  if ($signed($signed($unsigned((8'hb2)))))
                    begin
                      reg1424 <= ($unsigned(reg1421[(3'h4):(2'h2)]) ?
                          $signed(((wire1413 ? wire1416 : (8'hb6)) ?
                              (reg1417 - reg1421) : $signed(reg1419))) : (forvar1423 | (^~(8'ha3))));
                      reg1425 <= wire1415;
                      reg1426 <= reg1421[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg1424 <= reg1425[(2'h3):(1'h1)];
                      reg1425 <= ((-forvar1423[(4'ha):(3'h5)]) ?
                          {{(-wire1415)}} : reg1417);
                      reg1426 <= $signed(wire1416[(4'ha):(4'h8)]);
                    end
                  if (({(~$unsigned(wire1414))} && wire1416))
                    begin
                      reg1427 <= {(|$signed((wire1413 << reg1419)))};
                      reg1428 <= $unsigned({$unsigned(reg1421)});
                    end
                  else
                    begin
                      reg1427 <= $signed(($signed(((8'hba) ?
                          (8'hb1) : reg1425)) <= reg1421[(3'h5):(2'h2)]));
                      reg1428 <= forvar1417[(1'h0):(1'h0)];
                      reg1429 <= forvar1417[(3'h5):(3'h4)];
                      reg1430 <= reg1424[(2'h3):(2'h2)];
                    end
                  if (reg1418[(2'h3):(2'h3)])
                    begin
                      reg1431 <= (^~($unsigned(reg1427[(1'h1):(1'h0)]) >>> $unsigned({reg1425})));
                      reg1432 <= reg1430;
                    end
                  else
                    begin
                      reg1431 <= reg1420;
                      reg1432 <= wire1415[(1'h1):(1'h0)];
                      reg1433 <= wire1413[(2'h2):(1'h0)];
                    end
                  reg1434 <= (reg1421 >>> reg1433);
                end
            end
        end
      else
        begin
          if (((~&(8'hb0)) <= reg1432))
            begin
              for (forvar1417 = (1'h0); (forvar1417 < (1'h0)); forvar1417 = (forvar1417 + (1'h1)))
                begin
                  for (forvar1418 = (1'h0); (forvar1418 < (2'h3)); forvar1418 = (forvar1418 + (1'h1)))
                    begin
                      reg1419 <= {reg1418[(1'h0):(1'h0)]};
                    end
                  if (forvar1418[(3'h5):(1'h1)])
                    begin
                      reg1420 <= (wire1415 ?
                          ($unsigned($signed(reg1421)) < reg1420[(4'h9):(1'h0)]) : wire1415);
                      reg1421 <= (^wire1412);
                    end
                  else
                    begin
                      reg1420 <= $signed(reg1430[(1'h1):(1'h1)]);
                      reg1421 <= $unsigned((|((reg1427 <= reg1431) <= reg1426)));
                      reg1422 <= $unsigned($signed(($signed(reg1420) ?
                          ((8'haa) ? wire1414 : reg1419) : reg1430)));
                      reg1423 <= forvar1423[(4'hb):(1'h1)];
                    end
                  for (forvar1424 = (1'h0); (forvar1424 < (1'h1)); forvar1424 = (forvar1424 + (1'h1)))
                    begin
                      reg1425 <= (reg1422[(3'h6):(3'h6)] ?
                          reg1421 : $signed(((8'ha1) ?
                              ((8'haf) ? wire1414 : reg1432) : (8'ha9))));
                      reg1426 <= (&reg1428);
                      reg1427 <= $unsigned((((reg1425 ?
                              reg1423 : reg1424) >= (-reg1427)) ?
                          ((wire1412 + reg1424) < (reg1431 ?
                              reg1428 : forvar1417)) : {{reg1421}}));
                      reg1428 <= (~^(8'hae));
                    end
                end
              for (forvar1429 = (1'h0); (forvar1429 < (2'h2)); forvar1429 = (forvar1429 + (1'h1)))
                begin
                  for (forvar1430 = (1'h0); (forvar1430 < (2'h2)); forvar1430 = (forvar1430 + (1'h1)))
                    begin
                      reg1431 <= (-$unsigned($unsigned((reg1431 ?
                          forvar1417 : reg1425))));
                      reg1432 <= ((forvar1430 ?
                          reg1419 : forvar1418[(2'h3):(2'h3)]) >= $unsigned($unsigned((~|forvar1423))));
                    end
                end
              if (((~(reg1427[(1'h1):(1'h1)] ?
                      (reg1427 ^ wire1416) : $unsigned(reg1417))) ?
                  $unsigned((~^(reg1419 || wire1416))) : $unsigned(($unsigned(reg1423) ?
                      $signed(forvar1417) : $unsigned(reg1426)))))
                begin
                  if ($signed($signed(((reg1430 ? reg1434 : reg1433) ?
                      (reg1422 ? reg1434 : forvar1430) : (+(8'hae))))))
                    begin
                      reg1433 <= {(($unsigned(reg1418) <= $unsigned(reg1428)) << $unsigned($unsigned(reg1429)))};
                      reg1434 <= forvar1429;
                      reg1435 <= reg1426;
                    end
                  else
                    begin
                      reg1433 <= reg1425;
                      reg1434 <= $signed($unsigned(((reg1430 ?
                          reg1418 : forvar1430) >= (reg1423 ?
                          reg1431 : wire1416))));
                    end
                end
              else
                begin
                  reg1433 <= $signed(wire1414[(2'h2):(2'h2)]);
                end
            end
          else
            begin
              if ($signed($unsigned($signed(reg1432))))
                begin
                  for (forvar1417 = (1'h0); (forvar1417 < (1'h1)); forvar1417 = (forvar1417 + (1'h1)))
                    begin
                      reg1418 <= (|reg1427[(1'h0):(1'h0)]);
                      reg1419 <= reg1426[(4'h9):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar1417 = (1'h0); (forvar1417 < (2'h3)); forvar1417 = (forvar1417 + (1'h1)))
                    begin
                      reg1418 <= reg1423[(2'h2):(1'h0)];
                      reg1419 <= ((~{(forvar1430 >> reg1428)}) ?
                          (8'ha7) : (~|$signed($signed((8'hb8)))));
                    end
                end
              if (((-{(reg1425 & reg1420)}) ?
                  ($unsigned($unsigned(reg1435)) ?
                      reg1435 : forvar1430) : $signed($signed($signed(forvar1424)))))
                begin
                  if ((((~&$unsigned(wire1416)) ?
                          {(&reg1432)} : ({reg1426} >= (reg1427 | reg1428))) ?
                      (({(8'haf)} - (~forvar1430)) ~^ {$unsigned(reg1428)}) : $unsigned($signed((~forvar1423)))))
                    begin
                      reg1420 <= (-reg1419[(1'h0):(1'h0)]);
                      reg1421 <= (+forvar1417);
                      reg1422 <= (wire1415[(2'h2):(1'h1)] && reg1427[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg1420 <= {forvar1430};
                    end
                  for (forvar1423 = (1'h0); (forvar1423 < (2'h2)); forvar1423 = (forvar1423 + (1'h1)))
                    begin
                      reg1424 <= (8'hb9);
                      reg1425 <= reg1428[(1'h1):(1'h0)];
                      reg1426 <= (~$signed((~|reg1433[(1'h1):(1'h0)])));
                    end
                  for (forvar1427 = (1'h0); (forvar1427 < (1'h1)); forvar1427 = (forvar1427 + (1'h1)))
                    begin
                      reg1428 <= $unsigned(wire1415[(1'h0):(1'h0)]);
                      reg1429 <= (!reg1426[(3'h4):(2'h2)]);
                      reg1430 <= (^$unsigned((~^$signed(reg1431))));
                      reg1431 <= $unsigned($unsigned(reg1429[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  if ($unsigned((!reg1426[(3'h6):(2'h3)])))
                    begin
                      reg1420 <= (($unsigned(((8'haf) ? reg1422 : wire1415)) ?
                          reg1421 : (reg1428 ?
                              {reg1435} : reg1421[(2'h2):(1'h1)])) >= $unsigned((8'ha8)));
                      reg1421 <= $unsigned((forvar1418[(4'ha):(2'h2)] <<< $signed($unsigned(reg1427))));
                      reg1422 <= ((^reg1423) ?
                          $signed(reg1426[(4'h9):(2'h3)]) : (((reg1425 ?
                                  forvar1427 : wire1416) <<< {wire1413}) ?
                              $signed((8'ha9)) : $signed(forvar1417)));
                      reg1423 <= $signed(reg1432[(3'h7):(1'h1)]);
                    end
                  else
                    begin
                      reg1420 <= reg1424[(1'h0):(1'h0)];
                    end
                end
              if ((8'hb0))
                begin
                  if ({$signed({(forvar1430 ? reg1422 : reg1419)})})
                    begin
                      reg1432 <= (^reg1435[(3'h6):(1'h1)]);
                      reg1433 <= ((+$signed((-reg1421))) ?
                          $unsigned(reg1423[(1'h0):(1'h0)]) : (forvar1430[(1'h1):(1'h1)] ?
                              reg1422[(3'h5):(3'h5)] : $signed(((8'h9d) ?
                                  reg1418 : reg1431))));
                    end
                  else
                    begin
                      reg1432 <= reg1435[(1'h0):(1'h0)];
                    end
                  if (forvar1424[(3'h4):(1'h0)])
                    begin
                      reg1434 <= ((-$signed((^reg1424))) >= $unsigned(reg1425[(3'h5):(1'h0)]));
                    end
                  else
                    begin
                      reg1434 <= {(~^(reg1424[(2'h3):(1'h1)] ?
                              $signed(wire1412) : (reg1435 ~^ reg1421)))};
                      reg1435 <= (~^({wire1415} ? {(&wire1414)} : {{reg1432}}));
                      reg1436 <= wire1413;
                    end
                  reg1437 <= (reg1418 == $signed((reg1419[(1'h1):(1'h0)] > (reg1432 >> reg1422))));
                end
              else
                begin
                  for (forvar1432 = (1'h0); (forvar1432 < (2'h2)); forvar1432 = (forvar1432 + (1'h1)))
                    begin
                      reg1433 <= forvar1417;
                      reg1434 <= ((($unsigned(reg1424) ^~ $unsigned(wire1412)) + $signed((reg1426 ?
                              (8'haa) : forvar1418))) ?
                          reg1432[(3'h6):(1'h1)] : $unsigned((^reg1436)));
                    end
                  if (reg1433)
                    begin
                      reg1435 <= ((reg1427[(1'h1):(1'h1)] ?
                          (^~reg1434[(1'h1):(1'h0)]) : $signed(forvar1423)) & ($unsigned((forvar1424 <<< reg1431)) == (reg1419 ?
                          (^~(8'ha2)) : (8'h9c))));
                      reg1436 <= reg1420[(3'h4):(2'h2)];
                      reg1437 <= reg1427[(1'h0):(1'h0)];
                      reg1438 <= {($signed((8'ha0)) * reg1426)};
                    end
                  else
                    begin
                      reg1435 <= $signed((^~((^~reg1421) >>> $signed(reg1419))));
                    end
                end
            end
        end
      for (forvar1439 = (1'h0); (forvar1439 < (2'h2)); forvar1439 = (forvar1439 + (1'h1)))
        begin
          if (($signed({reg1435}) && wire1416[(2'h2):(1'h0)]))
            begin
              if (reg1427[(1'h0):(1'h0)])
                begin
                  for (forvar1440 = (1'h0); (forvar1440 < (1'h1)); forvar1440 = (forvar1440 + (1'h1)))
                    begin
                      reg1441 <= wire1412[(3'h4):(2'h3)];
                      reg1442 <= (~(8'hb1));
                      reg1443 <= $signed($signed({$unsigned(reg1432)}));
                      reg1444 <= (8'hba);
                    end
                  reg1445 <= $signed((($signed(wire1415) <<< $signed(reg1421)) ?
                      ($signed(reg1432) ?
                          (|forvar1440) : (reg1417 > reg1442)) : ((!reg1437) ?
                          (+reg1432) : $signed(reg1423))));
                  reg1446 <= ($unsigned((8'hb8)) ?
                      ((^reg1433) + reg1437) : $unsigned($unsigned((-forvar1430))));
                end
              else
                begin
                  if ($unsigned(({(reg1441 >= (8'ha8))} ?
                      (&(reg1421 == reg1433)) : ($unsigned(forvar1432) ?
                          (reg1442 ? reg1446 : reg1445) : $unsigned(reg1418)))))
                    begin
                      reg1440 <= reg1427[(1'h1):(1'h0)];
                      reg1441 <= forvar1424[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg1440 <= (reg1429[(1'h0):(1'h0)] || reg1444[(1'h0):(1'h0)]);
                      reg1441 <= $signed((&(8'had)));
                    end
                end
              if (($signed($unsigned((forvar1430 ? reg1425 : (8'ha6)))) ?
                  $unsigned($signed((~|reg1429))) : $signed((-reg1443[(3'h5):(2'h3)]))))
                begin
                  for (forvar1447 = (1'h0); (forvar1447 < (1'h1)); forvar1447 = (forvar1447 + (1'h1)))
                    begin
                      reg1448 <= $unsigned($unsigned({reg1424[(1'h0):(1'h0)]}));
                    end
                  for (forvar1449 = (1'h0); (forvar1449 < (1'h1)); forvar1449 = (forvar1449 + (1'h1)))
                    begin
                      reg1450 <= reg1420;
                      reg1451 <= (reg1432 ?
                          reg1441[(2'h3):(2'h2)] : $unsigned(forvar1439));
                    end
                end
              else
                begin
                  if ((forvar1417[(4'hb):(3'h6)] * (-$unsigned((8'hb3)))))
                    begin
                      reg1447 <= ((forvar1429 ~^ reg1429[(3'h6):(1'h0)]) ?
                          ((~|((8'ha6) > reg1421)) ^~ reg1450[(2'h2):(1'h1)]) : $signed(((8'had) + (reg1441 ?
                              reg1422 : reg1436))));
                    end
                  else
                    begin
                      reg1447 <= $signed($unsigned(($signed(wire1412) < (reg1431 * (8'ha1)))));
                    end
                  for (forvar1448 = (1'h0); (forvar1448 < (2'h3)); forvar1448 = (forvar1448 + (1'h1)))
                    begin
                      reg1449 <= ({(!(reg1428 + reg1426))} & $unsigned($signed((8'hb5))));
                      reg1450 <= (~|(({(8'hae)} == (forvar1423 + reg1450)) * reg1427[(1'h1):(1'h0)]));
                      reg1451 <= forvar1427;
                    end
                  if ({(~(reg1438[(3'h5):(3'h5)] ?
                          $unsigned(reg1445) : $signed(wire1416)))})
                    begin
                      reg1452 <= (+reg1429[(1'h0):(1'h0)]);
                      reg1453 <= reg1440;
                    end
                  else
                    begin
                      reg1452 <= ($unsigned(reg1437[(1'h1):(1'h0)]) - ($unsigned((-forvar1449)) + ((reg1418 ?
                          reg1450 : (8'ha8)) ^~ $unsigned(reg1450))));
                    end
                  if ($signed((reg1437[(1'h1):(1'h1)] ?
                      reg1437[(4'h8):(3'h7)] : reg1440[(1'h1):(1'h1)])))
                    begin
                      reg1454 <= reg1432;
                    end
                  else
                    begin
                      reg1454 <= ((($unsigned(forvar1439) ?
                          {reg1435} : (~reg1428)) >= ((reg1426 != reg1420) >> $signed(reg1426))) * $unsigned(forvar1424));
                      reg1455 <= ((+(reg1442[(3'h7):(3'h4)] + reg1421)) >= (-$unsigned(reg1434)));
                      reg1456 <= reg1451;
                      reg1457 <= ({reg1456[(3'h6):(3'h6)]} ?
                          $unsigned(reg1437) : (~reg1454[(1'h1):(1'h0)]));
                    end
                end
            end
          else
            begin
              for (forvar1440 = (1'h0); (forvar1440 < (1'h1)); forvar1440 = (forvar1440 + (1'h1)))
                begin
                  if ($unsigned(reg1442))
                    begin
                      reg1441 <= reg1444[(4'h8):(2'h3)];
                      reg1442 <= ((~^wire1416) - ((~^(reg1454 >= reg1444)) ?
                          ((reg1435 | reg1422) ?
                              $unsigned(forvar1424) : (reg1438 <= reg1423)) : reg1427[(1'h1):(1'h0)]));
                      reg1443 <= $unsigned($signed(reg1428));
                      reg1444 <= ($unsigned($signed(wire1414[(3'h7):(3'h7)])) & (forvar1429[(4'hf):(4'he)] ?
                          reg1457[(4'ha):(3'h5)] : forvar1423));
                    end
                  else
                    begin
                      reg1441 <= (reg1450[(1'h0):(1'h0)] >>> wire1413[(1'h1):(1'h0)]);
                      reg1442 <= forvar1449;
                    end
                  for (forvar1445 = (1'h0); (forvar1445 < (2'h3)); forvar1445 = (forvar1445 + (1'h1)))
                    begin
                      reg1446 <= forvar1429;
                      reg1447 <= reg1455[(3'h5):(1'h0)];
                      reg1448 <= {(reg1424 <= ((reg1433 ?
                              wire1415 : (8'ha9)) <<< reg1450[(2'h3):(2'h3)]))};
                      reg1449 <= ($signed(reg1452[(2'h2):(2'h2)]) <<< ({(forvar1424 + wire1414)} != (^reg1447)));
                    end
                  for (forvar1450 = (1'h0); (forvar1450 < (1'h1)); forvar1450 = (forvar1450 + (1'h1)))
                    begin
                      reg1451 <= (~(((forvar1424 && reg1447) ^~ forvar1439[(1'h1):(1'h0)]) <<< $unsigned((8'hb9))));
                      reg1452 <= ($signed($unsigned({reg1425})) ?
                          (((reg1447 ? (8'ha3) : reg1456) ?
                                  (~forvar1440) : (8'ha9)) ?
                              reg1456 : ((forvar1417 ? forvar1450 : reg1454) ?
                                  (reg1435 - reg1421) : (forvar1424 <= forvar1423))) : forvar1430);
                      reg1453 <= (!reg1427);
                    end
                end
              if ((+$signed($signed((forvar1429 ? reg1444 : reg1452)))))
                begin
                  reg1454 <= ({$unsigned($unsigned(reg1454))} || wire1414);
                  reg1455 <= ((reg1447 ?
                      (+(|forvar1449)) : (^forvar1429[(2'h3):(1'h1)])) ^~ (8'hb8));
                  for (forvar1456 = (1'h0); (forvar1456 < (2'h3)); forvar1456 = (forvar1456 + (1'h1)))
                    begin
                      reg1457 <= $unsigned(reg1451);
                      reg1458 <= forvar1439[(2'h2):(2'h2)];
                      reg1459 <= forvar1429[(1'h0):(1'h0)];
                      reg1460 <= $signed(reg1421[(3'h5):(1'h0)]);
                    end
                end
              else
                begin
                  if ((-(^(&$signed(reg1459)))))
                    begin
                      reg1454 <= (^(8'h9c));
                    end
                  else
                    begin
                      reg1454 <= (forvar1417[(3'h6):(3'h5)] ?
                          {reg1427} : ($unsigned($unsigned(reg1443)) + reg1433[(3'h5):(1'h1)]));
                      reg1455 <= ((reg1437[(3'h5):(1'h0)] && reg1442) && (reg1444 && ((forvar1430 ^~ forvar1449) - $signed(reg1443))));
                    end
                  if ((8'hba))
                    begin
                      reg1456 <= (^~reg1430);
                      reg1457 <= $signed($signed((~forvar1439[(1'h1):(1'h0)])));
                      reg1458 <= $signed(reg1425[(1'h0):(1'h0)]);
                      reg1459 <= reg1441;
                    end
                  else
                    begin
                      reg1456 <= $signed(forvar1456[(4'h8):(1'h1)]);
                      reg1457 <= $unsigned((forvar1429[(3'h4):(2'h3)] >> reg1448[(2'h3):(1'h1)]));
                      reg1458 <= (8'ha2);
                    end
                end
              if ($unsigned((8'ha3)))
                begin
                  if ((|(+(&wire1416[(2'h3):(2'h2)]))))
                    begin
                      reg1461 <= (($unsigned((reg1434 < reg1426)) <<< ((wire1416 ?
                              reg1424 : forvar1427) ?
                          reg1420 : {reg1450})) <<< ($signed((forvar1445 ?
                          forvar1424 : reg1454)) & ($signed(forvar1430) ?
                          reg1448[(3'h7):(2'h2)] : $unsigned((8'haf)))));
                    end
                  else
                    begin
                      reg1461 <= $unsigned($signed(((~&(8'hae)) != reg1438[(3'h7):(2'h2)])));
                      reg1462 <= reg1454;
                    end
                  if ((($signed((reg1455 ^~ (8'ha0))) ?
                          (&$unsigned(reg1454)) : ((8'hb4) ?
                              $signed(reg1433) : {reg1451})) ?
                      $signed($signed({reg1425})) : reg1417[(1'h0):(1'h0)]))
                    begin
                      reg1463 <= (reg1429 ? wire1416[(3'h6):(3'h4)] : reg1459);
                    end
                  else
                    begin
                      reg1463 <= (!reg1446[(4'h9):(3'h5)]);
                      reg1464 <= $signed($unsigned((8'hb6)));
                      reg1465 <= $signed((reg1460[(1'h1):(1'h0)] ?
                          (+reg1454[(1'h1):(1'h0)]) : $signed((~&forvar1424))));
                    end
                  for (forvar1466 = (1'h0); (forvar1466 < (1'h1)); forvar1466 = (forvar1466 + (1'h1)))
                    begin
                      reg1467 <= (^~(reg1431 ^~ forvar1466));
                      reg1468 <= {(&reg1432)};
                      reg1469 <= reg1422[(2'h3):(1'h1)];
                    end
                  for (forvar1470 = (1'h0); (forvar1470 < (2'h3)); forvar1470 = (forvar1470 + (1'h1)))
                    begin
                      reg1471 <= ($signed(($signed(reg1426) ?
                          (reg1420 ?
                              (8'hae) : reg1449) : forvar1418)) + ((&$signed(reg1458)) ?
                          reg1469 : $unsigned({reg1449})));
                      reg1472 <= ($unsigned($signed((8'ha2))) ?
                          (+$signed({(8'hb0)})) : (({reg1469} ~^ $unsigned(reg1471)) | (8'ha3)));
                      reg1473 <= $signed(reg1442);
                    end
                end
              else
                begin
                  reg1461 <= (reg1459 ?
                      ((|(+(8'hb2))) ?
                          (8'ha2) : $unsigned((forvar1456 != reg1426))) : reg1428[(1'h0):(1'h0)]);
                end
              for (forvar1474 = (1'h0); (forvar1474 < (2'h2)); forvar1474 = (forvar1474 + (1'h1)))
                begin
                  if ((reg1433[(3'h4):(2'h2)] ?
                      reg1430 : $signed(reg1441[(1'h1):(1'h1)])))
                    begin
                      reg1475 <= (~&reg1473[(3'h5):(3'h4)]);
                    end
                  else
                    begin
                      reg1475 <= forvar1424[(2'h3):(2'h3)];
                      reg1476 <= $unsigned((reg1458 & (+$signed((8'hb6)))));
                    end
                  if ({(^({reg1437} ? reg1471[(4'hb):(3'h6)] : reg1447))})
                    begin
                      reg1477 <= reg1476;
                      reg1478 <= $signed({$unsigned({reg1457})});
                      reg1479 <= {{($signed(reg1443) >= reg1448)}};
                    end
                  else
                    begin
                      reg1477 <= $unsigned((($unsigned((8'hb6)) & (~reg1460)) ?
                          ($signed(reg1452) ?
                              (reg1429 ?
                                  reg1420 : reg1472) : (reg1426 > reg1447)) : ($unsigned(reg1437) - (|reg1420))));
                    end
                end
            end
          reg1480 <= $signed(forvar1447);
          reg1481 <= ($unsigned(reg1459[(1'h1):(1'h0)]) ?
              ({$signed(forvar1474)} * (reg1457 >>> reg1479)) : (reg1460 ?
                  ({forvar1445} ? (~forvar1450) : reg1428) : (forvar1445 ?
                      $unsigned(reg1441) : {forvar1429})));
        end
      if ({({(reg1451 ? (8'hb5) : reg1476)} ?
              reg1457[(3'h6):(2'h2)] : $unsigned(reg1460[(2'h3):(1'h0)]))})
        begin
          reg1482 <= $signed((8'ha7));
          if ((^reg1443))
            begin
              for (forvar1483 = (1'h0); (forvar1483 < (2'h2)); forvar1483 = (forvar1483 + (1'h1)))
                begin
                  for (forvar1484 = (1'h0); (forvar1484 < (2'h3)); forvar1484 = (forvar1484 + (1'h1)))
                    begin
                      reg1485 <= {$signed((~|wire1414[(3'h6):(1'h0)]))};
                    end
                  if (reg1455)
                    begin
                      reg1486 <= $unsigned((|(8'hb9)));
                    end
                  else
                    begin
                      reg1486 <= ((($unsigned(reg1444) && $signed(reg1423)) - {$unsigned(reg1427)}) ^~ reg1426);
                      reg1487 <= $unsigned($signed(($signed((8'hb2)) <<< reg1453[(3'h7):(2'h3)])));
                      reg1488 <= reg1427[(2'h3):(2'h3)];
                    end
                end
              if ((~^($unsigned($signed(reg1485)) ?
                  (reg1456[(4'h9):(1'h0)] + forvar1423[(1'h0):(1'h0)]) : $signed({wire1414}))))
                begin
                  reg1489 <= forvar1430;
                  if ((reg1430 ?
                      reg1461[(4'h9):(1'h0)] : forvar1466[(3'h4):(1'h1)]))
                    begin
                      reg1490 <= reg1428;
                    end
                  else
                    begin
                      reg1490 <= forvar1417;
                      reg1491 <= $signed($signed($signed(forvar1474[(1'h0):(1'h0)])));
                      reg1492 <= forvar1440[(1'h0):(1'h0)];
                      reg1493 <= (reg1490 <= $signed((reg1428[(2'h3):(2'h3)] ?
                          (|wire1415) : $unsigned(reg1453))));
                    end
                  for (forvar1494 = (1'h0); (forvar1494 < (1'h0)); forvar1494 = (forvar1494 + (1'h1)))
                    begin
                      reg1495 <= $unsigned((8'ha9));
                      reg1496 <= (-{(~(~|reg1435))});
                    end
                end
              else
                begin
                  if ($signed((~|$signed(((8'hb9) ? reg1475 : wire1415)))))
                    begin
                      reg1489 <= $unsigned(reg1419);
                    end
                  else
                    begin
                      reg1489 <= $signed((~&(~&reg1491)));
                    end
                  for (forvar1490 = (1'h0); (forvar1490 < (2'h3)); forvar1490 = (forvar1490 + (1'h1)))
                    begin
                      reg1491 <= $unsigned($signed(reg1429));
                      reg1492 <= ($signed((|((8'ha7) + reg1492))) ?
                          $unsigned(($signed(reg1424) ?
                              (~^reg1434) : $unsigned(reg1427))) : ($unsigned(forvar1427) >> $signed((reg1435 >= reg1479))));
                      reg1493 <= reg1454[(2'h2):(2'h2)];
                    end
                  for (forvar1494 = (1'h0); (forvar1494 < (1'h0)); forvar1494 = (forvar1494 + (1'h1)))
                    begin
                      reg1495 <= {(~|forvar1470[(4'h8):(3'h5)])};
                      reg1496 <= ($unsigned((!forvar1449)) ?
                          ($signed((forvar1430 ?
                              reg1493 : forvar1424)) >>> reg1475) : reg1492[(1'h0):(1'h0)]);
                    end
                end
              if ((reg1459 >> $unsigned(reg1471[(1'h1):(1'h1)])))
                begin
                  for (forvar1497 = (1'h0); (forvar1497 < (2'h3)); forvar1497 = (forvar1497 + (1'h1)))
                    begin
                      reg1498 <= (~&reg1457[(4'h9):(4'h9)]);
                    end
                end
              else
                begin
                  for (forvar1497 = (1'h0); (forvar1497 < (2'h3)); forvar1497 = (forvar1497 + (1'h1)))
                    begin
                      reg1498 <= $unsigned(reg1462[(2'h2):(1'h1)]);
                      reg1499 <= $signed(forvar1418);
                      reg1500 <= reg1467[(1'h1):(1'h1)];
                    end
                  if ($signed($signed({$unsigned(forvar1432)})))
                    begin
                      reg1501 <= $unsigned($unsigned(forvar1440[(3'h6):(2'h2)]));
                      reg1502 <= $unsigned((($unsigned(wire1416) >>> (~|forvar1445)) >> {(forvar1466 >= reg1487)}));
                    end
                  else
                    begin
                      reg1501 <= (((~&((8'ha7) ?
                          forvar1494 : (8'hb0))) + $signed(reg1487)) << ((~|(~&(8'ha6))) ?
                          reg1476 : wire1413[(1'h0):(1'h0)]));
                      reg1502 <= $signed($signed(((8'hba) ?
                          reg1501[(4'h9):(2'h2)] : $unsigned(forvar1448))));
                      reg1503 <= forvar1449;
                      reg1504 <= {(8'h9f)};
                    end
                  if (forvar1440)
                    begin
                      reg1505 <= $unsigned(({reg1422[(2'h2):(2'h2)]} ?
                          ((-reg1504) ?
                              (forvar1490 ?
                                  reg1487 : reg1418) : (~reg1501)) : {$signed(forvar1424)}));
                      reg1506 <= (~&(8'hae));
                      reg1507 <= ((~|reg1427) ~^ $unsigned({forvar1418}));
                      reg1508 <= ({reg1456} ?
                          (8'ha0) : {$unsigned({forvar1456})});
                    end
                  else
                    begin
                      reg1505 <= reg1421;
                    end
                end
              reg1509 <= ({((reg1481 == reg1420) ?
                          reg1420 : $signed(reg1487))} ?
                  reg1502 : $signed({reg1508}));
            end
          else
            begin
              for (forvar1483 = (1'h0); (forvar1483 < (1'h1)); forvar1483 = (forvar1483 + (1'h1)))
                begin
                  reg1484 <= $unsigned({reg1509});
                end
            end
          if ((^~$unsigned(forvar1427)))
            begin
              for (forvar1510 = (1'h0); (forvar1510 < (1'h0)); forvar1510 = (forvar1510 + (1'h1)))
                begin
                  if ((reg1468[(2'h3):(2'h3)] ?
                      reg1499 : reg1444[(4'h9):(3'h7)]))
                    begin
                      reg1511 <= ((($unsigned(reg1444) ?
                          forvar1423 : (~^(8'ha5))) ^~ ((~forvar1497) ?
                          (8'ha6) : {(8'hb3)})) >>> (($unsigned(forvar1497) ^ $signed(reg1446)) - reg1432));
                      reg1512 <= ((&reg1489) ?
                          {reg1436} : $unsigned($signed({reg1501})));
                      reg1513 <= $unsigned((($signed(reg1451) * (^~reg1476)) * reg1482[(4'hb):(4'h8)]));
                    end
                  else
                    begin
                      reg1511 <= $signed($signed(((-reg1433) >= reg1493)));
                      reg1512 <= (reg1438 ?
                          {((reg1425 ? wire1412 : reg1493) ?
                                  {forvar1466} : {reg1441})} : reg1433);
                      reg1513 <= reg1453;
                    end
                end
              for (forvar1514 = (1'h0); (forvar1514 < (2'h3)); forvar1514 = (forvar1514 + (1'h1)))
                begin
                  reg1515 <= (|((reg1505[(2'h2):(2'h2)] - $signed(reg1461)) ?
                      (8'h9c) : ((reg1422 ^~ reg1445) ?
                          $unsigned(reg1424) : $signed(reg1431))));
                end
            end
          else
            begin
              for (forvar1510 = (1'h0); (forvar1510 < (1'h1)); forvar1510 = (forvar1510 + (1'h1)))
                begin
                  if ({{reg1512[(1'h0):(1'h0)]}})
                    begin
                      reg1511 <= (~forvar1490[(1'h0):(1'h0)]);
                      reg1512 <= {$signed(forvar1494)};
                    end
                  else
                    begin
                      reg1511 <= $unsigned({$unsigned($signed(forvar1440))});
                      reg1512 <= {$unsigned((+{(8'ha2)}))};
                      reg1513 <= (^reg1503[(1'h0):(1'h0)]);
                      reg1514 <= (|(8'hb2));
                    end
                end
              for (forvar1515 = (1'h0); (forvar1515 < (1'h1)); forvar1515 = (forvar1515 + (1'h1)))
                begin
                  if ($unsigned((~&$signed(reg1476[(1'h1):(1'h0)]))))
                    begin
                      reg1516 <= ({reg1432} >> {((~^reg1493) >= (!reg1435))});
                      reg1517 <= (~&$signed((!reg1500)));
                    end
                  else
                    begin
                      reg1516 <= $signed(((~|$unsigned(forvar1456)) < {(8'ha3)}));
                      reg1517 <= reg1464[(2'h2):(2'h2)];
                    end
                  for (forvar1518 = (1'h0); (forvar1518 < (1'h1)); forvar1518 = (forvar1518 + (1'h1)))
                    begin
                      reg1519 <= reg1423[(1'h0):(1'h0)];
                      reg1520 <= ({reg1461} ^ {reg1450[(1'h1):(1'h1)]});
                      reg1521 <= (reg1509 >> reg1487[(3'h7):(3'h4)]);
                      reg1522 <= {({forvar1447[(3'h5):(1'h0)]} ?
                              $unsigned((&reg1502)) : $unsigned((reg1514 << wire1413)))};
                    end
                  for (forvar1523 = (1'h0); (forvar1523 < (2'h2)); forvar1523 = (forvar1523 + (1'h1)))
                    begin
                      reg1524 <= $signed({(~|$signed(reg1501))});
                      reg1525 <= $unsigned((|$unsigned(forvar1418)));
                      reg1526 <= (($signed((reg1524 <<< reg1506)) << ({reg1457} * (forvar1523 ?
                              wire1415 : (8'hb4)))) ?
                          (~|forvar1430) : (~&(~&(forvar1447 ?
                              reg1471 : (8'ha3)))));
                      reg1527 <= $signed($signed($unsigned(forvar1418)));
                    end
                  for (forvar1528 = (1'h0); (forvar1528 < (1'h0)); forvar1528 = (forvar1528 + (1'h1)))
                    begin
                      reg1529 <= ($signed(reg1477[(1'h1):(1'h0)]) ?
                          $unsigned($signed(reg1517)) : ($signed((reg1515 ?
                                  forvar1447 : reg1520)) ?
                              wire1413[(2'h2):(1'h0)] : $signed(((8'ha3) ?
                                  reg1462 : (8'ha5)))));
                      reg1530 <= ($unsigned(({reg1442} - reg1520)) ?
                          ((((8'haf) ? (8'hae) : reg1498) ?
                                  (reg1529 ? reg1422 : reg1529) : (^wire1413)) ?
                              $unsigned(reg1438) : $unsigned((~|reg1456))) : reg1512[(3'h5):(1'h1)]);
                      reg1531 <= reg1450;
                      reg1532 <= ((+$unsigned($unsigned(reg1513))) && $unsigned(reg1452));
                    end
                end
              if (({reg1432[(3'h7):(1'h0)]} ?
                  (8'hb7) : ((^~reg1464) ?
                      $signed($signed(reg1512)) : reg1425[(1'h1):(1'h1)])))
                begin
                  for (forvar1533 = (1'h0); (forvar1533 < (2'h2)); forvar1533 = (forvar1533 + (1'h1)))
                    begin
                      reg1534 <= $signed(($signed((reg1527 - reg1488)) <= (+(reg1449 < reg1455))));
                    end
                  reg1535 <= reg1449[(2'h2):(1'h1)];
                  if ($unsigned(((~$signed(reg1522)) >>> {reg1516})))
                    begin
                      reg1536 <= ($signed(reg1434) <<< (8'h9c));
                      reg1537 <= reg1492;
                      reg1538 <= {$signed(reg1487)};
                      reg1539 <= {$unsigned($signed((reg1487 ?
                              forvar1439 : reg1461)))};
                    end
                  else
                    begin
                      reg1536 <= ($signed(({reg1454} ^ (+reg1437))) * (8'hb3));
                      reg1537 <= reg1520[(1'h1):(1'h1)];
                      reg1538 <= $unsigned(reg1467[(3'h4):(2'h2)]);
                      reg1539 <= ($unsigned($signed($signed(reg1499))) <<< reg1507[(2'h3):(2'h2)]);
                    end
                end
              else
                begin
                  reg1533 <= ($signed((^~$signed(forvar1418))) ?
                      (~$unsigned($signed((8'ha4)))) : reg1519[(2'h2):(1'h0)]);
                  for (forvar1534 = (1'h0); (forvar1534 < (2'h2)); forvar1534 = (forvar1534 + (1'h1)))
                    begin
                      reg1535 <= reg1452[(2'h2):(1'h0)];
                    end
                  for (forvar1536 = (1'h0); (forvar1536 < (1'h1)); forvar1536 = (forvar1536 + (1'h1)))
                    begin
                      reg1537 <= $unsigned(reg1425[(1'h1):(1'h1)]);
                      reg1538 <= $unsigned((reg1454 ?
                          (&$signed(reg1423)) : ($signed(reg1444) * (~&wire1416))));
                    end
                end
            end
        end
      else
        begin
          for (forvar1482 = (1'h0); (forvar1482 < (1'h1)); forvar1482 = (forvar1482 + (1'h1)))
            begin
              if ($signed({forvar1418}))
                begin
                  if (reg1426)
                    begin
                      reg1483 <= reg1519[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1483 <= $signed($signed(((reg1426 ~^ reg1496) | (8'hab))));
                      reg1484 <= $unsigned((~&reg1418[(1'h0):(1'h0)]));
                      reg1485 <= reg1501[(3'h7):(3'h7)];
                    end
                  for (forvar1486 = (1'h0); (forvar1486 < (1'h1)); forvar1486 = (forvar1486 + (1'h1)))
                    begin
                      reg1487 <= ((+{forvar1417[(3'h6):(1'h0)]}) ^ $unsigned($signed((~reg1469))));
                      reg1488 <= ($unsigned(reg1505[(3'h4):(1'h0)]) != (reg1419[(1'h1):(1'h1)] ?
                          $unsigned(((8'hb1) ?
                              reg1500 : (8'ha9))) : ($signed(wire1415) > forvar1439[(1'h0):(1'h0)])));
                      reg1489 <= (~^(reg1476 ?
                          $unsigned($signed(reg1531)) : reg1419));
                      reg1490 <= (($signed(reg1515[(4'h9):(4'h8)]) ^ (reg1467 ?
                          ((8'hba) > forvar1450) : reg1468[(2'h2):(1'h0)])) > ((8'hba) | $unsigned($unsigned(reg1437))));
                    end
                  if ((($signed(reg1450[(3'h4):(1'h0)]) ?
                          (&{reg1459}) : reg1429[(4'ha):(3'h4)]) ?
                      forvar1439[(1'h0):(1'h0)] : (^~(forvar1518 ?
                          (reg1449 ?
                              reg1433 : forvar1450) : $unsigned((8'hb1))))))
                    begin
                      reg1491 <= ({$signed((reg1428 ? reg1462 : forvar1466))} ?
                          reg1423 : ({(reg1496 ^~ (8'ha8))} ?
                              reg1487 : ($unsigned((8'ha8)) ?
                                  {reg1430} : (wire1413 ?
                                      reg1485 : forvar1483))));
                      reg1492 <= $signed((~|((reg1512 ^~ forvar1514) ?
                          (reg1524 ? reg1451 : reg1447) : forvar1424)));
                      reg1493 <= $signed($unsigned({reg1532[(4'h9):(1'h1)]}));
                      reg1494 <= (((forvar1418[(4'hc):(4'hc)] ?
                              $signed(reg1484) : reg1479[(3'h4):(2'h2)]) << $signed(reg1417[(4'ha):(3'h5)])) ?
                          (^~(forvar1536 - reg1493[(3'h7):(1'h1)])) : (wire1412[(1'h0):(1'h0)] ?
                              (8'ha9) : (reg1499 ^ reg1428)));
                    end
                  else
                    begin
                      reg1491 <= ((reg1486 & ($unsigned(reg1465) <= reg1452[(2'h3):(2'h2)])) ?
                          reg1421[(3'h4):(3'h4)] : $unsigned((((8'ha3) ^~ forvar1536) ~^ $unsigned(reg1437))));
                      reg1492 <= ({reg1450} ?
                          ($signed({(8'ha5)}) ?
                              (8'h9f) : (8'ha3)) : $unsigned(reg1443));
                    end
                end
              else
                begin
                  for (forvar1483 = (1'h0); (forvar1483 < (1'h1)); forvar1483 = (forvar1483 + (1'h1)))
                    begin
                      reg1484 <= $signed({reg1455});
                      reg1485 <= reg1425[(3'h4):(1'h1)];
                    end
                  for (forvar1486 = (1'h0); (forvar1486 < (2'h3)); forvar1486 = (forvar1486 + (1'h1)))
                    begin
                      reg1487 <= reg1509;
                      reg1488 <= reg1481;
                      reg1489 <= (($unsigned($unsigned(reg1517)) + ((|forvar1518) ?
                              (^forvar1417) : (reg1436 <<< forvar1497))) ?
                          (((wire1415 && reg1471) <= (8'hb2)) ?
                              ((reg1529 ?
                                  reg1431 : reg1469) >> reg1434) : ((|reg1471) ?
                                  (~reg1502) : $unsigned(reg1456))) : ($unsigned((|(8'hb4))) ?
                              {$signed(reg1489)} : reg1472));
                    end
                  reg1490 <= (reg1538[(4'h9):(3'h5)] ^~ ($signed($signed((8'hb7))) * forvar1482));
                  reg1491 <= ({((reg1419 ?
                              forvar1439 : forvar1456) ^ reg1454)} ?
                      {{((8'ha9) ?
                                  reg1475 : (8'ha0))}} : ($unsigned((+reg1515)) << (+$unsigned(reg1469))));
                end
              if (reg1457)
                begin
                  if (($signed((reg1430 ?
                          $signed((8'hb0)) : (forvar1523 <= reg1446))) ?
                      reg1472 : (^$unsigned(((8'haf) <= reg1538)))))
                    begin
                      reg1495 <= $signed(reg1513[(2'h2):(1'h0)]);
                      reg1496 <= ({forvar1497[(4'hf):(2'h3)]} ?
                          reg1433[(2'h2):(1'h1)] : {reg1431});
                      reg1497 <= (((((8'h9d) ? (8'hb7) : forvar1456) ?
                              (|reg1472) : {reg1532}) <= reg1532) ?
                          (reg1475[(2'h2):(1'h0)] != reg1477[(2'h3):(2'h3)]) : (reg1423 ?
                              (reg1516[(1'h1):(1'h0)] ?
                                  $unsigned(reg1533) : (^~reg1454)) : $signed(reg1452)));
                      reg1498 <= (!(|{(reg1489 ? reg1448 : reg1427)}));
                    end
                  else
                    begin
                      reg1495 <= (reg1450 ?
                          reg1420 : $unsigned($signed((reg1531 ?
                              reg1512 : reg1524))));
                      reg1496 <= ($unsigned(((-forvar1486) ?
                              $signed(reg1488) : reg1435[(1'h0):(1'h0)])) ?
                          {$signed(reg1448[(2'h3):(2'h3)])} : ($signed(reg1538) ?
                              (~|reg1481[(1'h1):(1'h1)]) : reg1493[(4'ha):(4'ha)]));
                      reg1497 <= ($signed(forvar1490[(4'h9):(4'h8)]) < reg1452[(3'h5):(3'h5)]);
                      reg1498 <= $signed($unsigned((reg1536[(4'hc):(2'h3)] >> (!reg1429))));
                    end
                  reg1499 <= forvar1432[(2'h3):(2'h3)];
                  reg1500 <= $unsigned(((reg1520[(2'h3):(1'h0)] ?
                          forvar1427 : $signed(forvar1486)) ?
                      $signed((reg1503 ?
                          forvar1424 : reg1487)) : {(~^reg1424)}));
                end
              else
                begin
                  for (forvar1495 = (1'h0); (forvar1495 < (1'h1)); forvar1495 = (forvar1495 + (1'h1)))
                    begin
                      reg1496 <= $signed(reg1501[(4'hc):(1'h1)]);
                      reg1497 <= reg1537;
                    end
                  for (forvar1498 = (1'h0); (forvar1498 < (2'h3)); forvar1498 = (forvar1498 + (1'h1)))
                    begin
                      reg1499 <= (reg1499 ?
                          {((reg1435 <<< reg1471) ~^ reg1430)} : {(((8'h9c) ~^ forvar1514) ?
                                  (wire1416 + reg1508) : (reg1441 ?
                                      reg1486 : reg1430))});
                    end
                end
              for (forvar1501 = (1'h0); (forvar1501 < (2'h3)); forvar1501 = (forvar1501 + (1'h1)))
                begin
                  for (forvar1502 = (1'h0); (forvar1502 < (1'h1)); forvar1502 = (forvar1502 + (1'h1)))
                    begin
                      reg1503 <= reg1486;
                      reg1504 <= forvar1518;
                    end
                end
            end
        end
    end
  module1540 #() modinst2028 (wire2027, clk, reg1520, wire1412, reg1535, reg1501, reg1469);
  assign wire2029 = {(&(reg1485 || (8'hb1)))};
  assign wire2030 = (reg1500 ?
                        ($unsigned(reg1486) + (reg1424 ?
                            $signed((8'ha8)) : (+reg1526))) : ($signed(reg1425) & (|(reg1491 ?
                            reg1515 : reg1532))));
  assign wire2031 = $unsigned($unsigned(reg1526));
  always
    @(posedge clk) begin
      if ($unsigned((~((reg1498 ?
          reg1448 : reg1533) & reg1484[(3'h5):(2'h3)]))))
        begin
          for (forvar2032 = (1'h0); (forvar2032 < (1'h0)); forvar2032 = (forvar2032 + (1'h1)))
            begin
              reg2033 <= $signed(reg1496);
            end
          for (forvar2034 = (1'h0); (forvar2034 < (1'h0)); forvar2034 = (forvar2034 + (1'h1)))
            begin
              for (forvar2035 = (1'h0); (forvar2035 < (1'h0)); forvar2035 = (forvar2035 + (1'h1)))
                begin
                  for (forvar2036 = (1'h0); (forvar2036 < (1'h1)); forvar2036 = (forvar2036 + (1'h1)))
                    begin
                      reg2037 <= reg1434[(2'h2):(2'h2)];
                      reg2038 <= ((($unsigned(reg1527) + $unsigned(reg1495)) ?
                          {(reg1489 ?
                                  wire1414 : reg1436)} : reg1506[(4'h9):(1'h0)]) && (~(reg1435 >> (reg1473 > reg1484))));
                      reg2039 <= reg1459[(2'h3):(2'h2)];
                      reg2040 <= $unsigned((8'hb1));
                    end
                  if (((({reg1447} == (8'ha4)) ?
                          ($unsigned(reg1427) == {reg1472}) : $unsigned(((8'ha1) < reg1524))) ?
                      (reg1490 ?
                          (^~$unsigned((8'hb6))) : (|(reg1492 - reg1502))) : reg1457[(2'h2):(1'h1)]))
                    begin
                      reg2041 <= {(~&($signed(reg1499) - ((8'had) >>> (8'ha6))))};
                      reg2042 <= (^~((reg1487 << reg1486[(2'h3):(2'h2)]) ?
                          wire2030 : reg1434[(3'h7):(3'h5)]));
                      reg2043 <= reg1507;
                    end
                  else
                    begin
                      reg2041 <= ((-((reg1467 >> (8'hab)) ?
                          $unsigned(reg1430) : forvar2032)) < $unsigned(((~|reg1429) >>> wire2031[(1'h0):(1'h0)])));
                      reg2042 <= $signed(reg1423[(1'h0):(1'h0)]);
                      reg2043 <= {(&$unsigned(reg1445))};
                    end
                end
              for (forvar2044 = (1'h0); (forvar2044 < (2'h2)); forvar2044 = (forvar2044 + (1'h1)))
                begin
                  reg2045 <= (~^((^{reg1535}) ?
                      (~&{reg1530}) : (-$unsigned(reg1473))));
                  if (reg1492[(4'h9):(3'h6)])
                    begin
                      reg2046 <= $unsigned({({reg1530} << ((8'hab) ?
                              reg1425 : reg1448))});
                      reg2047 <= (reg1475 ? reg1513 : $signed((+wire1414)));
                      reg2048 <= ($signed(reg1446[(1'h0):(1'h0)]) ?
                          reg1423[(1'h1):(1'h0)] : reg1462[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg2046 <= (reg1511[(2'h3):(1'h1)] ?
                          (~^forvar2036[(1'h1):(1'h0)]) : (!(8'haa)));
                      reg2047 <= $unsigned(((!$signed(reg1531)) ?
                          $unsigned(reg2043) : ($unsigned(reg1447) ?
                              (reg1449 ?
                                  reg1461 : reg2048) : $unsigned((8'ha6)))));
                    end
                  for (forvar2049 = (1'h0); (forvar2049 < (2'h2)); forvar2049 = (forvar2049 + (1'h1)))
                    begin
                      reg2050 <= $signed(reg2037);
                      reg2051 <= $unsigned((($signed(reg1463) ?
                              $unsigned(reg1460) : (~|reg1450)) ?
                          reg1524 : (8'had)));
                      reg2052 <= {$unsigned(forvar2035[(4'h9):(1'h1)])};
                    end
                end
            end
          reg2053 <= $unsigned((reg1485[(1'h1):(1'h0)] ?
              $unsigned((~^reg1449)) : (8'haf)));
          for (forvar2054 = (1'h0); (forvar2054 < (1'h1)); forvar2054 = (forvar2054 + (1'h1)))
            begin
              for (forvar2055 = (1'h0); (forvar2055 < (2'h3)); forvar2055 = (forvar2055 + (1'h1)))
                begin
                  for (forvar2056 = (1'h0); (forvar2056 < (2'h2)); forvar2056 = (forvar2056 + (1'h1)))
                    begin
                      reg2057 <= reg1537[(1'h1):(1'h1)];
                    end
                  if (($unsigned(reg1495) && $signed($unsigned((8'hb5)))))
                    begin
                      reg2058 <= $signed((|{(reg1534 & reg1538)}));
                    end
                  else
                    begin
                      reg2058 <= $signed($signed($unsigned($signed(reg1453))));
                      reg2059 <= forvar2044[(4'hf):(4'hf)];
                      reg2060 <= ($signed((~^$unsigned(reg1503))) == (reg1498[(3'h5):(2'h3)] <<< (-(reg1490 ?
                          (8'hb7) : reg2038))));
                      reg2061 <= ($unsigned((reg1484 ?
                          (reg1491 ?
                              reg1509 : reg1435) : reg1477[(4'h8):(3'h5)])) || $unsigned(reg1447));
                    end
                  for (forvar2062 = (1'h0); (forvar2062 < (1'h0)); forvar2062 = (forvar2062 + (1'h1)))
                    begin
                      reg2063 <= reg1525;
                      reg2064 <= (+$unsigned(((wire1414 ? (8'ha0) : reg1485) ?
                          reg1463[(1'h0):(1'h0)] : (8'ha7))));
                      reg2065 <= $unsigned($signed(((reg1521 ?
                              reg1478 : reg1445) ?
                          $unsigned(wire1412) : reg1527)));
                      reg2066 <= (&$signed({$signed(reg1472)}));
                    end
                end
            end
        end
      else
        begin
          for (forvar2032 = (1'h0); (forvar2032 < (1'h0)); forvar2032 = (forvar2032 + (1'h1)))
            begin
              for (forvar2033 = (1'h0); (forvar2033 < (2'h2)); forvar2033 = (forvar2033 + (1'h1)))
                begin
                  for (forvar2034 = (1'h0); (forvar2034 < (1'h1)); forvar2034 = (forvar2034 + (1'h1)))
                    begin
                      reg2035 <= reg1440;
                      reg2036 <= ($signed($signed(reg1508)) ?
                          (!$signed((!reg2047))) : $unsigned((!{reg1445})));
                      reg2037 <= reg1515[(3'h4):(1'h1)];
                      reg2038 <= ((forvar2032 ?
                          $unsigned($unsigned(reg1479)) : $unsigned((|reg2058))) + (+reg1473[(3'h4):(2'h3)]));
                    end
                end
              for (forvar2039 = (1'h0); (forvar2039 < (2'h3)); forvar2039 = (forvar2039 + (1'h1)))
                begin
                  for (forvar2040 = (1'h0); (forvar2040 < (1'h1)); forvar2040 = (forvar2040 + (1'h1)))
                    begin
                      reg2041 <= (~&$unsigned(((reg1428 ?
                          forvar2040 : reg1438) < (reg1497 <<< reg1492))));
                      reg2042 <= reg2060[(1'h1):(1'h1)];
                      reg2043 <= $signed((8'hb9));
                    end
                  for (forvar2044 = (1'h0); (forvar2044 < (2'h2)); forvar2044 = (forvar2044 + (1'h1)))
                    begin
                      reg2045 <= $signed(((reg1465[(1'h0):(1'h0)] >= reg1456[(1'h0):(1'h0)]) ?
                          reg1443 : reg2035[(1'h1):(1'h0)]));
                      reg2046 <= reg1436[(4'hc):(4'hc)];
                      reg2047 <= ((-(((8'ha9) ? reg1433 : reg1428) ?
                          ((8'hb5) <= reg2065) : $unsigned(reg1537))) && ($signed($unsigned(reg1539)) ?
                          (^~reg1437) : $signed(forvar2044)));
                    end
                  for (forvar2048 = (1'h0); (forvar2048 < (1'h1)); forvar2048 = (forvar2048 + (1'h1)))
                    begin
                      reg2049 <= $signed((reg1426 ?
                          (~^$unsigned(reg1434)) : $unsigned((~^reg1479))));
                      reg2050 <= reg2059[(2'h2):(1'h0)];
                    end
                end
              if ($unsigned($signed($signed((^(8'hb6))))))
                begin
                  reg2051 <= $unsigned($signed({reg2057}));
                  for (forvar2052 = (1'h0); (forvar2052 < (2'h2)); forvar2052 = (forvar2052 + (1'h1)))
                    begin
                      reg2053 <= $unsigned(((-(forvar2044 ?
                              (8'hae) : reg1517)) ?
                          ($signed((8'hac)) << (reg2045 ?
                              reg1469 : reg1450)) : $unsigned((!reg1501))));
                      reg2054 <= $signed((((~forvar2062) | reg1431[(3'h4):(2'h2)]) * reg1434[(4'h8):(3'h7)]));
                      reg2055 <= reg1514;
                    end
                  for (forvar2056 = (1'h0); (forvar2056 < (2'h2)); forvar2056 = (forvar2056 + (1'h1)))
                    begin
                      reg2057 <= (($signed(reg2038) ?
                          $unsigned($signed(forvar2033)) : $signed($unsigned(reg1442))) & reg1539[(1'h0):(1'h0)]);
                      reg2058 <= ($unsigned((!reg2065[(4'hb):(1'h1)])) ?
                          reg2060 : reg1464);
                      reg2059 <= forvar2062[(2'h3):(1'h0)];
                      reg2060 <= $signed((&reg1464));
                    end
                  for (forvar2061 = (1'h0); (forvar2061 < (1'h1)); forvar2061 = (forvar2061 + (1'h1)))
                    begin
                      reg2062 <= {reg1505};
                    end
                end
              else
                begin
                  for (forvar2051 = (1'h0); (forvar2051 < (2'h3)); forvar2051 = (forvar2051 + (1'h1)))
                    begin
                      reg2052 <= reg1512[(2'h3):(1'h1)];
                      reg2053 <= (((reg1507 + $unsigned(reg2045)) ?
                              (~&(+reg1491)) : reg1526[(2'h3):(1'h1)]) ?
                          ((reg2049 >> (|reg2040)) ?
                              (!forvar2055[(1'h1):(1'h1)]) : $unsigned({wire2031})) : (($signed((8'haa)) ?
                              (forvar2061 ?
                                  forvar2040 : reg1419) : $signed(reg1463)) <<< (|(forvar2033 ?
                              forvar2062 : reg1454))));
                    end
                  for (forvar2054 = (1'h0); (forvar2054 < (1'h1)); forvar2054 = (forvar2054 + (1'h1)))
                    begin
                      reg2055 <= reg1444;
                      reg2056 <= reg1485;
                      reg2057 <= (reg1492[(2'h2):(1'h0)] + ((reg1440[(2'h2):(2'h2)] ^ $signed(reg1440)) ?
                          reg1467 : $unsigned((~^reg1490))));
                    end
                  if ({$unsigned(reg2049[(3'h5):(3'h5)])})
                    begin
                      reg2058 <= $unsigned($unsigned(((forvar2040 <<< reg1447) ?
                          (reg1437 ? reg1432 : reg1489) : (reg1454 ?
                              reg1483 : forvar2040))));
                      reg2059 <= $unsigned($signed((reg2039 ?
                          $unsigned(reg1479) : (forvar2033 ^ reg1487))));
                      reg2060 <= (|reg2045[(2'h2):(1'h1)]);
                      reg2061 <= ((~^reg1497[(4'he):(4'hd)]) < ((reg1433[(2'h2):(1'h1)] ?
                              reg1472 : wire1416[(3'h5):(2'h2)]) ?
                          ($unsigned(reg2041) || ((8'hb4) ?
                              reg1524 : forvar2033)) : forvar2051[(5'h10):(4'hf)]));
                    end
                  else
                    begin
                      reg2058 <= (~&$unsigned((reg1515 >= $signed(reg1435))));
                      reg2059 <= ((~reg1423) - {(~&{reg1417})});
                    end
                end
              if (reg1423)
                begin
                  reg2063 <= ((((reg1426 ? forvar2035 : (8'ha2)) ?
                          $signed(reg1432) : reg2043[(3'h4):(2'h2)]) * (8'had)) ?
                      ($signed((reg1455 || reg1481)) ?
                          $unsigned((reg2046 ?
                              reg1519 : forvar2054)) : (~|$signed(reg1485))) : ($signed((~|reg1482)) ^ {((8'haf) + reg1475)}));
                  for (forvar2064 = (1'h0); (forvar2064 < (2'h2)); forvar2064 = (forvar2064 + (1'h1)))
                    begin
                      reg2065 <= $unsigned(reg1460);
                      reg2066 <= ((8'hb7) <= (~|$signed($unsigned(reg1445))));
                    end
                end
              else
                begin
                  reg2063 <= $signed($unsigned((^~$signed(reg1420))));
                  if (({(^$signed((8'ha0)))} | reg1493))
                    begin
                      reg2064 <= reg2046;
                      reg2065 <= reg1489;
                    end
                  else
                    begin
                      reg2064 <= $signed($signed($signed((reg1437 + forvar2040))));
                      reg2065 <= (^($signed(reg1492[(1'h0):(1'h0)]) << ($signed(reg2052) ?
                          $signed(reg1499) : (~&reg1420))));
                      reg2066 <= $signed({{(^~reg1524)}});
                      reg2067 <= forvar2061;
                    end
                end
            end
          reg2068 <= reg2055[(4'he):(4'hb)];
        end
      if (((~^({reg1441} <<< $unsigned((8'hb8)))) >>> {(8'hba)}))
        begin
          if (forvar2055)
            begin
              for (forvar2069 = (1'h0); (forvar2069 < (2'h2)); forvar2069 = (forvar2069 + (1'h1)))
                begin
                  reg2070 <= $signed((~|$signed((&reg1432))));
                end
              reg2071 <= reg1425;
              if ((((forvar2044[(3'h4):(1'h1)] ? (8'ha1) : reg1471) ?
                      {reg2047} : ($unsigned(forvar2034) != (reg1426 ?
                          reg1444 : reg1529))) ?
                  $unsigned($unsigned((forvar2048 <= forvar2061))) : $unsigned(forvar2052[(3'h5):(3'h5)])))
                begin
                  for (forvar2072 = (1'h0); (forvar2072 < (2'h3)); forvar2072 = (forvar2072 + (1'h1)))
                    begin
                      reg2073 <= (forvar2069[(2'h3):(2'h3)] ?
                          ((8'h9c) ?
                              {(&reg2062)} : reg1424[(1'h0):(1'h0)]) : reg2067);
                      reg2074 <= (wire2030 ?
                          (~(reg1448 & (|reg1534))) : (forvar2069 ?
                              $unsigned(reg1490[(3'h5):(1'h0)]) : (~&(forvar2040 != reg2051))));
                    end
                  if ((~reg2064[(2'h2):(1'h0)]))
                    begin
                      reg2075 <= reg1422[(2'h2):(1'h0)];
                      reg2076 <= $unsigned(((reg1444[(3'h4):(1'h0)] == $unsigned(reg1527)) && ($signed((8'ha2)) ?
                          $unsigned(reg1512) : (|reg1505))));
                      reg2077 <= (&reg1493);
                      reg2078 <= (^~reg1490[(3'h7):(3'h6)]);
                    end
                  else
                    begin
                      reg2075 <= ((reg1503[(2'h2):(1'h1)] ?
                          ((reg2078 & reg1421) ?
                              (&reg2041) : (reg1442 ?
                                  reg2074 : reg1494)) : reg1508) <<< ({$signed(reg1514)} ?
                          reg2060[(2'h2):(1'h1)] : (~&$signed(reg1538))));
                      reg2076 <= (~&({((8'hba) ?
                              forvar2051 : reg1443)} <= (reg1471 || (~reg1446))));
                      reg2077 <= (reg1486 >>> $unsigned(((reg1455 ?
                              reg2057 : reg1475) ?
                          {reg2051} : {reg1537})));
                      reg2078 <= reg2043;
                    end
                  if (reg1504)
                    begin
                      reg2079 <= (|$signed(reg2062));
                      reg2080 <= reg1496;
                      reg2081 <= ({{$signed(reg1468)}} > reg1480[(3'h4):(1'h1)]);
                      reg2082 <= (^$unsigned({$unsigned((8'ha5))}));
                    end
                  else
                    begin
                      reg2079 <= (8'h9c);
                      reg2080 <= reg1501[(4'he):(3'h4)];
                    end
                  reg2083 <= wire1414;
                end
              else
                begin
                  if ((^$signed(reg2082)))
                    begin
                      reg2072 <= (8'hb7);
                      reg2073 <= (forvar2034 ?
                          reg1438 : $signed(reg1513[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg2072 <= $unsigned((|(reg1497 ^ (reg2068 ?
                          reg1529 : reg2043))));
                      reg2073 <= $signed(reg1501[(4'hf):(4'hb)]);
                      reg2074 <= forvar2061[(3'h4):(2'h3)];
                      reg2075 <= {(~&(^forvar2061))};
                    end
                  for (forvar2076 = (1'h0); (forvar2076 < (1'h1)); forvar2076 = (forvar2076 + (1'h1)))
                    begin
                      reg2077 <= $signed((|{$signed(reg2039)}));
                      reg2078 <= $signed(($signed((reg1479 < reg2071)) == wire2029[(2'h3):(2'h2)]));
                    end
                end
            end
          else
            begin
              reg2069 <= (($signed(reg1536[(4'ha):(1'h1)]) != reg1531[(4'h8):(1'h1)]) ?
                  (8'hb8) : reg2062[(3'h6):(1'h1)]);
              for (forvar2070 = (1'h0); (forvar2070 < (2'h2)); forvar2070 = (forvar2070 + (1'h1)))
                begin
                  if (((^~reg1432) - ($signed((-reg2067)) * reg1422[(2'h2):(1'h0)])))
                    begin
                      reg2071 <= reg1418;
                      reg2072 <= forvar2072;
                      reg2073 <= ((wire1415 ?
                          reg1532 : (8'h9f)) ^~ $signed(reg2072[(2'h3):(2'h2)]));
                      reg2074 <= reg1487;
                    end
                  else
                    begin
                      reg2071 <= $unsigned((+$signed($unsigned(reg2080))));
                      reg2072 <= $signed((reg2071[(1'h1):(1'h1)] ?
                          reg1479 : reg1516[(4'hc):(4'hb)]));
                      reg2073 <= forvar2076;
                      reg2074 <= {($unsigned($unsigned(reg2064)) ?
                              (reg2045[(2'h2):(2'h2)] ?
                                  reg1447 : (~&reg2045)) : $unsigned((+reg1481)))};
                    end
                end
              for (forvar2075 = (1'h0); (forvar2075 < (1'h0)); forvar2075 = (forvar2075 + (1'h1)))
                begin
                  for (forvar2076 = (1'h0); (forvar2076 < (2'h2)); forvar2076 = (forvar2076 + (1'h1)))
                    begin
                      reg2077 <= {$unsigned(((|reg1444) ?
                              (-forvar2051) : $signed(forvar2062)))};
                    end
                  for (forvar2078 = (1'h0); (forvar2078 < (1'h1)); forvar2078 = (forvar2078 + (1'h1)))
                    begin
                      reg2079 <= reg2059;
                      reg2080 <= reg1516;
                    end
                end
              if ((~|reg2076[(1'h0):(1'h0)]))
                begin
                  for (forvar2081 = (1'h0); (forvar2081 < (1'h0)); forvar2081 = (forvar2081 + (1'h1)))
                    begin
                      reg2082 <= (^(reg2083[(3'h4):(2'h3)] ?
                          (&reg2080[(4'h8):(3'h6)]) : (((8'hb3) - (8'hb0)) ~^ (reg1461 ?
                              reg1505 : (8'hb8)))));
                    end
                end
              else
                begin
                  for (forvar2081 = (1'h0); (forvar2081 < (1'h0)); forvar2081 = (forvar2081 + (1'h1)))
                    begin
                      reg2082 <= ($signed((^~(^reg2080))) ?
                          ((-$unsigned(forvar2061)) * reg1486) : $unsigned(({reg2046} ?
                              ((8'had) ? reg1460 : (8'hae)) : (~^reg1531))));
                      reg2083 <= (~&($signed((!reg2078)) >>> {reg1502}));
                      reg2084 <= {reg2081};
                      reg2085 <= {$unsigned($unsigned({forvar2044}))};
                    end
                end
            end
          for (forvar2086 = (1'h0); (forvar2086 < (2'h3)); forvar2086 = (forvar2086 + (1'h1)))
            begin
              for (forvar2087 = (1'h0); (forvar2087 < (2'h3)); forvar2087 = (forvar2087 + (1'h1)))
                begin
                  if ({$signed($signed({forvar2040}))})
                    begin
                      reg2088 <= $signed(reg1465);
                      reg2089 <= (-$unsigned({$signed(forvar2039)}));
                    end
                  else
                    begin
                      reg2088 <= (~|reg2082);
                      reg2089 <= reg2048;
                      reg2090 <= reg1482;
                    end
                  for (forvar2091 = (1'h0); (forvar2091 < (2'h3)); forvar2091 = (forvar2091 + (1'h1)))
                    begin
                      reg2092 <= ((reg1441 ?
                          {$signed(reg1422)} : reg1525) >> reg1447[(1'h1):(1'h0)]);
                    end
                  if ($signed($unsigned(reg2082)))
                    begin
                      reg2093 <= reg2045[(1'h1):(1'h1)];
                      reg2094 <= $unsigned(forvar2032[(4'hd):(3'h5)]);
                    end
                  else
                    begin
                      reg2093 <= ((reg1535[(4'hc):(4'ha)] ?
                              (^(reg1495 ?
                                  (8'hb3) : reg1527)) : ($signed(reg1432) != $signed(reg1467))) ?
                          ($signed(reg2083[(2'h2):(2'h2)]) ?
                              reg1434[(1'h0):(1'h0)] : $signed({reg1495})) : (+{$unsigned((8'h9c))}));
                      reg2094 <= (((8'h9f) ^~ (-$unsigned(forvar2049))) ^~ $signed((~^(&(8'hb7)))));
                    end
                end
            end
          for (forvar2095 = (1'h0); (forvar2095 < (2'h3)); forvar2095 = (forvar2095 + (1'h1)))
            begin
              for (forvar2096 = (1'h0); (forvar2096 < (1'h1)); forvar2096 = (forvar2096 + (1'h1)))
                begin
                  for (forvar2097 = (1'h0); (forvar2097 < (1'h0)); forvar2097 = (forvar2097 + (1'h1)))
                    begin
                      reg2098 <= reg2079;
                    end
                  if (reg1481)
                    begin
                      reg2099 <= $unsigned($unsigned(((reg1430 ?
                          reg2045 : forvar2091) ^ $signed(reg1435))));
                      reg2100 <= reg1536;
                    end
                  else
                    begin
                      reg2099 <= {reg1532[(4'h9):(2'h3)]};
                    end
                  for (forvar2101 = (1'h0); (forvar2101 < (2'h2)); forvar2101 = (forvar2101 + (1'h1)))
                    begin
                      reg2102 <= ((!((~^reg1418) && $unsigned(reg1478))) <= (reg2088[(3'h4):(1'h1)] - reg2039[(3'h7):(1'h1)]));
                      reg2103 <= {(reg1421 << reg1463[(2'h2):(2'h2)])};
                      reg2104 <= (~$signed(reg2083));
                      reg2105 <= (-($signed((-reg2071)) * reg1486[(4'hb):(3'h6)]));
                    end
                end
            end
        end
      else
        begin
          if ((reg1421[(2'h2):(1'h0)] ^ $unsigned($unsigned(reg1437[(4'ha):(3'h5)]))))
            begin
              reg2069 <= ((((~|(8'hba)) ?
                      (forvar2044 ?
                          forvar2064 : forvar2035) : (forvar2044 + reg1497)) ?
                  reg1487 : ({reg2058} ?
                      (~&reg2046) : reg2100)) != reg1517[(5'h10):(4'h9)]);
              for (forvar2070 = (1'h0); (forvar2070 < (1'h1)); forvar2070 = (forvar2070 + (1'h1)))
                begin
                  reg2071 <= reg1531;
                  for (forvar2072 = (1'h0); (forvar2072 < (1'h1)); forvar2072 = (forvar2072 + (1'h1)))
                    begin
                      reg2073 <= {reg1483[(1'h0):(1'h0)]};
                      reg2074 <= (&(|(reg1464 ?
                          forvar2091[(3'h5):(3'h5)] : (~&reg1462))));
                      reg2075 <= $signed((8'ha6));
                      reg2076 <= forvar2078;
                    end
                  for (forvar2077 = (1'h0); (forvar2077 < (2'h3)); forvar2077 = (forvar2077 + (1'h1)))
                    begin
                      reg2078 <= reg1464;
                      reg2079 <= (reg2047 ?
                          $signed(($unsigned(reg2067) ?
                              reg1527[(2'h2):(1'h0)] : (reg2073 >>> (8'hb8)))) : (8'h9d));
                      reg2080 <= $signed(forvar2076[(1'h0):(1'h0)]);
                    end
                end
            end
          else
            begin
              if (reg1480)
                begin
                  if (reg1488)
                    begin
                      reg2069 <= $signed(({reg1462} ^~ $unsigned((8'ha1))));
                      reg2070 <= ((reg2071 ?
                              reg1485[(3'h7):(3'h5)] : (^forvar2062[(2'h2):(1'h0)])) ?
                          $unsigned(reg1520[(1'h0):(1'h0)]) : reg2061[(2'h2):(2'h2)]);
                      reg2071 <= reg1437;
                      reg2072 <= reg1530;
                    end
                  else
                    begin
                      reg2069 <= forvar2064[(4'h9):(3'h4)];
                    end
                  if (reg2098)
                    begin
                      reg2073 <= reg1488;
                      reg2074 <= (((^~(reg1513 && forvar2044)) ?
                          {$unsigned((8'ha4))} : wire2027) && (&((reg2054 ?
                          reg2069 : reg1487) != (~^(8'hb1)))));
                    end
                  else
                    begin
                      reg2073 <= $signed(reg1538[(4'h8):(3'h6)]);
                      reg2074 <= ($signed((!((8'ha3) || reg1500))) ?
                          (&((reg1496 - reg2082) == (reg1519 ?
                              reg2056 : reg1465))) : ((-$unsigned(reg1446)) ?
                              $unsigned((reg1432 <= forvar2095)) : $unsigned((reg1486 + reg2058))));
                      reg2075 <= wire2027[(1'h0):(1'h0)];
                      reg2076 <= (reg1529[(4'hb):(4'hb)] ?
                          ((forvar2097 ~^ (reg1495 ? forvar2078 : reg1459)) ?
                              (~|reg1530) : ((reg1450 ?
                                  forvar2097 : reg2036) >= $signed(reg1516))) : {{(reg2065 ?
                                      reg1447 : reg1438)}});
                    end
                end
              else
                begin
                  reg2069 <= forvar2054[(1'h1):(1'h1)];
                  for (forvar2070 = (1'h0); (forvar2070 < (2'h2)); forvar2070 = (forvar2070 + (1'h1)))
                    begin
                      reg2071 <= $unsigned(reg1432);
                      reg2072 <= (~^reg1432[(4'hb):(2'h2)]);
                      reg2073 <= (!($unsigned($unsigned(reg2071)) ?
                          {$unsigned(reg1434)} : $signed((reg1458 && forvar2039))));
                    end
                  if ($unsigned((|(reg2100 ?
                      reg1463[(3'h5):(2'h3)] : $unsigned((8'hb3))))))
                    begin
                      reg2074 <= ((8'hb0) << ($signed($unsigned(reg1446)) + (reg2045[(2'h2):(2'h2)] ?
                          (~^reg2047) : reg2042[(1'h1):(1'h1)])));
                      reg2075 <= ((^~$signed($signed(reg1532))) ?
                          (^$signed(forvar2033)) : $signed(reg1446[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg2074 <= reg1506;
                    end
                  if ($unsigned($unsigned(((^~forvar2072) ?
                      $unsigned(reg2045) : (~&reg1440)))))
                    begin
                      reg2076 <= ({(8'ha5)} > $signed($signed(reg1437)));
                      reg2077 <= $unsigned((~^$unsigned(reg1522[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg2076 <= $unsigned(forvar2101[(1'h1):(1'h0)]);
                    end
                end
              if (((((reg1471 == reg2037) && $unsigned(reg2068)) ?
                  forvar2061 : $signed(reg1434)) & forvar2101))
                begin
                  for (forvar2078 = (1'h0); (forvar2078 < (1'h0)); forvar2078 = (forvar2078 + (1'h1)))
                    begin
                      reg2079 <= forvar2032[(4'he):(4'hd)];
                      reg2080 <= reg2094;
                      reg2081 <= ((reg1522[(1'h1):(1'h0)] ?
                          $signed(reg1462[(2'h2):(1'h1)]) : (~^{reg1464})) >= $signed(((reg2074 ?
                          reg2033 : reg1499) & (!reg2082))));
                    end
                  reg2082 <= reg1456;
                end
              else
                begin
                  if ((~&reg1452))
                    begin
                      reg2078 <= $signed({($signed(reg2046) && ((8'ha3) ?
                              wire2030 : reg1436))});
                    end
                  else
                    begin
                      reg2078 <= {($signed(reg1473) ? (^~(8'hb2)) : reg1450)};
                      reg2079 <= $unsigned((^$unsigned($signed(reg1465))));
                      reg2080 <= ($unsigned(((8'hb2) && (reg1441 || reg1481))) - (+(~&$unsigned((8'hb9)))));
                      reg2081 <= ((!reg1526) - $unsigned((reg2067 <= $unsigned((8'hae)))));
                    end
                  for (forvar2082 = (1'h0); (forvar2082 < (2'h2)); forvar2082 = (forvar2082 + (1'h1)))
                    begin
                      reg2083 <= $unsigned(($unsigned((~reg1509)) ?
                          {$signed(reg1517)} : (8'ha0)));
                      reg2084 <= reg2051[(3'h6):(2'h2)];
                    end
                  for (forvar2085 = (1'h0); (forvar2085 < (2'h3)); forvar2085 = (forvar2085 + (1'h1)))
                    begin
                      reg2086 <= $signed((^~$unsigned($unsigned(wire1414))));
                      reg2087 <= forvar2034;
                      reg2088 <= $unsigned({$unsigned({reg1469})});
                      reg2089 <= (reg2057[(2'h3):(1'h1)] ?
                          $unsigned(((forvar2078 || reg1421) ?
                              reg1488[(2'h3):(1'h1)] : (reg2103 ?
                                  reg2051 : (8'hae)))) : {wire2030[(2'h3):(1'h0)]});
                    end
                end
              for (forvar2090 = (1'h0); (forvar2090 < (2'h3)); forvar2090 = (forvar2090 + (1'h1)))
                begin
                  for (forvar2091 = (1'h0); (forvar2091 < (2'h2)); forvar2091 = (forvar2091 + (1'h1)))
                    begin
                      reg2092 <= (^reg1434[(3'h6):(1'h0)]);
                    end
                  for (forvar2093 = (1'h0); (forvar2093 < (1'h1)); forvar2093 = (forvar2093 + (1'h1)))
                    begin
                      reg2094 <= (&$signed($unsigned($signed(reg2042))));
                      reg2095 <= {{((!reg2083) && reg1451[(4'h8):(3'h6)])}};
                    end
                  for (forvar2096 = (1'h0); (forvar2096 < (2'h2)); forvar2096 = (forvar2096 + (1'h1)))
                    begin
                      reg2097 <= reg2061;
                      reg2098 <= reg2050[(3'h4):(3'h4)];
                      reg2099 <= ($signed((~&reg2038[(3'h4):(1'h0)])) ?
                          ({{reg1519}} <<< {reg2042[(2'h3):(2'h2)]}) : $signed($unsigned((reg2047 ?
                              reg1449 : reg2045))));
                      reg2100 <= (~&(8'hb8));
                    end
                end
            end
          for (forvar2101 = (1'h0); (forvar2101 < (2'h3)); forvar2101 = (forvar2101 + (1'h1)))
            begin
              reg2102 <= ($signed($signed($signed(reg2058))) < wire2029);
              for (forvar2103 = (1'h0); (forvar2103 < (2'h2)); forvar2103 = (forvar2103 + (1'h1)))
                begin
                  reg2104 <= $signed(reg1527);
                  for (forvar2105 = (1'h0); (forvar2105 < (1'h0)); forvar2105 = (forvar2105 + (1'h1)))
                    begin
                      reg2106 <= wire2029;
                      reg2107 <= {forvar2093[(3'h6):(3'h4)]};
                    end
                end
              reg2108 <= ({reg1514[(2'h2):(1'h1)]} ?
                  (|$signed($unsigned(reg1441))) : ({$signed((8'ha4))} >>> $unsigned($signed((8'haa)))));
              for (forvar2109 = (1'h0); (forvar2109 < (2'h3)); forvar2109 = (forvar2109 + (1'h1)))
                begin
                  if (wire1412)
                    begin
                      reg2110 <= ($unsigned($signed($signed(reg1519))) ?
                          $signed($unsigned((~&reg1461))) : reg2065);
                      reg2111 <= reg1531;
                      reg2112 <= reg1432[(1'h1):(1'h0)];
                      reg2113 <= (~&((|$signed(reg1516)) ?
                          (reg1455[(2'h2):(1'h0)] + reg1430) : $signed((8'h9f))));
                    end
                  else
                    begin
                      reg2110 <= {(^((|reg1426) <= (reg1429 ?
                              reg1468 : reg1476)))};
                      reg2111 <= reg2098;
                      reg2112 <= (+{(~^(reg2106 ? (8'hb8) : reg2077))});
                    end
                  for (forvar2114 = (1'h0); (forvar2114 < (1'h1)); forvar2114 = (forvar2114 + (1'h1)))
                    begin
                      reg2115 <= ($signed({(~&reg1514)}) >> {reg1538[(3'h4):(2'h2)]});
                      reg2116 <= $unsigned(reg2055[(2'h2):(1'h0)]);
                      reg2117 <= (({$unsigned(reg1506)} ?
                          {reg1458[(2'h2):(1'h1)]} : ((8'hb7) <= $signed(reg2051))) >= (+$unsigned((reg1417 && (8'ha6)))));
                    end
                end
            end
        end
      if ((&(^~reg1506[(4'h9):(3'h5)])))
        begin
          reg2118 <= ($signed((8'ha0)) <= (wire1413 << $unsigned((~&(8'hba)))));
          for (forvar2119 = (1'h0); (forvar2119 < (1'h1)); forvar2119 = (forvar2119 + (1'h1)))
            begin
              if ((reg1427[(1'h1):(1'h1)] ?
                  ($signed((^reg1476)) <= (reg2100 - (reg1479 && reg1514))) : (^(reg2038[(4'h9):(3'h7)] ?
                      ((8'hab) >> forvar2062) : $signed(reg2115)))))
                begin
                  for (forvar2120 = (1'h0); (forvar2120 < (2'h3)); forvar2120 = (forvar2120 + (1'h1)))
                    begin
                      reg2121 <= ((!({reg2116} + $unsigned(reg1536))) ?
                          (reg2117 ?
                              {(-reg1501)} : reg2081[(3'h6):(1'h0)]) : {($unsigned(forvar2120) ^ {forvar2101})});
                      reg2122 <= (8'haf);
                      reg2123 <= reg1484;
                    end
                  for (forvar2124 = (1'h0); (forvar2124 < (2'h3)); forvar2124 = (forvar2124 + (1'h1)))
                    begin
                      reg2125 <= reg1502;
                      reg2126 <= $signed(reg2059);
                    end
                  for (forvar2127 = (1'h0); (forvar2127 < (2'h2)); forvar2127 = (forvar2127 + (1'h1)))
                    begin
                      reg2128 <= reg2043;
                      reg2129 <= reg1420[(4'ha):(1'h0)];
                      reg2130 <= (reg1476[(1'h1):(1'h0)] ?
                          $signed((!(reg2051 ?
                              reg1459 : reg1498))) : reg1524[(1'h1):(1'h0)]);
                    end
                  for (forvar2131 = (1'h0); (forvar2131 < (1'h1)); forvar2131 = (forvar2131 + (1'h1)))
                    begin
                      reg2132 <= reg1472;
                    end
                end
              else
                begin
                  reg2120 <= (8'ha0);
                  for (forvar2121 = (1'h0); (forvar2121 < (1'h0)); forvar2121 = (forvar2121 + (1'h1)))
                    begin
                      reg2122 <= ($signed($signed(reg1427[(2'h2):(1'h0)])) ?
                          $unsigned($unsigned((reg2104 ?
                              (8'ha7) : reg2126))) : $signed($unsigned(((8'had) >>> reg1477))));
                    end
                end
              reg2133 <= (8'hb3);
              if (reg1498)
                begin
                  for (forvar2134 = (1'h0); (forvar2134 < (2'h3)); forvar2134 = (forvar2134 + (1'h1)))
                    begin
                      reg2135 <= forvar2056[(1'h1):(1'h0)];
                    end
                  if ({forvar2035})
                    begin
                      reg2136 <= (reg1503 ?
                          $signed($unsigned((wire2031 ^ forvar2087))) : (reg2135 ?
                              reg1440[(2'h3):(2'h2)] : {(&reg1490)}));
                      reg2137 <= ((~|reg1445[(1'h0):(1'h0)]) ?
                          ({(reg2043 ?
                                  reg2072 : reg2113)} || $unsigned((reg1492 ?
                              forvar2069 : reg1502))) : ((!$signed(reg2086)) >> ((reg1452 != reg2080) >= reg1491[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg2136 <= ($signed((reg2083[(1'h0):(1'h0)] ?
                          $signed(reg2057) : {reg2099})) && (^~(|(~reg2073))));
                      reg2137 <= reg1456;
                      reg2138 <= {$unsigned(reg2076[(4'h9):(3'h7)])};
                      reg2139 <= (((8'hb5) ?
                              reg1453[(3'h7):(1'h0)] : (^reg1434[(3'h7):(3'h5)])) ?
                          ({forvar2054[(1'h0):(1'h0)]} ?
                              {{forvar2040}} : (forvar2103 - (+reg2085))) : reg1533);
                    end
                end
              else
                begin
                  reg2134 <= ((^$signed((forvar2082 ?
                      forvar2033 : reg2063))) | (8'ha2));
                  reg2135 <= ((($unsigned(reg1436) ?
                      forvar2056[(2'h3):(2'h2)] : $unsigned(forvar2076)) >>> $signed({forvar2033})) ~^ $unsigned((&(reg2083 - (8'hb4)))));
                end
              for (forvar2140 = (1'h0); (forvar2140 < (2'h3)); forvar2140 = (forvar2140 + (1'h1)))
                begin
                  if (reg2058[(1'h1):(1'h1)])
                    begin
                      reg2141 <= reg1497[(2'h2):(1'h1)];
                      reg2142 <= ({(~^(^~forvar2091))} - $signed(forvar2069));
                    end
                  else
                    begin
                      reg2141 <= $unsigned($signed((!{forvar2069})));
                      reg2142 <= (($signed(reg1519[(1'h0):(1'h0)]) ?
                          reg2048 : (^~(8'ha6))) * reg2093);
                    end
                  if (reg2047)
                    begin
                      reg2143 <= {reg2090};
                    end
                  else
                    begin
                      reg2143 <= $signed(forvar2044);
                      reg2144 <= (+$signed(($signed(reg2045) >>> $unsigned((8'hb0)))));
                      reg2145 <= reg2080[(2'h2):(1'h1)];
                    end
                  reg2146 <= $unsigned((+$signed((reg1513 ?
                      (8'ha1) : reg1462))));
                  for (forvar2147 = (1'h0); (forvar2147 < (1'h1)); forvar2147 = (forvar2147 + (1'h1)))
                    begin
                      reg2148 <= (~((reg2126 ?
                              $signed(reg1512) : reg2078[(1'h0):(1'h0)]) ?
                          reg2077[(1'h1):(1'h1)] : forvar2090[(3'h7):(3'h4)]));
                      reg2149 <= $signed(reg1461[(3'h5):(1'h1)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar2118 = (1'h0); (forvar2118 < (2'h2)); forvar2118 = (forvar2118 + (1'h1)))
            begin
              for (forvar2119 = (1'h0); (forvar2119 < (1'h0)); forvar2119 = (forvar2119 + (1'h1)))
                begin
                  reg2120 <= forvar2039;
                  if ($signed({(~(|forvar2086))}))
                    begin
                      reg2121 <= $unsigned(({forvar2147} ?
                          $signed(reg1436[(3'h5):(2'h3)]) : reg1422));
                      reg2122 <= $unsigned($signed((reg1477[(2'h2):(1'h1)] ?
                          $unsigned(reg1494) : wire2031[(2'h2):(2'h2)])));
                      reg2123 <= ($signed($unsigned(reg1516)) ?
                          ((~^reg2058) != $unsigned(reg1472)) : {{(reg2120 ?
                                      reg1422 : reg2138)}});
                      reg2124 <= forvar2052;
                    end
                  else
                    begin
                      reg2121 <= (^~reg2049);
                      reg2122 <= reg2041;
                      reg2123 <= $unsigned(reg1475);
                      reg2124 <= (((~^(reg2057 ? (8'ha7) : forvar2121)) ?
                          (forvar2097[(3'h7):(2'h3)] ?
                              $unsigned(reg1422) : reg1535[(3'h5):(2'h2)]) : $unsigned(reg2111[(2'h3):(2'h2)])) - reg1492[(1'h1):(1'h1)]);
                    end
                  if (($unsigned(((reg2121 ? reg2143 : (8'hb5)) * forvar2051)) ?
                      reg2112[(1'h1):(1'h1)] : $unsigned(forvar2035)))
                    begin
                      reg2125 <= (reg2095 ^ reg1524[(3'h4):(3'h4)]);
                      reg2126 <= ((-$unsigned($unsigned(reg2081))) ^~ (reg2086[(1'h1):(1'h0)] <<< forvar2039));
                      reg2127 <= reg1462[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2125 <= reg1429;
                      reg2126 <= $signed(forvar2093);
                      reg2127 <= (reg1463[(3'h4):(2'h2)] ?
                          ($unsigned($signed(reg1486)) ?
                              (!(reg2068 ?
                                  reg1443 : reg2051)) : $unsigned(reg2127)) : ($unsigned((8'hb6)) ?
                              $signed({reg1463}) : $signed({forvar2085})));
                    end
                end
              reg2128 <= reg1514;
              if ($signed(reg1508))
                begin
                  if (reg1423)
                    begin
                      reg2129 <= (8'hb8);
                      reg2130 <= forvar2118;
                    end
                  else
                    begin
                      reg2129 <= reg1464;
                      reg2130 <= (8'hb8);
                      reg2131 <= (wire2027 ? reg2126 : $signed(reg2064));
                      reg2132 <= {(reg2081 ? reg2107 : (|$signed(reg2049)))};
                    end
                  if ($unsigned({reg1504[(3'h5):(3'h5)]}))
                    begin
                      reg2133 <= reg1530[(3'h4):(1'h0)];
                      reg2134 <= (reg2069[(4'hd):(3'h6)] ?
                          (($signed(reg2073) ?
                              {reg1522} : {forvar2086}) * $unsigned($signed(forvar2120))) : (^((forvar2101 != (8'hb2)) ?
                              {(8'ha7)} : (reg2078 != reg2104))));
                      reg2135 <= $signed((~&$unsigned($unsigned(wire2031))));
                      reg2136 <= (^$signed(($signed(reg2117) ?
                          reg2039[(2'h2):(2'h2)] : (8'hae))));
                    end
                  else
                    begin
                      reg2133 <= $unsigned(($signed({forvar2077}) > $unsigned({reg1462})));
                    end
                  for (forvar2137 = (1'h0); (forvar2137 < (2'h2)); forvar2137 = (forvar2137 + (1'h1)))
                    begin
                      reg2138 <= forvar2069[(2'h3):(1'h1)];
                    end
                end
              else
                begin
                  reg2129 <= (reg1509 + reg2036);
                end
              reg2139 <= $signed($signed($signed((8'hae))));
            end
          for (forvar2140 = (1'h0); (forvar2140 < (1'h0)); forvar2140 = (forvar2140 + (1'h1)))
            begin
              if (reg2067[(1'h1):(1'h0)])
                begin
                  for (forvar2141 = (1'h0); (forvar2141 < (2'h3)); forvar2141 = (forvar2141 + (1'h1)))
                    begin
                      reg2142 <= $signed($signed($unsigned((+reg2137))));
                    end
                  for (forvar2143 = (1'h0); (forvar2143 < (2'h2)); forvar2143 = (forvar2143 + (1'h1)))
                    begin
                      reg2144 <= (reg2099[(4'h9):(2'h3)] >> ((~|$signed(reg2103)) ?
                          reg1504[(1'h0):(1'h0)] : ($unsigned((8'hb8)) >>> (reg2074 ?
                              reg2045 : (8'hba)))));
                      reg2145 <= (forvar2052 ?
                          (&(((8'hb7) ?
                              (8'hb0) : reg1536) == $signed((8'h9f)))) : (((reg1535 ?
                                  reg1487 : forvar2085) ?
                              (|(8'hb6)) : (&reg2063)) <= ((reg1468 ?
                                  forvar2118 : (8'hb4)) ?
                              $signed(reg1501) : (reg1532 ?
                                  (8'ha0) : reg1433))));
                    end
                  reg2146 <= reg1512[(2'h2):(1'h1)];
                  for (forvar2147 = (1'h0); (forvar2147 < (2'h3)); forvar2147 = (forvar2147 + (1'h1)))
                    begin
                      reg2148 <= $unsigned(forvar2120);
                      reg2149 <= $signed(((~^(~reg1420)) ?
                          reg1457[(2'h2):(2'h2)] : $unsigned((~^forvar2141))));
                    end
                end
              else
                begin
                  for (forvar2141 = (1'h0); (forvar2141 < (1'h0)); forvar2141 = (forvar2141 + (1'h1)))
                    begin
                      reg2142 <= (~&reg1526);
                      reg2143 <= ($unsigned(reg1516[(3'h6):(2'h2)]) * $signed({(reg2033 != reg2039)}));
                      reg2144 <= reg2042;
                      reg2145 <= reg2134[(3'h6):(1'h0)];
                    end
                  reg2146 <= (8'h9e);
                  if (reg1480)
                    begin
                      reg2147 <= ((&reg1429) ?
                          {reg2059[(1'h1):(1'h1)]} : (8'hb3));
                      reg2148 <= ((|({(8'hb7)} ?
                          {(8'ha8)} : $signed(reg1468))) != $signed(reg1500));
                      reg2149 <= reg1494[(2'h2):(2'h2)];
                      reg2150 <= $unsigned(reg1477[(4'hd):(4'ha)]);
                    end
                  else
                    begin
                      reg2147 <= (($signed((+reg1425)) + $signed(reg2148[(1'h0):(1'h0)])) ?
                          ({((8'hb1) ? forvar2131 : reg1506)} ?
                              forvar2081 : reg1529) : $signed($unsigned(reg2080[(3'h4):(3'h4)])));
                      reg2148 <= ({(((8'h9e) < reg1535) ?
                                  (|(8'h9e)) : reg1533)} ?
                          {(~(~^forvar2034))} : $signed(forvar2131[(3'h5):(3'h4)]));
                      reg2149 <= $signed($signed(reg1452));
                      reg2150 <= reg2065;
                    end
                  reg2151 <= ({((+reg1455) ^~ {reg1530})} ?
                      ($signed(reg2089) && {$unsigned(reg1489)}) : reg2117);
                end
            end
          for (forvar2152 = (1'h0); (forvar2152 < (1'h0)); forvar2152 = (forvar2152 + (1'h1)))
            begin
              if ({reg2125[(3'h7):(3'h4)]})
                begin
                  reg2153 <= $signed((8'hba));
                  for (forvar2154 = (1'h0); (forvar2154 < (1'h0)); forvar2154 = (forvar2154 + (1'h1)))
                    begin
                      reg2155 <= $signed(reg1499[(4'h8):(2'h3)]);
                    end
                  if ((^~forvar2078))
                    begin
                      reg2156 <= reg2104;
                      reg2157 <= (forvar2137[(1'h0):(1'h0)] > reg1500);
                      reg2158 <= $signed((($unsigned(reg2074) ?
                              $unsigned(reg2075) : reg2151[(3'h5):(1'h0)]) ?
                          forvar2147[(2'h3):(1'h1)] : reg1507[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg2156 <= (reg2117[(3'h6):(1'h1)] ?
                          $signed($signed(((8'ha6) ?
                              reg1530 : reg2095))) : (reg1517[(2'h3):(1'h0)] + forvar2131));
                      reg2157 <= $unsigned(reg1495[(2'h3):(1'h0)]);
                      reg2158 <= {(~|$signed(forvar2081[(2'h2):(1'h0)]))};
                    end
                end
              else
                begin
                  reg2153 <= (|(((reg2099 == reg2138) ?
                          (reg2055 ? forvar2141 : forvar2044) : (^~reg2038)) ?
                      reg1504[(4'hc):(4'h8)] : $unsigned($signed(reg1499))));
                  if ($unsigned(reg2060))
                    begin
                      reg2154 <= (^reg1483[(3'h6):(2'h2)]);
                      reg2155 <= reg1484[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg2154 <= (^~(($signed(forvar2147) & (reg2112 ?
                          reg1495 : reg1493)) ^ ((^(8'ha2)) < (reg1424 || reg1485))));
                      reg2155 <= ((forvar2124 + forvar2093) < (-($unsigned((8'had)) ?
                          (reg2042 ~^ reg1463) : {reg1487})));
                    end
                  for (forvar2156 = (1'h0); (forvar2156 < (2'h2)); forvar2156 = (forvar2156 + (1'h1)))
                    begin
                      reg2157 <= (8'h9e);
                      reg2158 <= ((reg1504 ?
                          reg1525 : $unsigned(((8'hba) > reg1453))) ^ (reg2106 > $unsigned((reg2102 << reg1530))));
                      reg2159 <= (forvar2056 ?
                          ($signed(reg2100) > (~(reg1463 >> reg1539))) : reg2073);
                      reg2160 <= {((~&$unsigned(forvar2096)) * (|(~&(8'hb9))))};
                    end
                  for (forvar2161 = (1'h0); (forvar2161 < (2'h3)); forvar2161 = (forvar2161 + (1'h1)))
                    begin
                      reg2162 <= $unsigned((^~(-$signed((8'hb4)))));
                      reg2163 <= (~^reg2079);
                    end
                end
              if (reg2159)
                begin
                  reg2164 <= {(($unsigned(reg2105) <= ((8'ha3) ?
                          reg1436 : reg1417)) && ((~reg2059) + (8'hb5)))};
                end
              else
                begin
                  if (($signed((-$signed(reg1529))) ^ (8'hba)))
                    begin
                      reg2164 <= (($unsigned(((8'haf) ? (8'hb8) : forvar2039)) ?
                          reg1500 : reg1524[(3'h4):(1'h0)]) ^~ reg2068);
                    end
                  else
                    begin
                      reg2164 <= $signed(({(reg2095 ?
                              reg1443 : reg2064)} != (reg2093 ?
                          (|reg2131) : $unsigned(reg2144))));
                    end
                  reg2165 <= $unsigned((^~$unsigned(reg2061)));
                end
              for (forvar2166 = (1'h0); (forvar2166 < (1'h0)); forvar2166 = (forvar2166 + (1'h1)))
                begin
                  for (forvar2167 = (1'h0); (forvar2167 < (1'h1)); forvar2167 = (forvar2167 + (1'h1)))
                    begin
                      reg2168 <= $unsigned($unsigned((!reg2106[(3'h4):(3'h4)])));
                      reg2169 <= $unsigned(reg1460[(3'h5):(3'h4)]);
                      reg2170 <= $unsigned($unsigned($unsigned(reg2115[(2'h3):(2'h2)])));
                    end
                  for (forvar2171 = (1'h0); (forvar2171 < (1'h0)); forvar2171 = (forvar2171 + (1'h1)))
                    begin
                      reg2172 <= $unsigned($unsigned($unsigned((reg1532 ^~ reg1539))));
                    end
                end
              for (forvar2173 = (1'h0); (forvar2173 < (2'h3)); forvar2173 = (forvar2173 + (1'h1)))
                begin
                  for (forvar2174 = (1'h0); (forvar2174 < (1'h1)); forvar2174 = (forvar2174 + (1'h1)))
                    begin
                      reg2175 <= reg2061[(3'h5):(3'h4)];
                      reg2176 <= reg1525[(2'h2):(1'h1)];
                      reg2177 <= ((($unsigned(reg1435) ?
                              ((8'ha0) & wire1416) : reg1450) <= (reg2106[(1'h1):(1'h1)] ?
                              (-reg2070) : $signed(forvar2049))) ?
                          $unsigned(reg2110) : {$unsigned($signed(forvar2096))});
                    end
                end
            end
          if ($unsigned(reg1464))
            begin
              reg2178 <= {reg2086};
              if ((reg2056[(2'h2):(1'h1)] ?
                  (^~((|forvar2131) ? $signed((8'hae)) : reg1526)) : reg1522))
                begin
                  for (forvar2179 = (1'h0); (forvar2179 < (2'h2)); forvar2179 = (forvar2179 + (1'h1)))
                    begin
                      reg2180 <= ({reg2074[(2'h2):(2'h2)]} ?
                          $unsigned((+(forvar2034 & reg2115))) : $unsigned((reg1491[(1'h0):(1'h0)] ?
                              $unsigned(forvar2054) : ((8'h9d) ~^ (8'hab)))));
                      reg2181 <= reg2056[(1'h0):(1'h0)];
                      reg2182 <= (forvar2061 ?
                          reg1502 : $signed((+(reg2090 ? (8'hb8) : reg1499))));
                    end
                  for (forvar2183 = (1'h0); (forvar2183 < (1'h1)); forvar2183 = (forvar2183 + (1'h1)))
                    begin
                      reg2184 <= (~^((reg1481[(1'h1):(1'h1)] ?
                          (|reg2049) : reg1450[(2'h3):(1'h1)]) >>> ((~&reg2099) ?
                          $unsigned(reg1431) : $unsigned((8'hb8)))));
                      reg2185 <= ($unsigned(((forvar2167 ? reg2132 : reg2118) ?
                              (8'haf) : $signed(reg2062))) ?
                          (~^$unsigned({(8'ha7)})) : (($unsigned(reg1438) - (reg1524 ?
                              reg2156 : reg2143)) <= (^$unsigned(reg2143))));
                    end
                end
              else
                begin
                  reg2179 <= reg2076;
                  reg2180 <= (^~(~^reg1469[(3'h4):(3'h4)]));
                  if ($signed((forvar2081[(2'h2):(1'h0)] ?
                      reg1476[(1'h1):(1'h0)] : (|reg2146))))
                    begin
                      reg2181 <= $signed(reg2041[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2181 <= $signed($unsigned(((!reg1445) ?
                          (reg1539 << (8'hba)) : $signed(reg1458))));
                      reg2182 <= $signed((&(~&(reg2122 == forvar2114))));
                      reg2183 <= reg2129;
                    end
                  for (forvar2184 = (1'h0); (forvar2184 < (1'h0)); forvar2184 = (forvar2184 + (1'h1)))
                    begin
                      reg2185 <= {forvar2078};
                      reg2186 <= $signed(($unsigned(reg2048[(3'h7):(3'h4)]) ^ (reg1494[(4'he):(1'h0)] == reg2138[(4'h9):(4'h8)])));
                    end
                end
              if ($signed({reg2181[(4'h8):(3'h6)]}))
                begin
                  if ((reg2159[(2'h2):(2'h2)] ~^ (reg2095 ?
                      (^reg2107) : $signed({forvar2034}))))
                    begin
                      reg2187 <= (reg2143 - $unsigned({(&reg1457)}));
                      reg2188 <= (~|{((reg2112 && reg2143) <<< (^(8'ha7)))});
                    end
                  else
                    begin
                      reg2187 <= (&$signed((-$signed(reg1500))));
                      reg2188 <= (~^{$signed((reg1482 ?
                              forvar2171 : reg2120))});
                      reg2189 <= {$unsigned(($signed(reg1534) ?
                              $unsigned(reg2082) : $unsigned(reg2110)))};
                      reg2190 <= $unsigned((^~reg2102[(2'h2):(1'h0)]));
                    end
                end
              else
                begin
                  reg2187 <= $unsigned({$signed(reg2188[(4'ha):(3'h6)])});
                  if ((~&((reg2179[(2'h2):(2'h2)] != forvar2064) <<< (+{reg1457}))))
                    begin
                      reg2188 <= $unsigned($unsigned(({wire2030} ?
                          (reg2168 ?
                              reg1475 : (8'hb3)) : ((8'hb4) << reg1446))));
                      reg2189 <= (({forvar2174} ?
                              $signed(forvar2143[(3'h4):(1'h1)]) : ((|forvar2076) * reg2175[(1'h0):(1'h0)])) ?
                          reg2135[(3'h6):(2'h2)] : (reg1423 >> $unsigned((-(8'hb3)))));
                      reg2190 <= $signed(reg2107);
                    end
                  else
                    begin
                      reg2188 <= {(+$unsigned(reg2048))};
                      reg2189 <= forvar2077[(1'h1):(1'h1)];
                      reg2190 <= (({(reg2127 ?
                                  reg1473 : reg1491)} <<< $unsigned($unsigned(reg2060))) ?
                          (^(|reg2041[(2'h2):(1'h0)])) : reg2082[(1'h1):(1'h1)]);
                      reg2191 <= $unsigned({reg2164[(1'h0):(1'h0)]});
                    end
                  for (forvar2192 = (1'h0); (forvar2192 < (1'h1)); forvar2192 = (forvar2192 + (1'h1)))
                    begin
                      reg2193 <= (^~forvar2090[(3'h7):(3'h6)]);
                    end
                  reg2194 <= forvar2118[(1'h0):(1'h0)];
                end
            end
          else
            begin
              for (forvar2178 = (1'h0); (forvar2178 < (2'h2)); forvar2178 = (forvar2178 + (1'h1)))
                begin
                  if ((^reg1435[(1'h1):(1'h1)]))
                    begin
                      reg2179 <= (reg2100[(1'h1):(1'h1)] ?
                          reg2191[(4'h8):(3'h5)] : reg1483);
                      reg2180 <= (($signed(reg1473) ?
                          $signed((reg2059 << reg2149)) : (^~$unsigned(reg2107))) ^~ reg1427[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg2179 <= forvar2093;
                      reg2180 <= $signed((8'ha9));
                    end
                  for (forvar2181 = (1'h0); (forvar2181 < (1'h0)); forvar2181 = (forvar2181 + (1'h1)))
                    begin
                      reg2182 <= ((&reg2084[(1'h0):(1'h0)]) ?
                          $signed(reg1506[(4'ha):(3'h7)]) : $unsigned($unsigned({(8'hb7)})));
                      reg2183 <= $unsigned((^~($signed(forvar2039) >> reg2131)));
                      reg2184 <= ($signed({{reg2064}}) * $unsigned(forvar2032));
                    end
                  if ($signed($signed((~|{(8'ha1)}))))
                    begin
                      reg2185 <= $signed({reg2189});
                      reg2186 <= reg1521[(4'hd):(1'h0)];
                      reg2187 <= {forvar2124[(2'h2):(1'h1)]};
                      reg2188 <= ({reg1421[(2'h3):(2'h3)]} ?
                          reg1521[(3'h4):(1'h1)] : ((|(forvar2076 ?
                                  reg2138 : reg2070)) ?
                              {(-forvar2078)} : $unsigned(reg1508[(4'hc):(2'h3)])));
                    end
                  else
                    begin
                      reg2185 <= ($unsigned($signed($signed((8'hb6)))) != (8'hb9));
                      reg2186 <= (reg2050 ?
                          reg1531[(4'hd):(4'hb)] : (&(~(reg2100 >> forvar2167))));
                    end
                  for (forvar2189 = (1'h0); (forvar2189 < (2'h2)); forvar2189 = (forvar2189 + (1'h1)))
                    begin
                      reg2190 <= reg1483[(3'h6):(3'h6)];
                      reg2191 <= (+($signed($signed(reg1421)) || $signed(reg2094[(2'h3):(2'h2)])));
                    end
                end
            end
        end
      for (forvar2195 = (1'h0); (forvar2195 < (1'h0)); forvar2195 = (forvar2195 + (1'h1)))
        begin
          if ((|$signed(((reg1445 << reg2045) ~^ reg1498))))
            begin
              for (forvar2196 = (1'h0); (forvar2196 < (2'h3)); forvar2196 = (forvar2196 + (1'h1)))
                begin
                  reg2197 <= $signed((8'hba));
                  for (forvar2198 = (1'h0); (forvar2198 < (2'h3)); forvar2198 = (forvar2198 + (1'h1)))
                    begin
                      reg2199 <= reg2100[(2'h2):(2'h2)];
                      reg2200 <= reg2094[(4'hc):(2'h3)];
                      reg2201 <= $unsigned({reg2057});
                      reg2202 <= $signed((^~(~|(reg2042 ? reg1537 : reg1421))));
                    end
                end
              for (forvar2203 = (1'h0); (forvar2203 < (1'h1)); forvar2203 = (forvar2203 + (1'h1)))
                begin
                  reg2204 <= $unsigned(($signed({(8'haf)}) <<< ($signed(forvar2109) ?
                      reg1420[(1'h1):(1'h1)] : reg1467[(1'h1):(1'h0)])));
                  if (forvar2178)
                    begin
                      reg2205 <= $unsigned($unsigned((~reg2162)));
                      reg2206 <= {(forvar2077[(3'h6):(2'h3)] == reg2188)};
                      reg2207 <= (forvar2072 ?
                          $unsigned($signed($signed(reg1525))) : $signed((~(~^(8'hb4)))));
                      reg2208 <= (reg2082 ?
                          reg2148[(2'h2):(1'h1)] : (~reg2033[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg2205 <= (forvar2076[(1'h1):(1'h0)] ?
                          ($signed($unsigned(reg1444)) ?
                              (~forvar2096[(3'h4):(1'h1)]) : (8'ha6)) : reg2191[(3'h6):(3'h4)]);
                      reg2206 <= (~|$signed($signed($signed(forvar2081))));
                    end
                end
              for (forvar2209 = (1'h0); (forvar2209 < (2'h2)); forvar2209 = (forvar2209 + (1'h1)))
                begin
                  if ((&(!forvar2034[(4'hd):(1'h1)])))
                    begin
                      reg2210 <= ($unsigned(reg2070) < (-{(~|forvar2095)}));
                    end
                  else
                    begin
                      reg2210 <= (~|(8'h9e));
                      reg2211 <= {$unsigned($unsigned(reg1456[(3'h6):(3'h5)]))};
                      reg2212 <= reg2061;
                      reg2213 <= $unsigned(($unsigned((reg2126 ?
                              reg1442 : reg2061)) ?
                          ((reg2048 ^ reg1448) ?
                              ((8'hb8) ?
                                  reg1471 : reg1468) : forvar2101) : {$unsigned(forvar2203)}));
                    end
                  reg2214 <= $signed((^((-reg1483) ?
                      (!reg1447) : $signed(reg1534))));
                end
            end
          else
            begin
              if ($signed((forvar2183[(4'he):(3'h5)] == $signed(reg2095))))
                begin
                  reg2196 <= (($unsigned(reg2052) >= wire1416[(3'h4):(2'h2)]) ?
                      ({(reg2180 >>> reg2045)} ~^ (8'ha0)) : (-$unsigned($signed(reg2199))));
                  for (forvar2197 = (1'h0); (forvar2197 < (1'h0)); forvar2197 = (forvar2197 + (1'h1)))
                    begin
                      reg2198 <= reg1420[(4'h8):(3'h6)];
                    end
                  for (forvar2199 = (1'h0); (forvar2199 < (2'h2)); forvar2199 = (forvar2199 + (1'h1)))
                    begin
                      reg2200 <= $unsigned(reg2105);
                      reg2201 <= (({(~&(8'had))} ^ reg2212) ?
                          reg1440[(3'h5):(1'h1)] : (8'haa));
                      reg2202 <= $unsigned((reg2058[(2'h2):(2'h2)] || $signed(reg1521)));
                    end
                  if (reg1521[(2'h3):(1'h0)])
                    begin
                      reg2203 <= reg2055;
                      reg2204 <= forvar2171;
                      reg2205 <= (-(forvar2062[(2'h3):(1'h1)] ?
                          $signed($unsigned((8'hb7))) : ((!reg2072) + reg2083)));
                    end
                  else
                    begin
                      reg2203 <= reg2102;
                      reg2204 <= ((~^(!reg1428[(1'h0):(1'h0)])) ?
                          forvar2131 : reg2130);
                    end
                end
              else
                begin
                  if ((forvar2077[(2'h3):(2'h3)] ? reg2214 : forvar2036))
                    begin
                      reg2196 <= reg1460[(3'h7):(3'h5)];
                      reg2197 <= ((&($signed(forvar2093) ?
                              (~|reg1488) : $signed(reg2181))) ?
                          {$unsigned((~|reg1477))} : (!(reg1449[(1'h0):(1'h0)] ^~ (reg1436 >> reg1444))));
                    end
                  else
                    begin
                      reg2196 <= $unsigned((reg1498[(1'h1):(1'h0)] <= $signed(reg2199[(3'h5):(2'h2)])));
                      reg2197 <= reg2143[(4'h8):(3'h5)];
                      reg2198 <= ((~|{$unsigned(reg2156)}) + (-((reg1480 >= reg1498) ?
                          forvar2052[(4'h9):(2'h3)] : reg1490)));
                    end
                  for (forvar2199 = (1'h0); (forvar2199 < (1'h0)); forvar2199 = (forvar2199 + (1'h1)))
                    begin
                      reg2200 <= (($signed((-reg2212)) >>> ($unsigned(reg2214) > (reg2170 - reg1481))) <<< reg2130);
                    end
                  for (forvar2201 = (1'h0); (forvar2201 < (1'h1)); forvar2201 = (forvar2201 + (1'h1)))
                    begin
                      reg2202 <= (~|(forvar2184 ? (-reg2118) : forvar2203));
                      reg2203 <= forvar2049[(1'h0):(1'h0)];
                    end
                  for (forvar2204 = (1'h0); (forvar2204 < (1'h0)); forvar2204 = (forvar2204 + (1'h1)))
                    begin
                      reg2205 <= forvar2082;
                      reg2206 <= $unsigned(((~^{(8'h9c)}) ~^ reg2213[(2'h3):(2'h2)]));
                      reg2207 <= {(+($unsigned(reg2090) ?
                              (~&forvar2082) : {reg2075}))};
                      reg2208 <= {reg2053[(3'h7):(1'h1)]};
                    end
                end
              if ((($unsigned(reg2149[(2'h2):(1'h0)]) ?
                      $signed(reg1527[(4'h8):(4'h8)]) : {(reg2053 > forvar2061)}) ?
                  reg2137 : ($unsigned((-reg2052)) ?
                      $unsigned((reg2051 != (8'ha6))) : {reg2094[(4'he):(3'h7)]})))
                begin
                  for (forvar2209 = (1'h0); (forvar2209 < (1'h1)); forvar2209 = (forvar2209 + (1'h1)))
                    begin
                      reg2210 <= $unsigned(reg1447);
                      reg2211 <= (!$unsigned(reg2131[(3'h4):(1'h0)]));
                      reg2212 <= reg2127[(4'h9):(1'h0)];
                      reg2213 <= (reg1433[(3'h4):(3'h4)] <<< reg2038);
                    end
                  for (forvar2214 = (1'h0); (forvar2214 < (2'h2)); forvar2214 = (forvar2214 + (1'h1)))
                    begin
                      reg2215 <= {({$unsigned(reg1430)} ?
                              {reg2078} : $signed((~^reg2065)))};
                      reg2216 <= ((~($signed(reg2190) ?
                              $unsigned(reg2060) : $unsigned((8'ha7)))) ?
                          $signed($signed((reg1484 ?
                              reg1454 : reg2069))) : (reg2127 ?
                              ((reg1495 ? reg2054 : reg1508) ?
                                  $unsigned(reg1426) : $signed(reg1433)) : $unsigned($unsigned(wire2029))));
                    end
                  for (forvar2217 = (1'h0); (forvar2217 < (1'h1)); forvar2217 = (forvar2217 + (1'h1)))
                    begin
                      reg2218 <= $signed(reg2068);
                    end
                  if ((reg2072 ?
                      $unsigned((forvar2086[(4'h8):(2'h3)] ?
                          (reg1425 ?
                              forvar2124 : reg1438) : $unsigned(reg2194))) : (reg2088[(2'h2):(1'h1)] ?
                          $signed((reg1475 ? (8'had) : reg2164)) : reg1503)))
                    begin
                      reg2219 <= $signed(reg1526[(2'h3):(2'h3)]);
                      reg2220 <= $unsigned(reg1427[(1'h0):(1'h0)]);
                      reg2221 <= $unsigned(($unsigned($unsigned(reg2039)) == reg2155));
                    end
                  else
                    begin
                      reg2219 <= $unsigned(($unsigned((~|reg1464)) < $unsigned(reg2212)));
                      reg2220 <= $unsigned(forvar2072);
                      reg2221 <= (!(-(8'hb7)));
                      reg2222 <= reg2072;
                    end
                end
              else
                begin
                  if ($unsigned($unsigned((reg2194 == $signed(reg2147)))))
                    begin
                      reg2209 <= (-(!(~$signed(reg1447))));
                      reg2210 <= reg1429[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg2209 <= $signed($signed((!forvar2049[(2'h2):(1'h0)])));
                      reg2210 <= $unsigned((~^(-reg2049[(3'h7):(2'h2)])));
                      reg2211 <= (|(~(wire2029 + $signed(reg1508))));
                    end
                end
              reg2223 <= reg2219[(4'hb):(1'h0)];
              for (forvar2224 = (1'h0); (forvar2224 < (2'h3)); forvar2224 = (forvar2224 + (1'h1)))
                begin
                  if ($unsigned({{$signed(reg1452)}}))
                    begin
                      reg2225 <= (~&($unsigned((~reg1497)) ?
                          (reg1514 ?
                              reg2057[(4'hc):(1'h0)] : $unsigned(forvar2198)) : reg2178[(1'h0):(1'h0)]));
                      reg2226 <= ((-{{reg2135}}) ?
                          reg2047 : (wire2031 || reg1464[(1'h1):(1'h0)]));
                      reg2227 <= (^~(-((reg1539 ?
                          (8'h9d) : reg1513) == (8'hb2))));
                    end
                  else
                    begin
                      reg2225 <= $signed((&$signed((reg1456 & reg2075))));
                      reg2226 <= reg2132;
                      reg2227 <= (^~(({(8'hb2)} ?
                          forvar2034 : {(8'ha5)}) >> (reg1509[(2'h3):(1'h0)] ?
                          (~&reg2049) : ((8'hb6) ? forvar2201 : reg2136))));
                      reg2228 <= forvar2078[(1'h0):(1'h0)];
                    end
                  for (forvar2229 = (1'h0); (forvar2229 < (1'h0)); forvar2229 = (forvar2229 + (1'h1)))
                    begin
                      reg2230 <= forvar2152;
                      reg2231 <= (-$signed(reg1475[(2'h2):(1'h1)]));
                      reg2232 <= $signed(forvar2181[(1'h1):(1'h0)]);
                      reg2233 <= (reg1507[(2'h2):(1'h1)] ?
                          {((^reg1422) ?
                                  (8'h9e) : (|(8'hb5)))} : reg1418[(2'h3):(2'h3)]);
                    end
                  if (reg2105[(2'h3):(1'h0)])
                    begin
                      reg2234 <= {$unsigned($signed(reg2067))};
                      reg2235 <= $unsigned({{reg1471[(3'h4):(1'h1)]}});
                    end
                  else
                    begin
                      reg2234 <= $signed($signed($unsigned((~|reg1460))));
                    end
                end
            end
          for (forvar2236 = (1'h0); (forvar2236 < (2'h2)); forvar2236 = (forvar2236 + (1'h1)))
            begin
              for (forvar2237 = (1'h0); (forvar2237 < (2'h2)); forvar2237 = (forvar2237 + (1'h1)))
                begin
                  reg2238 <= ($unsigned((((8'hb4) && forvar2183) >>> {reg2078})) + (-(&$unsigned((8'h9c)))));
                  for (forvar2239 = (1'h0); (forvar2239 < (2'h2)); forvar2239 = (forvar2239 + (1'h1)))
                    begin
                      reg2240 <= reg2146;
                      reg2241 <= {forvar2201[(4'h8):(4'h8)]};
                      reg2242 <= (($signed((wire1413 ?
                              (8'h9d) : reg1536)) | {(reg1502 >>> reg2095)}) ?
                          {$unsigned((~|(8'ha0)))} : (~^forvar2141[(3'h4):(1'h0)]));
                    end
                end
            end
          for (forvar2243 = (1'h0); (forvar2243 < (1'h0)); forvar2243 = (forvar2243 + (1'h1)))
            begin
              if ((forvar2087 ?
                  ($unsigned(forvar2237[(1'h1):(1'h0)]) && (reg2062 >= $unsigned(reg2069))) : $signed($signed((forvar2096 - reg1495)))))
                begin
                  reg2244 <= (-reg2087);
                end
              else
                begin
                  reg2244 <= (-reg2121);
                end
              if (forvar2127)
                begin
                  for (forvar2245 = (1'h0); (forvar2245 < (2'h3)); forvar2245 = (forvar2245 + (1'h1)))
                    begin
                      reg2246 <= $unsigned(reg2068[(3'h4):(1'h0)]);
                      reg2247 <= $unsigned(((|$signed(reg1460)) * ($signed(reg1417) <<< (reg1473 > (8'hb8)))));
                      reg2248 <= forvar2183[(4'ha):(3'h7)];
                      reg2249 <= $signed((forvar2109 ?
                          forvar2192[(1'h0):(1'h0)] : (^(reg2115 < reg1532))));
                    end
                end
              else
                begin
                  reg2245 <= forvar2034[(4'hb):(3'h5)];
                  for (forvar2246 = (1'h0); (forvar2246 < (1'h1)); forvar2246 = (forvar2246 + (1'h1)))
                    begin
                      reg2247 <= reg2191;
                    end
                end
            end
        end
    end
  assign wire2250 = (^~reg2210[(2'h2):(1'h1)]);
  assign wire2251 = ({(|{(8'hb5)})} < $signed(($signed(reg2242) && $unsigned(reg1454))));
  assign wire2252 = ($signed((&$unsigned((8'h9c)))) ?
                        (~((reg1427 ?
                            reg2138 : reg1445) >= reg1531)) : reg2176);
  assign wire2253 = $unsigned($unsigned(wire2030));
  always
    @(posedge clk) begin
      reg2254 <= (&(|(^~{reg2094})));
      reg2255 <= {reg2242};
      if ((reg1428[(1'h0):(1'h0)] ?
          reg1498[(1'h0):(1'h0)] : $unsigned(reg2040)))
        begin
          if ({$signed(((reg2177 - reg1438) > $signed(reg2054)))})
            begin
              if ($unsigned((+$unsigned($signed((8'haf))))))
                begin
                  if (($unsigned($unsigned($signed(reg2215))) ?
                      (8'hab) : {(~|(reg2158 < (8'hab)))}))
                    begin
                      reg2256 <= $signed(($signed(((8'hb1) ?
                              reg1486 : reg2106)) ?
                          (&(reg1471 && reg2083)) : (~&$unsigned(reg2061))));
                      reg2257 <= $signed(reg2052);
                      reg2258 <= (8'ha6);
                      reg2259 <= reg1443[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2256 <= (&reg2249[(4'hd):(1'h1)]);
                    end
                  for (forvar2260 = (1'h0); (forvar2260 < (1'h1)); forvar2260 = (forvar2260 + (1'h1)))
                    begin
                      reg2261 <= $signed(reg1483[(2'h3):(1'h0)]);
                      reg2262 <= (~^$unsigned($unsigned((8'hb2))));
                    end
                  for (forvar2263 = (1'h0); (forvar2263 < (2'h3)); forvar2263 = (forvar2263 + (1'h1)))
                    begin
                      reg2264 <= ($unsigned(reg1472) ?
                          $signed($signed($unsigned(reg1436))) : $signed(reg1529[(5'h10):(4'h9)]));
                      reg2265 <= ((~^({reg2143} ?
                          $signed(reg2156) : (reg2139 - reg1519))) & (^(~^reg1458)));
                      reg2266 <= {reg1437[(4'hf):(4'h8)]};
                      reg2267 <= ((!reg1463) >= reg1469[(3'h5):(3'h4)]);
                    end
                end
              else
                begin
                  if ((^~(-$unsigned(reg2095[(3'h6):(3'h6)]))))
                    begin
                      reg2256 <= $signed($signed($unsigned($signed(wire2031))));
                      reg2257 <= ($signed($unsigned((reg2241 ?
                          reg2147 : reg2180))) >> $unsigned({$unsigned(reg2145)}));
                      reg2258 <= (^~reg2188[(1'h1):(1'h0)]);
                      reg2259 <= {{$unsigned((reg2168 ? wire1416 : reg1437))}};
                    end
                  else
                    begin
                      reg2256 <= (reg1446 | (-(~|(reg1468 ?
                          (8'hb4) : reg1519))));
                      reg2257 <= reg1504[(3'h7):(3'h7)];
                    end
                  if ({reg2058})
                    begin
                      reg2260 <= ({{(reg1501 | (8'had))}} | $signed($signed(reg2262[(4'hc):(2'h3)])));
                      reg2261 <= (|((reg2138[(1'h0):(1'h0)] <<< (reg2267 | reg2093)) + $unsigned((8'h9d))));
                      reg2262 <= ((((reg2199 != (8'ha1)) >> $signed(reg1446)) <<< $unsigned((~&reg2187))) ?
                          wire1414 : $unsigned(reg2194[(4'he):(3'h4)]));
                      reg2263 <= wire1414;
                    end
                  else
                    begin
                      reg2260 <= reg1513;
                      reg2261 <= {((reg1435 ?
                                  wire2027[(3'h5):(1'h1)] : $signed((8'hab))) ?
                              $unsigned((reg2067 & reg2201)) : $signed($signed(reg2075)))};
                    end
                  for (forvar2264 = (1'h0); (forvar2264 < (2'h3)); forvar2264 = (forvar2264 + (1'h1)))
                    begin
                      reg2265 <= reg2118[(4'h9):(2'h2)];
                    end
                  for (forvar2266 = (1'h0); (forvar2266 < (1'h0)); forvar2266 = (forvar2266 + (1'h1)))
                    begin
                      reg2267 <= reg1424;
                      reg2268 <= ((reg2245 | $unsigned((reg1423 - reg2100))) ?
                          $unsigned(((~|reg1475) ?
                              (+reg2139) : (^~(8'h9d)))) : $signed($signed(reg1447)));
                      reg2269 <= (8'hb1);
                    end
                end
              if ({{(^$unsigned((8'ha0)))}})
                begin
                  for (forvar2270 = (1'h0); (forvar2270 < (1'h1)); forvar2270 = (forvar2270 + (1'h1)))
                    begin
                      reg2271 <= (reg1511[(2'h2):(1'h1)] - (~|reg1484[(2'h3):(2'h3)]));
                    end
                  if (reg2231)
                    begin
                      reg2272 <= $signed(({(^~reg1493)} ? reg2049 : reg2260));
                      reg2273 <= {$unsigned((reg1526[(1'h0):(1'h0)] >= (&(8'ha9))))};
                      reg2274 <= $unsigned(($signed((reg1478 && reg2257)) ?
                          (((8'hb3) <<< reg2269) | $unsigned(reg2186)) : reg2131));
                      reg2275 <= (+$unsigned((reg2103[(3'h6):(1'h0)] != {(8'h9e)})));
                    end
                  else
                    begin
                      reg2272 <= (reg2219[(2'h3):(1'h1)] ?
                          (^{reg2107}) : ((~&{reg2201}) ?
                              reg1417[(1'h0):(1'h0)] : $unsigned($unsigned(reg2124))));
                    end
                  if ($unsigned($signed(({(8'hb6)} ?
                      $signed(reg2154) : (~&reg2155)))))
                    begin
                      reg2276 <= (!{reg1438[(4'h9):(3'h5)]});
                      reg2277 <= (reg1462 >= reg2154[(3'h4):(2'h3)]);
                      reg2278 <= reg2222;
                      reg2279 <= ($unsigned(($signed(reg2271) * (-(8'ha1)))) ?
                          $unsigned(reg2271[(2'h2):(2'h2)]) : (($unsigned((8'ha9)) ?
                              (reg2078 ?
                                  (8'h9d) : reg1524) : reg1539) >>> {reg2183[(2'h2):(1'h1)]}));
                    end
                  else
                    begin
                      reg2276 <= (~&$unsigned(((reg1534 != reg1449) * wire1416[(4'ha):(2'h3)])));
                      reg2277 <= ((&$unsigned((reg2194 | reg2210))) ?
                          {(^(reg1493 ?
                                  reg2235 : wire2027))} : ($signed(reg2131[(3'h5):(1'h0)]) > ($signed(reg2154) ?
                              {reg1497} : (^reg1496))));
                      reg2278 <= reg2158;
                    end
                  if (reg2183)
                    begin
                      reg2280 <= reg2145[(1'h0):(1'h0)];
                      reg2281 <= $unsigned(reg2116);
                      reg2282 <= ($signed(reg2036[(2'h2):(2'h2)]) * ((((8'hba) & reg2083) ?
                              $unsigned(reg2189) : reg2078[(1'h1):(1'h0)]) ?
                          $signed({reg1511}) : ((&reg2260) >= (reg2267 ?
                              (8'ha2) : reg2122))));
                      reg2283 <= ($unsigned(reg2189) ?
                          $unsigned($unsigned($unsigned(reg2102))) : ((reg2052[(4'hb):(2'h2)] - forvar2264) >> $unsigned(((8'haf) ?
                              reg1477 : reg2188))));
                    end
                  else
                    begin
                      reg2280 <= wire2027[(3'h6):(3'h4)];
                      reg2281 <= reg1469;
                    end
                end
              else
                begin
                  reg2270 <= (reg2137[(2'h2):(1'h0)] - (8'ha1));
                  for (forvar2271 = (1'h0); (forvar2271 < (1'h0)); forvar2271 = (forvar2271 + (1'h1)))
                    begin
                      reg2272 <= ((reg1419 * (|(reg2214 ?
                          (8'hb8) : reg2158))) ~^ (-{$signed(reg2142)}));
                      reg2273 <= reg2123;
                      reg2274 <= {$signed($unsigned(reg2191))};
                    end
                  for (forvar2275 = (1'h0); (forvar2275 < (2'h2)); forvar2275 = (forvar2275 + (1'h1)))
                    begin
                      reg2276 <= ((+{reg2249[(3'h7):(2'h2)]}) ?
                          $signed($unsigned(reg2221[(1'h0):(1'h0)])) : reg1446);
                    end
                  for (forvar2277 = (1'h0); (forvar2277 < (1'h0)); forvar2277 = (forvar2277 + (1'h1)))
                    begin
                      reg2278 <= $signed((-(-$signed(reg1462))));
                      reg2279 <= (^~((reg2052 ~^ (wire2250 ?
                              (8'h9d) : reg1501)) ?
                          reg1430 : reg1450));
                      reg2280 <= reg2149[(1'h0):(1'h0)];
                    end
                end
            end
          else
            begin
              if ($signed(reg1452))
                begin
                  reg2256 <= (~|$signed(((reg2107 >= (8'ha1)) >>> reg1517)));
                  if (($signed(({reg2064} - (reg2097 ?
                      reg1428 : (8'hae)))) == reg2200[(4'hb):(4'hb)]))
                    begin
                      reg2257 <= ($unsigned($unsigned(reg2205)) ?
                          $unsigned((|(reg2143 - reg2197))) : (($unsigned(reg2035) ?
                              (~&(8'hb5)) : (-reg1516)) << $signed((reg2245 >>> reg1425))));
                      reg2258 <= ((((~reg2235) ?
                          $signed(forvar2275) : (~reg1436)) << reg1496[(3'h6):(3'h4)]) << ($signed($signed(reg1533)) ?
                          (8'hba) : {reg2190[(3'h7):(3'h7)]}));
                    end
                  else
                    begin
                      reg2257 <= reg1455;
                      reg2258 <= reg2053[(3'h6):(3'h5)];
                    end
                  for (forvar2259 = (1'h0); (forvar2259 < (2'h2)); forvar2259 = (forvar2259 + (1'h1)))
                    begin
                      reg2260 <= reg2259;
                      reg2261 <= reg1442;
                      reg2262 <= reg1477;
                      reg2263 <= reg2183[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  reg2256 <= $unsigned($signed($signed($unsigned(reg2141))));
                  for (forvar2257 = (1'h0); (forvar2257 < (2'h3)); forvar2257 = (forvar2257 + (1'h1)))
                    begin
                      reg2258 <= ((($unsigned(reg2211) ?
                                  $signed(reg2157) : (reg2244 ?
                                      wire2027 : reg2279)) ?
                              ((reg1509 ? reg2124 : reg2248) ?
                                  (reg2102 <<< (8'ha3)) : $unsigned(reg1420)) : $unsigned((~&reg2059))) ?
                          $unsigned(reg2075) : {$unsigned($unsigned(reg2205))});
                      reg2259 <= (^~$signed($signed(reg1433[(2'h3):(1'h0)])));
                      reg2260 <= ((+((reg2104 ?
                              reg2069 : reg2123) <<< (reg1422 == (8'hb9)))) ?
                          $unsigned(reg2043) : $unsigned($unsigned((~^reg2100))));
                    end
                end
            end
        end
      else
        begin
          if ((~$unsigned(reg2273)))
            begin
              if ({reg2208[(3'h7):(3'h5)]})
                begin
                  for (forvar2256 = (1'h0); (forvar2256 < (2'h3)); forvar2256 = (forvar2256 + (1'h1)))
                    begin
                      reg2257 <= $signed(reg2258[(1'h1):(1'h0)]);
                      reg2258 <= (reg2215 ?
                          reg2056 : $signed($unsigned(reg1534[(1'h0):(1'h0)])));
                      reg2259 <= $unsigned($signed($unsigned(reg2172[(2'h3):(1'h1)])));
                      reg2260 <= ((^~((+(8'h9f)) | reg2206)) * ((~&(~reg2169)) >> reg2108[(1'h0):(1'h0)]));
                    end
                  if ({((+((8'ha9) >> reg1446)) ?
                          reg2033[(2'h3):(1'h0)] : $signed({reg2244}))})
                    begin
                      reg2261 <= {reg2278};
                    end
                  else
                    begin
                      reg2261 <= (~(reg2186[(1'h1):(1'h1)] & ((reg2227 && reg2168) ?
                          $signed(reg1539) : reg2143)));
                      reg2262 <= $unsigned(reg1493);
                      reg2263 <= {forvar2266};
                    end
                  reg2264 <= $signed(((+$unsigned(forvar2257)) ?
                      $signed((reg2210 != reg2106)) : (!$unsigned((8'hb9)))));
                  for (forvar2265 = (1'h0); (forvar2265 < (1'h1)); forvar2265 = (forvar2265 + (1'h1)))
                    begin
                      reg2266 <= (^~($signed((8'had)) ?
                          (reg1514 ^ (reg2097 >>> wire2253)) : reg2146[(4'h8):(4'h8)]));
                      reg2267 <= (-reg1520[(4'h8):(2'h2)]);
                      reg2268 <= (~&reg2085);
                      reg2269 <= reg1532;
                    end
                end
              else
                begin
                  if ($signed((~&reg2220[(3'h5):(1'h0)])))
                    begin
                      reg2256 <= $unsigned($signed($unsigned(reg2235)));
                    end
                  else
                    begin
                      reg2256 <= ((({reg1445} <= (~(8'hb6))) ?
                          $signed((8'ha4)) : (|((8'ha3) ?
                              reg1502 : reg2214))) <<< reg1465);
                    end
                  if (reg1451)
                    begin
                      reg2257 <= $unsigned($unsigned($signed(((8'hb5) >> reg1461))));
                    end
                  else
                    begin
                      reg2257 <= ((reg2170 ?
                          $unsigned((reg2037 * reg2271)) : $signed($unsigned(reg1509))) >> $signed($signed((+reg2231))));
                      reg2258 <= ($unsigned((~^(!reg2257))) * reg1420[(2'h2):(2'h2)]);
                      reg2259 <= (wire2029[(1'h0):(1'h0)] >>> reg1475[(1'h0):(1'h0)]);
                      reg2260 <= wire1415[(2'h2):(1'h1)];
                    end
                  for (forvar2261 = (1'h0); (forvar2261 < (2'h3)); forvar2261 = (forvar2261 + (1'h1)))
                    begin
                      reg2262 <= $unsigned($unsigned(reg1478));
                      reg2263 <= ((!$unsigned((!reg1490))) ~^ reg2072);
                    end
                end
              if ({{($signed(wire2030) ? reg1501[(4'h8):(2'h3)] : (-reg1492))}})
                begin
                  reg2270 <= reg1509;
                  for (forvar2271 = (1'h0); (forvar2271 < (1'h1)); forvar2271 = (forvar2271 + (1'h1)))
                    begin
                      reg2272 <= $signed((reg1485[(4'h9):(2'h2)] ?
                          ((reg1494 ? reg2213 : reg2228) ?
                              $signed(reg2276) : {(8'ha8)}) : wire1416[(1'h0):(1'h0)]));
                      reg2273 <= (reg2087[(3'h7):(1'h1)] && (($unsigned((8'ha3)) > (reg2141 ?
                              (8'hab) : reg1512)) ?
                          {reg2055[(2'h3):(1'h1)]} : reg2233[(1'h1):(1'h1)]));
                      reg2274 <= wire2250;
                    end
                end
              else
                begin
                  for (forvar2270 = (1'h0); (forvar2270 < (2'h3)); forvar2270 = (forvar2270 + (1'h1)))
                    begin
                      reg2271 <= wire1412;
                      reg2272 <= $unsigned(((^~forvar2265) ?
                          (reg2120 * (reg2083 == forvar2261)) : reg2083[(1'h1):(1'h0)]));
                    end
                  reg2273 <= reg2169;
                  for (forvar2274 = (1'h0); (forvar2274 < (1'h0)); forvar2274 = (forvar2274 + (1'h1)))
                    begin
                      reg2275 <= (^(($unsigned((8'h9f)) <= $unsigned(reg1512)) >= ((reg1452 >= reg1418) ?
                          reg2272 : (reg2045 ? reg1444 : reg1457))));
                      reg2276 <= $unsigned((reg2055 + $signed((reg1514 << reg2162))));
                      reg2277 <= (($signed((8'h9c)) ?
                          reg1444 : reg2121) <= reg2060);
                      reg2278 <= reg2199;
                    end
                  if (reg2272)
                    begin
                      reg2279 <= (~&$signed(reg2281[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg2279 <= (^~(^{(~reg1417)}));
                    end
                end
              for (forvar2280 = (1'h0); (forvar2280 < (1'h1)); forvar2280 = (forvar2280 + (1'h1)))
                begin
                  if ((+$unsigned({$unsigned(reg2070)})))
                    begin
                      reg2281 <= ($unsigned((~^{reg1459})) <<< (reg1489 ?
                          (!reg2121[(2'h2):(1'h0)]) : ($signed(reg2274) >> (reg2059 <<< reg1534))));
                    end
                  else
                    begin
                      reg2281 <= (8'ha5);
                    end
                  if (($signed((reg2212 && (~^reg1467))) ?
                      (~^reg1520[(3'h4):(2'h2)]) : {{reg2223[(2'h3):(1'h0)]}}))
                    begin
                      reg2282 <= {(((^reg2223) != $signed(reg2144)) ?
                              reg2260 : $signed({(8'hb5)}))};
                      reg2283 <= reg1465;
                    end
                  else
                    begin
                      reg2282 <= ({reg2226} >= $signed((reg2090 ?
                          reg1464[(1'h0):(1'h0)] : reg2218)));
                      reg2283 <= $signed(reg1465[(3'h4):(2'h3)]);
                    end
                end
            end
          else
            begin
              if ((reg1471[(4'h8):(2'h2)] < {$signed(reg2164)}))
                begin
                  for (forvar2256 = (1'h0); (forvar2256 < (2'h3)); forvar2256 = (forvar2256 + (1'h1)))
                    begin
                      reg2257 <= (reg1431 ?
                          (&($unsigned(reg2060) ?
                              (reg2278 - reg2148) : ((8'ha6) ?
                                  reg1539 : reg2125))) : reg2261);
                      reg2258 <= (~^($signed((^reg1503)) ?
                          $signed($unsigned((8'ha3))) : (^(+reg2099))));
                      reg2259 <= reg1448[(3'h5):(3'h5)];
                    end
                  if ($signed(reg2083[(3'h5):(3'h4)]))
                    begin
                      reg2260 <= ({(8'ha4)} ?
                          $signed($unsigned({reg2120})) : {(~{(8'h9d)})});
                    end
                  else
                    begin
                      reg2260 <= ($unsigned($signed((reg1442 < reg2084))) ?
                          (~($unsigned(reg1499) * (~|reg2124))) : (reg2139[(1'h1):(1'h0)] ?
                              $unsigned({reg2033}) : ((&(8'hae)) <= $signed(reg2162))));
                    end
                end
              else
                begin
                  for (forvar2256 = (1'h0); (forvar2256 < (2'h2)); forvar2256 = (forvar2256 + (1'h1)))
                    begin
                      reg2257 <= $signed(reg2134[(2'h3):(1'h0)]);
                      reg2258 <= ($unsigned(reg2279[(3'h5):(2'h2)]) ?
                          ((reg1495 ~^ reg2268[(4'he):(1'h0)]) * (reg2108[(3'h7):(3'h5)] * reg1500[(2'h2):(1'h0)])) : $unsigned(reg1453[(4'hc):(4'hc)]));
                      reg2259 <= wire2251[(2'h2):(2'h2)];
                      reg2260 <= ($signed(reg1467[(3'h5):(2'h2)]) ?
                          (8'ha6) : reg2063);
                    end
                end
              for (forvar2261 = (1'h0); (forvar2261 < (1'h1)); forvar2261 = (forvar2261 + (1'h1)))
                begin
                  reg2262 <= ((reg1420 && reg2225) - $signed({(reg2127 <= reg2184)}));
                  if ((reg2263 ?
                      reg1433 : (wire2253 ?
                          (((8'hb1) ? reg2246 : reg2280) ?
                              $signed(reg1454) : reg2277[(3'h6):(1'h0)]) : (8'hb5))))
                    begin
                      reg2263 <= (!reg2216[(4'he):(4'ha)]);
                      reg2264 <= $signed((8'ha1));
                      reg2265 <= $signed($unsigned({reg1534[(2'h2):(1'h0)]}));
                    end
                  else
                    begin
                      reg2263 <= reg2219;
                    end
                end
              reg2266 <= $signed($signed((&(~|(8'hb5)))));
            end
          for (forvar2284 = (1'h0); (forvar2284 < (2'h2)); forvar2284 = (forvar2284 + (1'h1)))
            begin
              if ((reg2095[(3'h7):(2'h3)] ?
                  $signed(reg1450) : {(reg2157[(1'h0):(1'h0)] ?
                          wire2030[(3'h5):(3'h4)] : ((8'ha5) == reg1422))}))
                begin
                  if ((reg2235[(2'h2):(2'h2)] + {$signed(reg1477[(3'h7):(1'h0)])}))
                    begin
                      reg2285 <= (^(^~((8'ha8) ?
                          (reg1513 ? wire1414 : reg1527) : $signed(reg1468))));
                      reg2286 <= reg2057;
                    end
                  else
                    begin
                      reg2285 <= (($signed(reg2112) >> $signed($unsigned((8'hb3)))) ?
                          $signed(($signed(reg2213) < $unsigned(reg1526))) : (~(+$unsigned((8'h9e)))));
                      reg2286 <= $unsigned((|reg2122));
                      reg2287 <= {reg1512};
                      reg2288 <= (($signed({reg1529}) ?
                              reg2130[(3'h4):(1'h1)] : (reg2157 + (~^reg1455))) ?
                          (~^{(~|reg2155)}) : {((reg2046 + reg2103) >>> (reg1502 != reg1525))});
                    end
                  reg2289 <= $signed(($signed(reg2083[(4'h9):(3'h6)]) ^~ (8'hac)));
                  if ($signed(reg2139[(4'hb):(4'hb)]))
                    begin
                      reg2290 <= {reg1492};
                    end
                  else
                    begin
                      reg2290 <= (~^({((8'ha6) ?
                              reg2136 : reg1432)} - $unsigned(reg2076[(1'h1):(1'h0)])));
                      reg2291 <= (reg2242 ?
                          reg2117[(2'h3):(2'h3)] : reg1513[(1'h1):(1'h0)]);
                      reg2292 <= reg2156[(4'h8):(1'h1)];
                      reg2293 <= ($signed(reg2278[(4'hd):(2'h2)]) ?
                          $signed(reg1476[(1'h0):(1'h0)]) : $unsigned(reg2068));
                    end
                  for (forvar2294 = (1'h0); (forvar2294 < (2'h2)); forvar2294 = (forvar2294 + (1'h1)))
                    begin
                      reg2295 <= $signed($unsigned(reg2280));
                      reg2296 <= (~|{(reg2295[(3'h7):(2'h3)] + (reg2182 < (8'hb2)))});
                      reg2297 <= $unsigned(reg2209);
                    end
                end
              else
                begin
                  reg2285 <= $signed(reg2165);
                end
              reg2298 <= reg2038;
              for (forvar2299 = (1'h0); (forvar2299 < (2'h3)); forvar2299 = (forvar2299 + (1'h1)))
                begin
                  for (forvar2300 = (1'h0); (forvar2300 < (1'h1)); forvar2300 = (forvar2300 + (1'h1)))
                    begin
                      reg2301 <= $signed(reg2205);
                      reg2302 <= (~|$signed((reg1498 ?
                          (8'ha9) : (reg2205 ? reg2112 : reg1468))));
                      reg2303 <= (^~reg1529[(3'h5):(2'h2)]);
                      reg2304 <= reg2085;
                    end
                  reg2305 <= (^$unsigned((reg2069[(2'h3):(2'h2)] ?
                      reg1480[(3'h5):(2'h3)] : (reg2172 - reg1468))));
                  if ((reg2115 + ($signed(reg2142) ^ ((~&reg2177) >> (8'hb8)))))
                    begin
                      reg2306 <= {{($signed((8'h9c)) && (reg2278 ?
                                  reg1516 : reg1500))}};
                      reg2307 <= reg2201;
                      reg2308 <= ((~^$unsigned(((8'h9f) ?
                          reg2246 : (8'hab)))) ^~ $signed({$unsigned(reg2072)}));
                    end
                  else
                    begin
                      reg2306 <= ($unsigned(reg2139) ~^ (((reg1497 >= reg2164) ?
                          (8'hab) : $signed(forvar2261)) || reg2093[(3'h5):(1'h0)]));
                    end
                end
            end
          reg2309 <= reg2214;
          for (forvar2310 = (1'h0); (forvar2310 < (1'h0)); forvar2310 = (forvar2310 + (1'h1)))
            begin
              if ({reg2186[(2'h3):(1'h1)]})
                begin
                  reg2311 <= reg2194[(4'he):(2'h2)];
                  for (forvar2312 = (1'h0); (forvar2312 < (2'h3)); forvar2312 = (forvar2312 + (1'h1)))
                    begin
                      reg2313 <= $unsigned(reg2061);
                    end
                end
              else
                begin
                  for (forvar2311 = (1'h0); (forvar2311 < (2'h3)); forvar2311 = (forvar2311 + (1'h1)))
                    begin
                      reg2312 <= reg2221;
                      reg2313 <= (^~$unsigned((8'hb4)));
                      reg2314 <= reg2190[(4'h8):(1'h1)];
                    end
                  if ((~(-forvar2312[(3'h4):(2'h3)])))
                    begin
                      reg2315 <= ($signed(reg1444) ?
                          (8'had) : $signed($unsigned(reg2042[(2'h3):(1'h0)])));
                      reg2316 <= reg2055;
                    end
                  else
                    begin
                      reg2315 <= {wire2251[(3'h5):(1'h0)]};
                      reg2316 <= (($unsigned((reg2281 ?
                          reg2303 : (8'h9e))) >> (!(8'hb3))) ~^ reg1481[(2'h2):(2'h2)]);
                    end
                  if ((|(~|reg2035[(4'h8):(4'h8)])))
                    begin
                      reg2317 <= (!((~&reg2110[(3'h5):(2'h3)]) ?
                          (reg2307[(2'h3):(1'h0)] >>> {reg2201}) : ((8'ha1) ?
                              {reg1464} : {(8'haf)})));
                      reg2318 <= reg2198[(3'h7):(3'h5)];
                    end
                  else
                    begin
                      reg2317 <= (|(+$unsigned({reg2187})));
                      reg2318 <= $signed(wire1412);
                    end
                  reg2319 <= reg1463;
                end
              reg2320 <= ((((~(8'hb7)) ?
                  reg1535[(4'h8):(3'h5)] : (reg1502 ?
                      reg1480 : reg1509)) + (reg1521 ?
                  ((8'ha0) ? reg1457 : reg2054) : (reg2233 ?
                      reg2317 : reg2168))) << (~|(+reg2308)));
              for (forvar2321 = (1'h0); (forvar2321 < (2'h2)); forvar2321 = (forvar2321 + (1'h1)))
                begin
                  if ((reg1450 << (reg2060 ?
                      $signed((reg1488 ?
                          reg2153 : reg2197)) : reg2063[(3'h4):(1'h1)])))
                    begin
                      reg2322 <= reg2065;
                      reg2323 <= $signed((^(reg2287 >= $unsigned(forvar2299))));
                      reg2324 <= reg2087[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg2322 <= (reg2297[(2'h2):(2'h2)] ?
                          {{reg1482}} : (-(^~(reg2197 ? reg2160 : (8'hab)))));
                      reg2323 <= reg2136;
                    end
                  if ((reg2142 ?
                      {reg1483[(3'h5):(3'h5)]} : forvar2256[(2'h2):(1'h0)]))
                    begin
                      reg2325 <= ($signed((reg2263 ? reg2297 : reg1536)) ?
                          ($signed(reg1434) == {$unsigned(reg2311)}) : $signed($unsigned(reg2255)));
                    end
                  else
                    begin
                      reg2325 <= reg1538[(3'h5):(1'h1)];
                      reg2326 <= (~|$signed(reg2156[(2'h2):(2'h2)]));
                    end
                  if (reg2130[(3'h6):(1'h0)])
                    begin
                      reg2327 <= ((~|((+reg1426) ?
                              $unsigned((8'hb5)) : reg2293)) ?
                          ($unsigned(forvar2311[(1'h0):(1'h0)]) ?
                              (~&reg2045[(1'h1):(1'h0)]) : ((reg2241 ?
                                  (8'had) : reg1458) << (reg2082 && reg2180))) : ($signed((reg1533 & reg1462)) ?
                              $unsigned({reg2172}) : (~&(reg2124 ?
                                  reg2196 : reg1461))));
                      reg2328 <= reg2153[(4'hf):(4'he)];
                      reg2329 <= reg1517[(4'hb):(1'h0)];
                      reg2330 <= $signed($unsigned({{(8'h9f)}}));
                    end
                  else
                    begin
                      reg2327 <= (((&(|reg1504)) ~^ $signed(reg2041[(1'h1):(1'h0)])) ?
                          $unsigned(reg1432[(3'h5):(1'h0)]) : reg1472);
                      reg2328 <= (reg2136 ?
                          (^~(+(reg1499 ? reg2216 : (8'ha8)))) : (8'hb5));
                    end
                end
            end
        end
    end
  assign wire2331 = (+(reg1505 ?
                        {$unsigned(reg2219)} : (reg1524 ~^ $unsigned(reg2186))));
  always
    @(posedge clk) begin
      if (($signed(reg1524) == reg2313))
        begin
          for (forvar2332 = (1'h0); (forvar2332 < (1'h1)); forvar2332 = (forvar2332 + (1'h1)))
            begin
              if (($unsigned((((8'hb1) >= reg1459) != ((8'ha3) > reg2142))) ?
                  reg1459 : (reg2309 ?
                      (reg2330 ? (reg2139 ^ (8'h9e)) : (^~reg1417)) : reg1503)))
                begin
                  if (({((reg2149 ? reg1434 : reg1529) * (reg1419 * (8'hb6)))} ?
                      reg1448 : (^~($signed(reg2262) << reg1465))))
                    begin
                      reg2333 <= ($signed($unsigned((8'ha2))) ?
                          reg2107[(2'h2):(1'h1)] : $unsigned(reg2228[(3'h4):(1'h0)]));
                    end
                  else
                    begin
                      reg2333 <= (reg2269 ?
                          $unsigned(($signed((8'hb3)) >= ((8'ha4) ^~ reg1457))) : $signed((8'ha3)));
                      reg2334 <= $signed(((~&{reg1480}) || $signed(reg2289)));
                      reg2335 <= {reg2150[(3'h5):(2'h3)]};
                      reg2336 <= $signed((((^(8'h9e)) ?
                          (+reg1461) : (reg2278 ?
                              (8'ha2) : (8'had))) != ($unsigned((8'ha6)) ?
                          {reg2055} : $signed(reg2169))));
                    end
                end
              else
                begin
                  for (forvar2333 = (1'h0); (forvar2333 < (2'h3)); forvar2333 = (forvar2333 + (1'h1)))
                    begin
                      reg2334 <= {reg2262};
                      reg2335 <= reg2082[(1'h1):(1'h0)];
                      reg2336 <= {reg2073};
                    end
                  for (forvar2337 = (1'h0); (forvar2337 < (1'h1)); forvar2337 = (forvar2337 + (1'h1)))
                    begin
                      reg2338 <= (-$unsigned($signed((-reg1524))));
                      reg2339 <= (&reg2200[(2'h2):(1'h1)]);
                    end
                end
              for (forvar2340 = (1'h0); (forvar2340 < (1'h1)); forvar2340 = (forvar2340 + (1'h1)))
                begin
                  for (forvar2341 = (1'h0); (forvar2341 < (1'h0)); forvar2341 = (forvar2341 + (1'h1)))
                    begin
                      reg2342 <= (^$unsigned((reg1516[(4'h8):(2'h2)] ?
                          {reg2200} : $unsigned(reg2259))));
                      reg2343 <= (~reg1454[(1'h1):(1'h1)]);
                      reg2344 <= (+({(reg2181 || reg2329)} ?
                          {reg2207} : reg1517));
                      reg2345 <= (-$signed({reg2290[(1'h0):(1'h0)]}));
                    end
                end
              if ((+(reg2274 ?
                  (~&$signed(reg2262)) : $signed(((8'haf) ?
                      reg2297 : reg2260)))))
                begin
                  reg2346 <= $unsigned($unsigned(forvar2332));
                  if ($unsigned((reg1421 < (~|(reg2139 & (8'hb3))))))
                    begin
                      reg2347 <= reg2176[(2'h3):(2'h2)];
                      reg2348 <= reg2172;
                      reg2349 <= (($signed((reg2206 ?
                          (8'hb9) : reg2317)) * reg2077[(2'h3):(1'h1)]) & (~^reg2094[(4'hd):(4'hc)]));
                    end
                  else
                    begin
                      reg2347 <= ((~$unsigned(reg2106[(3'h4):(2'h3)])) ?
                          ($unsigned(reg2268) ?
                              reg2037 : ((!wire2252) ?
                                  $signed(reg2227) : $signed(forvar2333))) : $signed($signed($signed(reg1481))));
                      reg2348 <= $signed($unsigned($signed({reg2264})));
                    end
                  if (reg1427)
                    begin
                      reg2350 <= $unsigned((((^~reg2214) ?
                              $signed(reg2290) : (reg2198 ?
                                  reg2270 : reg1460)) ?
                          $unsigned((reg2150 && reg2154)) : (((8'hae) ?
                                  reg2343 : reg2147) ?
                              (reg2329 & (8'haf)) : reg2150)));
                      reg2351 <= ({reg2323[(3'h4):(1'h0)]} >= {$unsigned(((8'ha9) >= (8'ha2)))});
                    end
                  else
                    begin
                      reg2350 <= (8'had);
                      reg2351 <= reg2063[(3'h5):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar2346 = (1'h0); (forvar2346 < (2'h3)); forvar2346 = (forvar2346 + (1'h1)))
                    begin
                      reg2347 <= (~&(~^reg2175));
                      reg2348 <= reg2157[(3'h5):(3'h5)];
                    end
                  for (forvar2349 = (1'h0); (forvar2349 < (2'h2)); forvar2349 = (forvar2349 + (1'h1)))
                    begin
                      reg2350 <= (~(($signed(reg1482) || {reg1488}) | reg2062));
                      reg2351 <= $signed($signed($unsigned((reg2170 ?
                          reg1495 : reg2246))));
                      reg2352 <= reg2097[(3'h4):(1'h0)];
                    end
                  reg2353 <= reg2199[(4'ha):(1'h0)];
                end
            end
          reg2354 <= $signed(reg2095);
          for (forvar2355 = (1'h0); (forvar2355 < (2'h2)); forvar2355 = (forvar2355 + (1'h1)))
            begin
              for (forvar2356 = (1'h0); (forvar2356 < (2'h2)); forvar2356 = (forvar2356 + (1'h1)))
                begin
                  if (reg1418)
                    begin
                      reg2357 <= reg2063[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg2357 <= (~$unsigned(($unsigned(reg2297) ?
                          {reg1489} : reg2105)));
                      reg2358 <= reg1501[(4'he):(3'h5)];
                      reg2359 <= $signed(({reg2297[(1'h1):(1'h0)]} ?
                          $signed($signed(reg2133)) : reg2215[(3'h4):(2'h3)]));
                      reg2360 <= reg2060;
                    end
                  for (forvar2361 = (1'h0); (forvar2361 < (1'h1)); forvar2361 = (forvar2361 + (1'h1)))
                    begin
                      reg2362 <= $signed($unsigned(reg2078[(1'h1):(1'h0)]));
                      reg2363 <= ($signed((|(reg1452 ?
                          reg2040 : reg2079))) ^ (|(^~(reg2048 ?
                          reg2176 : reg2245))));
                    end
                  for (forvar2364 = (1'h0); (forvar2364 < (2'h2)); forvar2364 = (forvar2364 + (1'h1)))
                    begin
                      reg2365 <= (reg2324 ?
                          (reg2357[(2'h3):(2'h3)] ?
                              reg2292[(4'he):(2'h3)] : (~^(reg2219 & reg2285))) : $unsigned($unsigned((|reg2318))));
                      reg2366 <= reg2363;
                      reg2367 <= (8'ha9);
                    end
                  if ((&reg1505))
                    begin
                      reg2368 <= reg1459;
                      reg2369 <= ($signed($unsigned((+reg2315))) ?
                          reg1433[(1'h0):(1'h0)] : $signed(($signed(reg1527) ?
                              (reg1517 ? reg1467 : reg1476) : (+(8'hb0)))));
                      reg2370 <= reg2086[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg2368 <= reg2342;
                      reg2369 <= ((~|((+(8'hb4)) ~^ reg2273[(4'ha):(2'h3)])) << $unsigned(reg2206[(3'h6):(2'h3)]));
                    end
                end
              if ($signed(reg1524[(3'h6):(3'h5)]))
                begin
                  if ($unsigned(reg1490[(3'h5):(3'h4)]))
                    begin
                      reg2371 <= {$signed((&$unsigned((8'hb4))))};
                      reg2372 <= ((({reg2051} << (reg1437 ?
                              reg2057 : reg1465)) ?
                          ($unsigned(reg2136) ?
                              {(8'ha2)} : reg1457) : (((8'haa) * reg2075) != reg2057[(1'h1):(1'h0)])) ~^ $signed($signed((^reg2199))));
                    end
                  else
                    begin
                      reg2371 <= (!$signed(reg2082));
                      reg2372 <= reg2157[(2'h2):(1'h0)];
                    end
                  for (forvar2373 = (1'h0); (forvar2373 < (2'h3)); forvar2373 = (forvar2373 + (1'h1)))
                    begin
                      reg2374 <= ((~^reg2159[(3'h6):(1'h1)]) << reg1472);
                      reg2375 <= (~$unsigned({(|reg1501)}));
                    end
                  if ({reg2036})
                    begin
                      reg2376 <= reg2198;
                      reg2377 <= ((reg2187 ? reg2219 : (|reg2113)) & reg2369);
                    end
                  else
                    begin
                      reg2376 <= $signed(reg1427[(1'h0):(1'h0)]);
                      reg2377 <= (reg2082 << {$signed($unsigned(reg2349))});
                      reg2378 <= (^($signed(reg2376) ?
                          (8'hb1) : $unsigned(reg2157)));
                    end
                end
              else
                begin
                  for (forvar2371 = (1'h0); (forvar2371 < (2'h3)); forvar2371 = (forvar2371 + (1'h1)))
                    begin
                      reg2372 <= reg1486;
                      reg2373 <= (~forvar2371);
                      reg2374 <= ((-reg1460) ?
                          $unsigned(reg2090) : (({(8'h9d)} ?
                              $signed(reg2070) : reg2064) >> ($signed(reg2311) ?
                              (8'ha2) : ((8'hb6) <= (8'hb8)))));
                    end
                  for (forvar2375 = (1'h0); (forvar2375 < (2'h2)); forvar2375 = (forvar2375 + (1'h1)))
                    begin
                      reg2376 <= (reg2131[(2'h2):(2'h2)] * {wire2251});
                      reg2377 <= $signed($signed(reg2241));
                      reg2378 <= (~^(+(+(|reg1457))));
                    end
                  reg2379 <= (($signed($signed(reg2266)) << reg2293) ?
                      reg2089[(2'h3):(1'h1)] : reg2262[(3'h6):(1'h0)]);
                  for (forvar2380 = (1'h0); (forvar2380 < (2'h3)); forvar2380 = (forvar2380 + (1'h1)))
                    begin
                      reg2381 <= (!reg2121);
                      reg2382 <= reg1443[(2'h2):(1'h1)];
                      reg2383 <= reg2378[(3'h5):(3'h4)];
                      reg2384 <= ((~|reg2354) && $signed({$signed(forvar2337)}));
                    end
                end
              for (forvar2385 = (1'h0); (forvar2385 < (2'h2)); forvar2385 = (forvar2385 + (1'h1)))
                begin
                  for (forvar2386 = (1'h0); (forvar2386 < (2'h3)); forvar2386 = (forvar2386 + (1'h1)))
                    begin
                      reg2387 <= $signed((reg1535 ^~ $signed(reg2106[(2'h2):(1'h0)])));
                      reg2388 <= (8'hae);
                      reg2389 <= $signed($unsigned(reg1453));
                    end
                  reg2390 <= ((8'ha7) ^ (({reg2099} ?
                          (reg1536 + reg1420) : $signed(reg2233)) ?
                      $signed(reg1447[(1'h0):(1'h0)]) : $signed(wire2031)));
                  if ({($signed((reg1446 >= reg2232)) ^~ reg2275[(3'h5):(1'h0)])})
                    begin
                      reg2391 <= reg1422[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2391 <= $signed($signed($unsigned(((8'hae) & reg2138))));
                      reg2392 <= reg2221;
                      reg2393 <= ({{(~&reg1479)}} - reg2257);
                    end
                  for (forvar2394 = (1'h0); (forvar2394 < (1'h0)); forvar2394 = (forvar2394 + (1'h1)))
                    begin
                      reg2395 <= (^reg2068);
                      reg2396 <= reg1469;
                    end
                end
            end
          if ($signed(reg2326))
            begin
              reg2397 <= reg2072[(1'h0):(1'h0)];
              for (forvar2398 = (1'h0); (forvar2398 < (1'h1)); forvar2398 = (forvar2398 + (1'h1)))
                begin
                  for (forvar2399 = (1'h0); (forvar2399 < (1'h1)); forvar2399 = (forvar2399 + (1'h1)))
                    begin
                      reg2400 <= (reg2142[(1'h0):(1'h0)] + ($unsigned((reg2384 * reg2191)) != (reg2182[(3'h5):(2'h3)] != {reg2170})));
                    end
                end
            end
          else
            begin
              reg2397 <= $unsigned(reg2228);
              for (forvar2398 = (1'h0); (forvar2398 < (1'h1)); forvar2398 = (forvar2398 + (1'h1)))
                begin
                  for (forvar2399 = (1'h0); (forvar2399 < (2'h3)); forvar2399 = (forvar2399 + (1'h1)))
                    begin
                      reg2400 <= (reg1513[(3'h6):(3'h5)] + reg2283);
                      reg2401 <= {(&(reg1460[(3'h4):(3'h4)] ?
                              {forvar2337} : reg1448))};
                    end
                  if (reg1469[(4'ha):(3'h4)])
                    begin
                      reg2402 <= {(8'ha0)};
                      reg2403 <= reg2347[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg2402 <= ($unsigned((reg1494[(1'h0):(1'h0)] || $unsigned(reg2163))) ?
                          reg2278[(1'h0):(1'h0)] : reg2263[(1'h0):(1'h0)]);
                    end
                  for (forvar2404 = (1'h0); (forvar2404 < (2'h2)); forvar2404 = (forvar2404 + (1'h1)))
                    begin
                      reg2405 <= ($unsigned(forvar2333[(2'h2):(2'h2)]) | $signed(($signed(reg2115) ?
                          {reg1511} : (reg2209 ? (8'hb8) : reg2391))));
                      reg2406 <= reg2244;
                    end
                end
              if ({(reg1443 ?
                      $unsigned((reg2038 <<< reg2070)) : ((reg1464 ?
                          reg1441 : reg2049) + reg2291))})
                begin
                  for (forvar2407 = (1'h0); (forvar2407 < (2'h3)); forvar2407 = (forvar2407 + (1'h1)))
                    begin
                      reg2408 <= {$unsigned((~|reg1422[(3'h5):(1'h1)]))};
                      reg2409 <= $signed($unsigned(((reg2375 + reg2375) ^ ((8'ha9) ?
                          reg1505 : reg1455))));
                    end
                  if ($signed(reg2401[(3'h5):(3'h4)]))
                    begin
                      reg2410 <= (((|$signed(reg2367)) ?
                          {reg2051} : reg2319) >= ($unsigned((~|reg2228)) ?
                          $unsigned(reg1534[(1'h1):(1'h1)]) : ($signed(reg2228) ?
                              (8'h9f) : $signed(reg2053))));
                    end
                  else
                    begin
                      reg2410 <= $signed(({reg2098} ? (^{reg2170}) : reg2147));
                      reg2411 <= (&reg2264);
                      reg2412 <= (+(8'hb9));
                    end
                end
              else
                begin
                  if ($unsigned(($signed((reg1500 ^ reg2221)) ?
                      ((reg2071 ^~ reg2131) ?
                          $unsigned(reg2308) : (~|reg2084)) : ((+forvar2386) ?
                          (~^reg1468) : reg2183))))
                    begin
                      reg2407 <= reg2244[(3'h5):(2'h2)];
                      reg2408 <= reg1498;
                      reg2409 <= $signed($unsigned({(^reg1514)}));
                      reg2410 <= reg1499[(3'h6):(3'h4)];
                    end
                  else
                    begin
                      reg2407 <= (8'ha0);
                      reg2408 <= (|($unsigned(reg2194[(4'ha):(4'h9)]) ?
                          $unsigned($unsigned(reg2067)) : ((8'ha5) >> $signed(reg2240))));
                    end
                  if (($unsigned((reg2302[(4'h8):(4'h8)] ?
                          (reg1526 ? reg1524 : (8'ha6)) : (reg1434 ?
                              reg1483 : reg2055))) ?
                      reg2209 : $signed(($signed((8'h9c)) && (reg2218 ?
                          (8'ha0) : reg1482)))))
                    begin
                      reg2411 <= ((reg2084[(1'h1):(1'h0)] ?
                              reg2342 : (~^reg1469[(3'h6):(2'h2)])) ?
                          (8'hb0) : $signed(($signed(reg2378) - (-reg2041))));
                      reg2412 <= ((!($unsigned((8'hb0)) ?
                          (|reg2350) : (reg2210 * (8'haf)))) + reg2408);
                      reg2413 <= reg2201;
                    end
                  else
                    begin
                      reg2411 <= {(8'ha6)};
                      reg2412 <= reg2366;
                      reg2413 <= (reg2097 > (reg2124 >> ((reg2258 >>> reg2040) << forvar2373)));
                      reg2414 <= reg2379[(1'h1):(1'h0)];
                    end
                  if (reg2360[(2'h2):(2'h2)])
                    begin
                      reg2415 <= (^~(^{(reg1506 ? reg1535 : reg1445)}));
                      reg2416 <= ($unsigned(reg1503[(1'h0):(1'h0)]) ?
                          reg2194[(4'ha):(4'h9)] : (!reg2177));
                      reg2417 <= ($unsigned(reg2329) != reg2155[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2415 <= $unsigned((reg2246[(1'h0):(1'h0)] ?
                          reg2357[(1'h0):(1'h0)] : $signed((reg2222 ?
                              reg2111 : reg2209))));
                      reg2416 <= reg2051;
                      reg2417 <= ((~^(|forvar2356[(2'h2):(1'h0)])) ?
                          {$signed((reg2241 ^~ reg2233))} : (($signed(reg1433) != reg1424[(2'h2):(1'h1)]) >= forvar2371[(1'h1):(1'h0)]));
                    end
                end
              for (forvar2418 = (1'h0); (forvar2418 < (2'h3)); forvar2418 = (forvar2418 + (1'h1)))
                begin
                  for (forvar2419 = (1'h0); (forvar2419 < (2'h3)); forvar2419 = (forvar2419 + (1'h1)))
                    begin
                      reg2420 <= ((^$unsigned($signed((8'hb4)))) ^ (~^reg2105[(3'h7):(1'h0)]));
                      reg2421 <= reg2141;
                    end
                  if ($unsigned(reg2103[(1'h0):(1'h0)]))
                    begin
                      reg2422 <= $signed((~|((~reg2377) ?
                          reg1419[(1'h0):(1'h0)] : {reg2080})));
                      reg2423 <= (8'hb1);
                    end
                  else
                    begin
                      reg2422 <= ((8'ha2) ? $signed(forvar2399) : reg1448);
                      reg2423 <= (~^($signed($signed(reg2168)) <<< $unsigned(reg1539)));
                      reg2424 <= (((reg2406 ?
                              (8'hba) : ((8'hae) ?
                                  wire2030 : (8'haa))) ~^ ((~&reg1467) ?
                              wire1415[(1'h0):(1'h0)] : reg1536)) ?
                          wire2252 : reg2232[(3'h6):(3'h6)]);
                      reg2425 <= (+{$signed($signed(reg1447))});
                    end
                  for (forvar2426 = (1'h0); (forvar2426 < (2'h2)); forvar2426 = (forvar2426 + (1'h1)))
                    begin
                      reg2427 <= $signed((forvar2419[(2'h2):(2'h2)] || $unsigned((reg1519 ?
                          (8'haf) : reg1501))));
                      reg2428 <= (~|reg2069);
                      reg2429 <= (~|(^~(^~(reg2402 ? reg2099 : reg1455))));
                    end
                  for (forvar2430 = (1'h0); (forvar2430 < (1'h0)); forvar2430 = (forvar2430 + (1'h1)))
                    begin
                      reg2431 <= (reg2308[(1'h0):(1'h0)] ?
                          reg2144 : ($signed((reg2388 & reg2103)) ?
                              ((~&reg2387) * reg1477[(4'hc):(1'h1)]) : ((^~reg2429) ?
                                  $unsigned(reg2262) : reg2081)));
                      reg2432 <= ((|reg1507) == (8'haf));
                    end
                end
            end
        end
      else
        begin
          for (forvar2332 = (1'h0); (forvar2332 < (1'h1)); forvar2332 = (forvar2332 + (1'h1)))
            begin
              for (forvar2333 = (1'h0); (forvar2333 < (1'h1)); forvar2333 = (forvar2333 + (1'h1)))
                begin
                  if ((((~^reg2143[(3'h4):(2'h3)]) ?
                      $signed(reg2351[(1'h1):(1'h0)]) : reg2107) | $unsigned($unsigned($unsigned(reg2170)))))
                    begin
                      reg2334 <= ($signed(reg2179) ?
                          $unsigned(reg2270) : reg2187[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg2334 <= (~|reg2333[(4'h9):(3'h6)]);
                      reg2335 <= reg1443;
                    end
                end
              if ($unsigned($signed(($signed(wire1412) > $signed(reg1462)))))
                begin
                  for (forvar2336 = (1'h0); (forvar2336 < (1'h1)); forvar2336 = (forvar2336 + (1'h1)))
                    begin
                      reg2337 <= ((~|((reg1537 >>> reg2190) ~^ $unsigned(reg2391))) >= reg2348[(4'h8):(3'h6)]);
                      reg2338 <= $unsigned(($signed((reg1505 ?
                              reg2374 : forvar2361)) ?
                          $unsigned(reg2106) : ({(8'hb6)} >>> reg2337[(1'h0):(1'h0)])));
                    end
                  for (forvar2339 = (1'h0); (forvar2339 < (2'h3)); forvar2339 = (forvar2339 + (1'h1)))
                    begin
                      reg2340 <= (reg2350 <= (|$unsigned((reg2349 ~^ (8'hab)))));
                    end
                  reg2341 <= reg1435;
                end
              else
                begin
                  if ($unsigned((8'ha8)))
                    begin
                      reg2336 <= reg2333;
                      reg2337 <= reg2074[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg2336 <= (($unsigned(forvar2398[(1'h1):(1'h1)]) ?
                          $unsigned(reg1484) : (-(+forvar2394))) >> $signed((~reg2046)));
                      reg2337 <= (^$signed(reg2055));
                      reg2338 <= {$unsigned($signed({reg1449}))};
                    end
                end
              if ((8'h9f))
                begin
                  if (reg2065)
                    begin
                      reg2342 <= $signed((~&($unsigned(reg2264) << (8'hb2))));
                    end
                  else
                    begin
                      reg2342 <= $unsigned((((8'ha5) & (reg2100 ?
                          (8'ha5) : reg2102)) ^~ (reg2402[(2'h3):(1'h1)] <<< (~|reg2058))));
                    end
                  reg2343 <= $signed(reg2154);
                  if (($signed($signed((^reg2134))) ?
                      $unsigned(reg2118[(2'h3):(1'h1)]) : reg2071))
                    begin
                      reg2344 <= {$unsigned(({forvar2364} >>> $signed((8'ha6))))};
                      reg2345 <= reg2184[(4'ha):(1'h0)];
                      reg2346 <= $signed({$signed(reg2122[(1'h1):(1'h1)])});
                    end
                  else
                    begin
                      reg2344 <= reg1473[(1'h1):(1'h1)];
                      reg2345 <= reg2207[(1'h0):(1'h0)];
                      reg2346 <= ($signed({reg2313}) == $signed((8'hac)));
                      reg2347 <= $signed(reg2168[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  reg2342 <= $signed((reg2304 < (+$signed(reg2381))));
                end
              reg2348 <= {reg2272};
            end
          if (reg2415[(2'h2):(2'h2)])
            begin
              if ($signed(reg2307))
                begin
                  for (forvar2349 = (1'h0); (forvar2349 < (2'h3)); forvar2349 = (forvar2349 + (1'h1)))
                    begin
                      reg2350 <= $signed(($unsigned((|(8'ha8))) == ((reg2428 >> reg1446) ?
                          reg2314 : $unsigned(reg2070))));
                      reg2351 <= $signed(reg2255);
                    end
                  reg2352 <= forvar2399[(4'hb):(3'h6)];
                  reg2353 <= ($unsigned((-$signed(reg1434))) ?
                      (8'hb5) : forvar2418);
                  if ({reg2198[(3'h4):(2'h2)]})
                    begin
                      reg2354 <= $signed(reg2189);
                    end
                  else
                    begin
                      reg2354 <= reg2371;
                      reg2355 <= $signed(reg2407[(1'h1):(1'h0)]);
                      reg2356 <= {(reg2035 > (~&{reg2379}))};
                      reg2357 <= reg1419[(2'h2):(1'h1)];
                    end
                end
              else
                begin
                  if ($signed((((reg2297 ?
                      reg1423 : reg1491) <= $unsigned(reg2153)) | reg1457)))
                    begin
                      reg2349 <= $unsigned(((-{reg2258}) <= $unsigned(reg1492)));
                      reg2350 <= $unsigned(($unsigned($unsigned(reg1526)) >>> forvar2373[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg2349 <= (-(+$signed(reg1535[(4'h9):(1'h0)])));
                      reg2350 <= ((8'hb6) ?
                          reg1434 : $signed(reg1496[(2'h3):(2'h3)]));
                      reg2351 <= ($signed((~^$unsigned(reg2336))) ?
                          $signed($unsigned((~&forvar2430))) : ($unsigned($signed((8'ha4))) + (((8'ha0) && reg1492) != $signed(reg1504))));
                    end
                  reg2352 <= $unsigned(reg2402);
                  if ((reg1503 ?
                      ((-$signed(reg1432)) <= $unsigned($signed(reg2160))) : ((|$signed(forvar2419)) ?
                          $signed((reg2335 && reg2312)) : ((|reg2033) * (^reg2346)))))
                    begin
                      reg2353 <= (reg2424[(3'h6):(2'h2)] | $unsigned((+(reg2100 | reg2424))));
                      reg2354 <= $unsigned((reg1481[(2'h2):(1'h0)] && (((8'hb2) ?
                              (8'ha0) : reg2093) ?
                          reg2346 : $signed(reg1501))));
                    end
                  else
                    begin
                      reg2353 <= (reg1483[(1'h1):(1'h1)] << reg1418);
                    end
                end
              if (reg2144[(3'h5):(3'h4)])
                begin
                  for (forvar2358 = (1'h0); (forvar2358 < (1'h0)); forvar2358 = (forvar2358 + (1'h1)))
                    begin
                      reg2359 <= (8'hba);
                      reg2360 <= reg1462[(1'h1):(1'h1)];
                      reg2361 <= {reg1498};
                    end
                  for (forvar2362 = (1'h0); (forvar2362 < (1'h0)); forvar2362 = (forvar2362 + (1'h1)))
                    begin
                      reg2363 <= (-$signed($signed(reg2209)));
                      reg2364 <= (8'h9e);
                      reg2365 <= ($signed($signed($unsigned(reg1488))) ?
                          $signed({$unsigned(reg2052)}) : $signed($signed((8'hb3))));
                      reg2366 <= reg1524[(3'h7):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar2358 = (1'h0); (forvar2358 < (2'h2)); forvar2358 = (forvar2358 + (1'h1)))
                    begin
                      reg2359 <= reg2375[(2'h2):(1'h0)];
                    end
                  for (forvar2360 = (1'h0); (forvar2360 < (1'h1)); forvar2360 = (forvar2360 + (1'h1)))
                    begin
                      reg2361 <= reg2423[(2'h3):(2'h3)];
                      reg2362 <= (reg2256 && (reg2421[(1'h1):(1'h0)] ?
                          ($unsigned(reg2306) ?
                              {reg2357} : $signed(reg2074)) : reg2102[(2'h2):(1'h0)]));
                      reg2363 <= ($unsigned($signed((reg1522 ?
                              reg2158 : reg2062))) ?
                          (|($unsigned(reg1417) ?
                              (wire2251 ?
                                  reg1456 : reg2067) : reg2306)) : $signed($unsigned(reg1431[(4'ha):(3'h5)])));
                      reg2364 <= (reg2421 ?
                          (($signed(wire2029) >>> (reg2149 ?
                              (8'hb7) : reg2323)) || (reg1440[(3'h6):(3'h6)] ?
                              $unsigned((8'haa)) : $signed(reg2156))) : (~^$unsigned($unsigned(reg2392))));
                    end
                  if ((((+(8'h9f)) ?
                          ($signed((8'h9f)) ?
                              (^~reg2215) : (reg1484 ?
                                  reg1534 : reg2222)) : (&((8'ha7) * reg2242))) ?
                      (+$signed($unsigned((8'ha1)))) : $signed($signed((reg2068 ?
                          reg2390 : reg2200)))))
                    begin
                      reg2365 <= $signed($signed(({reg2318} != (reg2288 ?
                          reg2407 : (8'hb1)))));
                      reg2366 <= reg1503;
                      reg2367 <= $signed((~(&{(8'had)})));
                    end
                  else
                    begin
                      reg2365 <= (~&$unsigned(reg2078[(2'h2):(1'h1)]));
                    end
                  for (forvar2368 = (1'h0); (forvar2368 < (1'h1)); forvar2368 = (forvar2368 + (1'h1)))
                    begin
                      reg2369 <= {reg2062};
                      reg2370 <= wire2251[(1'h1):(1'h1)];
                      reg2371 <= reg2287[(1'h0):(1'h0)];
                      reg2372 <= reg2361[(3'h7):(2'h3)];
                    end
                end
              if (reg2396)
                begin
                  for (forvar2373 = (1'h0); (forvar2373 < (1'h1)); forvar2373 = (forvar2373 + (1'h1)))
                    begin
                      reg2374 <= ({$signed(((8'ha5) * reg2172))} ?
                          ($unsigned((reg2085 > reg2354)) ?
                              reg2136[(2'h2):(2'h2)] : (|(|reg1417))) : (reg2366[(2'h3):(2'h3)] ?
                              $unsigned((8'had)) : ({reg1430} > (reg2305 != reg1506))));
                    end
                  for (forvar2375 = (1'h0); (forvar2375 < (2'h3)); forvar2375 = (forvar2375 + (1'h1)))
                    begin
                      reg2376 <= ($signed(reg1432) >>> (($unsigned(reg2392) ?
                          (^~(8'haf)) : reg1463[(2'h3):(1'h1)]) <<< reg1475[(2'h2):(1'h0)]));
                      reg2377 <= reg2154[(3'h7):(3'h7)];
                      reg2378 <= ((~&(((8'ha4) || reg2041) > $unsigned(reg2082))) ~^ $unsigned({(wire2252 * reg2185)}));
                    end
                end
              else
                begin
                  if ((($signed($signed((8'h9f))) ?
                          ((forvar2419 & (8'hb7)) || (^(8'hb5))) : reg2147[(1'h0):(1'h0)]) ?
                      reg2205[(4'ha):(4'h9)] : {((reg2107 & reg2285) >= $signed(reg2346))}))
                    begin
                      reg2373 <= $unsigned($signed(reg2035));
                      reg2374 <= (^~(|reg2342[(4'hb):(1'h0)]));
                      reg2375 <= (~|$unsigned(($unsigned(forvar2394) ?
                          (&reg2297) : (reg2201 ? reg2245 : reg1462))));
                    end
                  else
                    begin
                      reg2373 <= (-(~^((|reg2203) >>> (~|reg2053))));
                      reg2374 <= $signed(($signed(reg2392) ?
                          $unsigned($signed(reg2412)) : $signed((~^(8'had)))));
                    end
                  if ((^~(!reg1437[(4'hb):(3'h6)])))
                    begin
                      reg2376 <= (($unsigned($signed((8'hb4))) ?
                              reg2255[(3'h6):(3'h5)] : $signed(reg2278[(3'h6):(2'h2)])) ?
                          $unsigned((~|(^~forvar2426))) : $signed($signed($unsigned(reg2129))));
                      reg2377 <= {(reg2225[(3'h7):(3'h5)] ?
                              (((8'ha5) && reg1525) ?
                                  (reg2389 == (8'h9d)) : reg2080[(3'h4):(1'h1)]) : $signed($signed(reg2254)))};
                    end
                  else
                    begin
                      reg2376 <= {$signed($signed((reg2125 || reg1539)))};
                    end
                  for (forvar2378 = (1'h0); (forvar2378 < (1'h1)); forvar2378 = (forvar2378 + (1'h1)))
                    begin
                      reg2379 <= (~^reg1512[(3'h5):(1'h1)]);
                    end
                end
              if (reg2136[(3'h5):(2'h2)])
                begin
                  for (forvar2380 = (1'h0); (forvar2380 < (1'h0)); forvar2380 = (forvar2380 + (1'h1)))
                    begin
                      reg2381 <= reg2223;
                      reg2382 <= (((|reg2180) ?
                          ($signed(reg2158) ^ (reg2047 > (8'hae))) : (~$unsigned(reg2359))) | ((&(reg2052 ^ reg2094)) ?
                          (!$signed(forvar2430)) : (8'hb6)));
                      reg2383 <= reg2287;
                    end
                  for (forvar2384 = (1'h0); (forvar2384 < (2'h3)); forvar2384 = (forvar2384 + (1'h1)))
                    begin
                      reg2385 <= $unsigned({(reg2221[(1'h1):(1'h0)] & (~&reg1508))});
                      reg2386 <= reg2197;
                      reg2387 <= reg2258[(3'h4):(1'h1)];
                      reg2388 <= reg2292[(1'h1):(1'h0)];
                    end
                  reg2389 <= ($unsigned((~|(reg2356 || reg2172))) ?
                      reg2076 : $unsigned((|$unsigned(reg2054))));
                end
              else
                begin
                  for (forvar2380 = (1'h0); (forvar2380 < (2'h3)); forvar2380 = (forvar2380 + (1'h1)))
                    begin
                      reg2381 <= $signed((reg1475[(2'h3):(2'h2)] ^~ {$unsigned(reg2190)}));
                      reg2382 <= (($unsigned(reg1507[(3'h7):(1'h0)]) << reg1448[(3'h7):(3'h4)]) < $unsigned(reg2372[(3'h4):(2'h2)]));
                      reg2383 <= ((reg1485 ?
                          reg2051[(3'h6):(1'h0)] : (+(reg2396 ?
                              reg2271 : reg2138))) == ((|$signed(reg1449)) ?
                          $unsigned($unsigned(reg2216)) : (8'hb7)));
                      reg2384 <= reg2153;
                    end
                  for (forvar2385 = (1'h0); (forvar2385 < (1'h1)); forvar2385 = (forvar2385 + (1'h1)))
                    begin
                      reg2386 <= $unsigned(reg2144);
                    end
                  reg2387 <= $signed($signed((8'hb9)));
                end
            end
          else
            begin
              for (forvar2349 = (1'h0); (forvar2349 < (1'h1)); forvar2349 = (forvar2349 + (1'h1)))
                begin
                  for (forvar2350 = (1'h0); (forvar2350 < (2'h3)); forvar2350 = (forvar2350 + (1'h1)))
                    begin
                      reg2351 <= $unsigned($signed($signed(reg1481)));
                      reg2352 <= $unsigned(($unsigned(reg2308) <<< {(reg1471 ~^ reg2037)}));
                    end
                  reg2353 <= reg2281[(1'h1):(1'h1)];
                end
              reg2354 <= $unsigned(reg2169[(3'h4):(1'h0)]);
            end
          if ((reg2349[(3'h6):(1'h0)] ?
              $unsigned(reg2260[(1'h0):(1'h0)]) : $signed(((reg2351 & reg2359) ?
                  (reg2135 & (8'hac)) : {reg2337}))))
            begin
              for (forvar2390 = (1'h0); (forvar2390 < (1'h0)); forvar2390 = (forvar2390 + (1'h1)))
                begin
                  for (forvar2391 = (1'h0); (forvar2391 < (1'h1)); forvar2391 = (forvar2391 + (1'h1)))
                    begin
                      reg2392 <= (($signed((reg2223 ? reg2222 : reg2185)) ?
                              ({reg1437} && (!reg2335)) : (^reg2341[(2'h2):(1'h0)])) ?
                          reg2098[(2'h2):(2'h2)] : (!$signed((reg2278 ?
                              reg2320 : (8'hb0)))));
                      reg2393 <= (((+(reg2202 ? reg2368 : reg2087)) ?
                              $unsigned((reg1469 | reg2223)) : (^reg2377)) ?
                          $signed($signed(reg2356)) : reg2212[(4'hb):(2'h3)]);
                    end
                end
            end
          else
            begin
              for (forvar2390 = (1'h0); (forvar2390 < (2'h3)); forvar2390 = (forvar2390 + (1'h1)))
                begin
                  for (forvar2391 = (1'h0); (forvar2391 < (2'h2)); forvar2391 = (forvar2391 + (1'h1)))
                    begin
                      reg2392 <= (+reg1508[(4'hb):(2'h3)]);
                      reg2393 <= $unsigned(({(reg1485 ? reg1534 : reg2187)} ?
                          ((8'h9c) ?
                              reg1452 : $unsigned(reg2339)) : $signed(reg2241)));
                    end
                  for (forvar2394 = (1'h0); (forvar2394 < (1'h1)); forvar2394 = (forvar2394 + (1'h1)))
                    begin
                      reg2395 <= reg2046;
                      reg2396 <= reg2325;
                    end
                  if ({{$unsigned((reg2401 ? (8'hab) : reg2071))}})
                    begin
                      reg2397 <= (8'h9c);
                      reg2398 <= reg1440;
                      reg2399 <= reg1430;
                      reg2400 <= (8'ha4);
                    end
                  else
                    begin
                      reg2397 <= (8'hb7);
                      reg2398 <= $signed(reg2147[(1'h0):(1'h0)]);
                      reg2399 <= reg2254;
                    end
                end
            end
          for (forvar2401 = (1'h0); (forvar2401 < (1'h1)); forvar2401 = (forvar2401 + (1'h1)))
            begin
              if ((~&(((~reg2364) ? $unsigned((8'hab)) : (~^(8'ha9))) ?
                  ($signed(forvar2360) == $signed(reg2289)) : reg2163[(3'h6):(3'h4)])))
                begin
                  if ({reg2142[(1'h0):(1'h0)]})
                    begin
                      reg2402 <= $signed((~&$signed((~^reg2061))));
                      reg2403 <= (!(reg1487[(3'h7):(2'h2)] | ({(8'hba)} ?
                          $signed(reg2431) : reg2209)));
                      reg2404 <= (reg1418[(1'h1):(1'h0)] ?
                          $unsigned(reg2309) : (forvar2333 ?
                              ((8'ha1) ?
                                  (^~reg2228) : $unsigned(wire1414)) : reg2301));
                    end
                  else
                    begin
                      reg2402 <= $unsigned($unsigned(reg2147));
                      reg2403 <= (wire1416[(3'h6):(3'h5)] == $signed((reg2200 && (reg2363 >= reg2057))));
                      reg2404 <= {$unsigned(reg2352)};
                      reg2405 <= $unsigned(((8'ha0) ?
                          (((8'h9e) + reg1477) << reg2235) : ($signed((8'hb1)) ?
                              (reg1485 ?
                                  reg2298 : (8'hab)) : $signed(reg1485))));
                    end
                  if ($unsigned(((((8'ha1) ? reg2179 : reg1535) ?
                      reg2261[(3'h6):(2'h3)] : $signed(reg1482)) >= reg1524[(2'h2):(2'h2)])))
                    begin
                      reg2406 <= (+(((reg2328 ?
                              reg1456 : reg2172) > {reg1534}) ?
                          reg2148[(1'h1):(1'h1)] : ((reg2267 ?
                              reg2208 : reg2231) | reg1464)));
                      reg2407 <= (reg2255 ?
                          (reg2283[(2'h2):(2'h2)] ^ $signed(reg1437)) : reg2266[(4'ha):(3'h5)]);
                      reg2408 <= (~(~&($unsigned((8'h9e)) ^~ {reg2181})));
                    end
                  else
                    begin
                      reg2406 <= reg1420;
                      reg2407 <= $signed(({{reg1432}} > ((^reg2077) ?
                          {reg2326} : (reg2104 < (8'hb2)))));
                      reg2408 <= reg2218[(4'ha):(3'h7)];
                    end
                end
              else
                begin
                  reg2402 <= forvar2340[(3'h4):(2'h2)];
                  for (forvar2403 = (1'h0); (forvar2403 < (2'h2)); forvar2403 = (forvar2403 + (1'h1)))
                    begin
                      reg2404 <= (reg2076 <= ((reg2357 <= $unsigned(reg2357)) ?
                          (reg2334[(4'hf):(4'hc)] ?
                              reg2339[(1'h0):(1'h0)] : ((8'ha9) ?
                                  reg2093 : (8'hb3))) : (^~$unsigned(reg2344))));
                    end
                  reg2405 <= $unsigned((forvar2364[(1'h0):(1'h0)] ?
                      reg2305 : reg2338[(2'h3):(2'h2)]));
                end
              for (forvar2409 = (1'h0); (forvar2409 < (1'h1)); forvar2409 = (forvar2409 + (1'h1)))
                begin
                  for (forvar2410 = (1'h0); (forvar2410 < (1'h1)); forvar2410 = (forvar2410 + (1'h1)))
                    begin
                      reg2411 <= reg2387[(3'h5):(2'h3)];
                    end
                  if (((~|{$unsigned((8'hb7))}) ?
                      ((reg2190[(3'h4):(1'h0)] ?
                              reg2271[(3'h7):(1'h1)] : $signed(reg2355)) ?
                          (forvar2346[(1'h0):(1'h0)] && (-(8'hb8))) : reg2266[(4'h8):(2'h3)]) : reg1441[(2'h2):(1'h1)]))
                    begin
                      reg2412 <= (|(+$signed((wire1414 ^ reg1485))));
                    end
                  else
                    begin
                      reg2412 <= (($unsigned($unsigned((8'ha3))) ?
                          forvar2385[(3'h4):(3'h4)] : $unsigned((!reg2289))) && (^reg2248[(1'h0):(1'h0)]));
                      reg2413 <= $signed((~&((reg1536 ?
                          reg1469 : (8'ha3)) == {reg2182})));
                    end
                  for (forvar2414 = (1'h0); (forvar2414 < (2'h3)); forvar2414 = (forvar2414 + (1'h1)))
                    begin
                      reg2415 <= $unsigned(reg2105[(2'h3):(2'h2)]);
                      reg2416 <= reg2412;
                      reg2417 <= ($signed(((forvar2362 >= reg2163) ~^ $signed(reg2396))) ?
                          ($signed($unsigned(reg2345)) * $unsigned($signed(reg1515))) : (((reg2145 ?
                                  reg1467 : reg2136) * (^reg2277)) ?
                              reg2130[(4'hd):(4'hc)] : {((8'ha1) ?
                                      reg2124 : (8'hab))}));
                    end
                  reg2418 <= $signed({reg2126});
                end
            end
        end
      if (($unsigned($signed($unsigned(reg2235))) ?
          $signed((+(reg2384 || reg1489))) : ((8'hb8) ^~ (8'h9f))))
        begin
          reg2433 <= $unsigned(reg2208);
          for (forvar2434 = (1'h0); (forvar2434 < (2'h2)); forvar2434 = (forvar2434 + (1'h1)))
            begin
              for (forvar2435 = (1'h0); (forvar2435 < (1'h1)); forvar2435 = (forvar2435 + (1'h1)))
                begin
                  for (forvar2436 = (1'h0); (forvar2436 < (1'h0)); forvar2436 = (forvar2436 + (1'h1)))
                    begin
                      reg2437 <= $signed($unsigned(reg2326[(4'hb):(1'h1)]));
                      reg2438 <= reg1446;
                      reg2439 <= ((!{reg1426}) ?
                          forvar2409[(4'h9):(1'h1)] : $unsigned($unsigned(reg2068[(3'h4):(1'h1)])));
                      reg2440 <= ((~&($signed((8'hb5)) ?
                              (-reg2058) : (+reg2221))) ?
                          (reg1536[(2'h3):(1'h0)] <= reg1509) : (+$signed((reg2141 ?
                              (8'hba) : (8'ha2)))));
                    end
                  for (forvar2441 = (1'h0); (forvar2441 < (2'h2)); forvar2441 = (forvar2441 + (1'h1)))
                    begin
                      reg2442 <= ((((|reg1517) ?
                                  $signed(reg2298) : (forvar2350 ^~ reg2132)) ?
                              (8'had) : ((reg1477 >> forvar2349) ?
                                  reg2293[(1'h0):(1'h0)] : {reg1464})) ?
                          reg2200[(2'h2):(1'h1)] : (^(reg2364[(1'h0):(1'h0)] * (reg2182 >> reg2184))));
                    end
                  for (forvar2443 = (1'h0); (forvar2443 < (2'h3)); forvar2443 = (forvar2443 + (1'h1)))
                    begin
                      reg2444 <= (&(reg2352[(1'h1):(1'h1)] ?
                          $signed((reg2106 ^ wire1416)) : $unsigned($unsigned(reg2308))));
                      reg2445 <= (~|(!$signed((~|(8'hb2)))));
                      reg2446 <= ((^~wire2252[(4'hc):(1'h0)]) ?
                          reg2128 : $signed($signed({reg2442})));
                    end
                  if (($signed(reg2338[(2'h3):(1'h0)]) - reg2194[(2'h3):(2'h3)]))
                    begin
                      reg2447 <= ((+((!reg2326) <= (-reg2442))) * reg2368[(1'h0):(1'h0)]);
                      reg2448 <= ({(-(reg1472 ?
                              reg2135 : reg1471))} ^ reg2333[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg2447 <= (+(~$signed(reg2213)));
                      reg2448 <= ($unsigned({(~|reg1445)}) <<< ($unsigned((~&reg1478)) ?
                          reg2370 : (reg1472[(2'h2):(1'h0)] ^ (reg2116 * (8'ha0)))));
                      reg2449 <= forvar2386;
                      reg2450 <= $signed($unsigned({(forvar2410 ?
                              reg2271 : forvar2430)}));
                    end
                end
              reg2451 <= $unsigned((((reg2092 & reg1495) <= $signed(reg2274)) ~^ ($unsigned((8'h9c)) && $unsigned(reg2138))));
              for (forvar2452 = (1'h0); (forvar2452 < (2'h3)); forvar2452 = (forvar2452 + (1'h1)))
                begin
                  if ((($signed($unsigned(reg2094)) > reg2033[(4'hc):(3'h5)]) + reg2343))
                    begin
                      reg2453 <= reg1485;
                    end
                  else
                    begin
                      reg2453 <= (8'ha9);
                    end
                end
            end
          for (forvar2454 = (1'h0); (forvar2454 < (2'h3)); forvar2454 = (forvar2454 + (1'h1)))
            begin
              for (forvar2455 = (1'h0); (forvar2455 < (2'h2)); forvar2455 = (forvar2455 + (1'h1)))
                begin
                  for (forvar2456 = (1'h0); (forvar2456 < (1'h1)); forvar2456 = (forvar2456 + (1'h1)))
                    begin
                      reg2457 <= reg2303;
                      reg2458 <= reg2075[(1'h0):(1'h0)];
                      reg2459 <= {{(8'haa)}};
                      reg2460 <= reg2102;
                    end
                  for (forvar2461 = (1'h0); (forvar2461 < (1'h1)); forvar2461 = (forvar2461 + (1'h1)))
                    begin
                      reg2462 <= (!(reg2302 ?
                          ($unsigned(reg2231) ?
                              (reg1532 + reg2301) : (+reg2448)) : (^((8'haa) ^ (8'ha2)))));
                      reg2463 <= $signed((+reg1507[(4'ha):(1'h0)]));
                    end
                end
              if ((|$unsigned(($unsigned(reg2169) >> $unsigned(reg2222)))))
                begin
                  reg2464 <= {reg2135[(2'h3):(1'h0)]};
                  for (forvar2465 = (1'h0); (forvar2465 < (2'h2)); forvar2465 = (forvar2465 + (1'h1)))
                    begin
                      reg2466 <= (~|reg2127);
                      reg2467 <= reg1453[(2'h2):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar2464 = (1'h0); (forvar2464 < (2'h3)); forvar2464 = (forvar2464 + (1'h1)))
                    begin
                      reg2465 <= (8'haa);
                      reg2466 <= {(^~($unsigned(reg1526) ? (8'haa) : reg2199))};
                    end
                  if (reg2420[(3'h5):(2'h2)])
                    begin
                      reg2467 <= (reg2410[(2'h3):(1'h1)] ?
                          (reg2373 << $unsigned($unsigned(reg2457))) : $unsigned((((8'hb4) || forvar2426) ?
                              {reg2232} : (~|(8'hb5)))));
                      reg2468 <= reg2188[(2'h3):(2'h2)];
                      reg2469 <= (reg2378[(2'h3):(2'h3)] ?
                          reg1431 : reg2225[(2'h3):(1'h0)]);
                    end
                  else
                    begin
                      reg2467 <= $signed(forvar2455);
                      reg2468 <= (reg2347 ?
                          reg2180 : (reg1427 >= reg2041[(1'h1):(1'h1)]));
                      reg2469 <= ({(|{reg2319})} >= (~|{(8'had)}));
                      reg2470 <= reg1456[(3'h5):(3'h5)];
                    end
                  reg2471 <= $unsigned($signed(reg2046[(3'h7):(3'h4)]));
                end
              for (forvar2472 = (1'h0); (forvar2472 < (1'h1)); forvar2472 = (forvar2472 + (1'h1)))
                begin
                  reg2473 <= reg2198[(1'h1):(1'h1)];
                  for (forvar2474 = (1'h0); (forvar2474 < (1'h0)); forvar2474 = (forvar2474 + (1'h1)))
                    begin
                      reg2475 <= $signed($signed({(~|reg1532)}));
                    end
                  reg2476 <= (~$unsigned({$signed(reg2244)}));
                end
              if ((^~(reg2143 ?
                  (|reg2051[(1'h1):(1'h0)]) : $unsigned(reg2125[(3'h4):(1'h0)]))))
                begin
                  if ($signed((!(^((8'hb6) <<< (8'h9c))))))
                    begin
                      reg2477 <= $signed((reg2115[(2'h3):(1'h1)] ?
                          (^~$signed(reg1422)) : $unsigned($signed(reg1431))));
                    end
                  else
                    begin
                      reg2477 <= reg2038[(3'h5):(3'h5)];
                      reg2478 <= $signed(reg2345[(2'h2):(1'h1)]);
                      reg2479 <= $unsigned((reg2397 ?
                          $unsigned($signed(wire2030)) : $unsigned(reg2116[(3'h5):(3'h5)])));
                    end
                end
              else
                begin
                  for (forvar2477 = (1'h0); (forvar2477 < (1'h1)); forvar2477 = (forvar2477 + (1'h1)))
                    begin
                      reg2478 <= forvar2390[(4'h9):(3'h4)];
                      reg2479 <= ((~&reg2043) ? $signed(reg2320) : reg2106);
                    end
                  if ((reg2371 >>> $unsigned((^~reg2365))))
                    begin
                      reg2480 <= (($unsigned((^reg2466)) ?
                          forvar2384[(1'h0):(1'h0)] : ({reg2465} - (reg2246 + reg1536))) > $signed($signed($unsigned(reg2304))));
                      reg2481 <= ($signed(($unsigned(reg1526) <<< reg2105[(3'h5):(3'h4)])) ?
                          {{(&reg2355)}} : {(reg2368 ?
                                  ((8'ha7) << reg2147) : reg2086[(4'hc):(3'h4)])});
                      reg2482 <= $unsigned($unsigned(reg2100));
                      reg2483 <= (^reg2071);
                    end
                  else
                    begin
                      reg2480 <= forvar2441[(4'h9):(3'h6)];
                    end
                  for (forvar2484 = (1'h0); (forvar2484 < (2'h3)); forvar2484 = (forvar2484 + (1'h1)))
                    begin
                      reg2485 <= forvar2350;
                      reg2486 <= $signed({($unsigned(reg1493) ?
                              (reg2267 ^~ reg2305) : reg2473)});
                      reg2487 <= $signed(reg2147[(1'h0):(1'h0)]);
                    end
                end
            end
        end
      else
        begin
          reg2433 <= (^({$unsigned(reg2425)} * ($signed(reg2333) ~^ {(8'ha9)})));
          for (forvar2434 = (1'h0); (forvar2434 < (1'h1)); forvar2434 = (forvar2434 + (1'h1)))
            begin
              for (forvar2435 = (1'h0); (forvar2435 < (2'h2)); forvar2435 = (forvar2435 + (1'h1)))
                begin
                  for (forvar2436 = (1'h0); (forvar2436 < (1'h1)); forvar2436 = (forvar2436 + (1'h1)))
                    begin
                      reg2437 <= $signed(reg2129[(2'h3):(1'h1)]);
                      reg2438 <= (((^~(reg2429 ? (8'hb5) : (8'hb5))) ?
                              $unsigned((reg2235 >= reg2048)) : forvar2336[(3'h7):(3'h6)]) ?
                          (+$unsigned((reg2146 == reg2408))) : $signed(wire2031[(2'h2):(1'h0)]));
                    end
                  reg2439 <= $unsigned(($signed((wire2252 >> reg2324)) - reg2256));
                end
            end
        end
      for (forvar2488 = (1'h0); (forvar2488 < (2'h2)); forvar2488 = (forvar2488 + (1'h1)))
        begin
          for (forvar2489 = (1'h0); (forvar2489 < (2'h2)); forvar2489 = (forvar2489 + (1'h1)))
            begin
              for (forvar2490 = (1'h0); (forvar2490 < (2'h2)); forvar2490 = (forvar2490 + (1'h1)))
                begin
                  reg2491 <= (8'hb1);
                end
              for (forvar2492 = (1'h0); (forvar2492 < (1'h1)); forvar2492 = (forvar2492 + (1'h1)))
                begin
                  if ($unsigned($signed(((8'hb0) << $signed(reg2381)))))
                    begin
                      reg2493 <= (~^reg2433[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg2493 <= reg1491[(3'h4):(2'h3)];
                      reg2494 <= (($signed((reg1451 ?
                              reg2432 : (8'haa))) >> reg2247) ?
                          ($unsigned((&forvar2465)) > ((reg2364 ?
                              reg2345 : reg2145) ~^ $signed(reg2265))) : $signed(($unsigned(reg2206) & $unsigned(reg2052))));
                      reg2495 <= ({$signed($unsigned((8'hb8)))} ?
                          reg2314[(1'h1):(1'h0)] : $signed(reg1534));
                      reg2496 <= (reg2420[(2'h2):(1'h1)] >= ((8'haf) << $unsigned(((8'had) == (8'hb8)))));
                    end
                end
              for (forvar2497 = (1'h0); (forvar2497 < (1'h0)); forvar2497 = (forvar2497 + (1'h1)))
                begin
                  if (((({reg2232} ?
                          (~|reg2137) : ((8'ha2) ? forvar2394 : (8'hac))) ?
                      reg2480 : $signed($signed(reg2054))) <= reg2058))
                    begin
                      reg2498 <= $unsigned(reg2421[(1'h0):(1'h0)]);
                      reg2499 <= $signed((8'hb9));
                    end
                  else
                    begin
                      reg2498 <= ($signed((!(!reg1448))) ?
                          ((|$unsigned(reg2359)) ?
                              reg2278[(1'h0):(1'h0)] : $unsigned(reg2124)) : (reg2298[(3'h6):(3'h5)] ?
                              (~^(^reg1475)) : $signed((8'hb5))));
                      reg2499 <= (8'ha3);
                      reg2500 <= {reg2107[(1'h1):(1'h1)]};
                      reg2501 <= (^(reg1514 ?
                          reg1423[(1'h1):(1'h0)] : (-{reg2172})));
                    end
                end
            end
          if (((!reg1457[(1'h0):(1'h0)]) ?
              $unsigned($unsigned((+reg2039))) : reg2143))
            begin
              if ($unsigned(((^~(reg2131 >> reg2305)) ?
                  $signed(reg2369[(4'hd):(4'hb)]) : reg2216[(4'h8):(3'h7)])))
                begin
                  if ($unsigned(reg1440[(3'h5):(3'h4)]))
                    begin
                      reg2502 <= (~((reg2067 ?
                          reg1427 : (reg2341 ?
                              reg1451 : reg2467)) + ({reg2264} ?
                          (reg1499 != reg1423) : $signed(reg2056))));
                      reg2503 <= $signed(reg1454[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg2502 <= ({reg2417[(1'h0):(1'h0)]} >>> reg2198[(1'h0):(1'h0)]);
                      reg2503 <= reg2112;
                      reg2504 <= reg2501;
                      reg2505 <= (reg2401[(3'h6):(2'h3)] || (|$signed($signed(reg2368))));
                    end
                  if (reg2235)
                    begin
                      reg2506 <= $signed($signed($signed((~^forvar2414))));
                      reg2507 <= reg1477;
                    end
                  else
                    begin
                      reg2506 <= reg2068[(3'h5):(3'h4)];
                      reg2507 <= ({reg2060} <= $unsigned(($unsigned(reg2372) ?
                          $unsigned((8'hb5)) : reg2485[(1'h0):(1'h0)])));
                      reg2508 <= ($signed(($unsigned(reg2503) ^ (!reg2163))) ?
                          $unsigned(({reg2387} ^~ reg2425[(3'h7):(3'h6)])) : forvar2484);
                      reg2509 <= (wire2027[(2'h3):(2'h3)] ?
                          ($signed($signed(reg2097)) ?
                              reg1449[(1'h1):(1'h1)] : ((^(8'hb7)) || reg2201[(3'h7):(3'h4)])) : $unsigned($unsigned($signed(reg2464))));
                    end
                  if (reg2437[(4'hb):(3'h5)])
                    begin
                      reg2510 <= $signed($unsigned($unsigned((8'ha9))));
                      reg2511 <= (($signed($unsigned(reg2244)) >> (forvar2332[(4'hb):(3'h5)] & {reg2069})) != {{(reg2120 ?
                                  reg2442 : (8'hb6))}});
                      reg2512 <= reg2447[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2510 <= $unsigned((reg1531 > $unsigned((reg2276 > reg2147))));
                      reg2511 <= $unsigned(($unsigned((reg2106 ?
                          reg2504 : reg2376)) | $signed((reg1524 ?
                          reg2442 : reg2170))));
                      reg2512 <= (($unsigned($unsigned(reg2478)) ?
                              (^~reg2427[(2'h3):(1'h1)]) : $signed((!reg2183))) ?
                          (~reg2204[(1'h1):(1'h1)]) : (&reg2317[(1'h0):(1'h0)]));
                    end
                  for (forvar2513 = (1'h0); (forvar2513 < (1'h0)); forvar2513 = (forvar2513 + (1'h1)))
                    begin
                      reg2514 <= $unsigned((reg1471 ?
                          ($signed(reg2504) ?
                              (~reg2457) : (forvar2336 ?
                                  reg2427 : (8'hb8))) : {$signed(reg2365)}));
                      reg2515 <= (!(!reg2470[(4'ha):(4'h9)]));
                      reg2516 <= (~^(wire2253[(1'h1):(1'h1)] ?
                          (^~((8'hb9) ? reg1483 : reg2162)) : reg2306));
                      reg2517 <= reg2511;
                    end
                end
              else
                begin
                  reg2502 <= {$signed($signed($signed(reg1507)))};
                  if (reg2346[(3'h6):(1'h1)])
                    begin
                      reg2503 <= (~&(reg2339[(1'h1):(1'h0)] << reg1444));
                      reg2504 <= ($unsigned({reg2478[(1'h1):(1'h0)]}) ?
                          ($unsigned({(8'had)}) > reg2041[(2'h3):(2'h2)]) : {($unsigned(reg2287) ?
                                  (reg2401 ?
                                      reg2134 : forvar2356) : {reg1526})});
                    end
                  else
                    begin
                      reg2503 <= wire2027[(2'h2):(2'h2)];
                    end
                end
            end
          else
            begin
              for (forvar2502 = (1'h0); (forvar2502 < (1'h0)); forvar2502 = (forvar2502 + (1'h1)))
                begin
                  reg2503 <= $unsigned($unsigned((reg1501 ?
                      {reg2458} : (&reg2157))));
                  if ($signed($unsigned(((|reg2210) < (8'hba)))))
                    begin
                      reg2504 <= $unsigned(((~&{(8'h9c)}) << $unsigned(reg2255[(2'h3):(1'h1)])));
                    end
                  else
                    begin
                      reg2504 <= {reg2371[(1'h0):(1'h0)]};
                      reg2505 <= ($unsigned((8'hab)) ?
                          (($signed(reg2510) ?
                              {reg2469} : (^reg2080)) && $signed((8'hb2))) : (8'hb6));
                    end
                  for (forvar2506 = (1'h0); (forvar2506 < (2'h3)); forvar2506 = (forvar2506 + (1'h1)))
                    begin
                      reg2507 <= ((~^(8'h9c)) ?
                          $unsigned((reg2458 ?
                              $signed(reg1526) : (reg2225 ?
                                  reg2344 : (8'hb0)))) : $unsigned($signed(reg2095)));
                      reg2508 <= (reg2088 ?
                          (+($signed(forvar2513) ~^ $signed(reg2099))) : $signed($signed(reg1511)));
                      reg2509 <= reg1459[(1'h0):(1'h0)];
                      reg2510 <= $signed($signed((reg1458[(2'h3):(2'h2)] ?
                          reg2099 : forvar2401)));
                    end
                end
            end
        end
      for (forvar2518 = (1'h0); (forvar2518 < (2'h2)); forvar2518 = (forvar2518 + (1'h1)))
        begin
          for (forvar2519 = (1'h0); (forvar2519 < (2'h3)); forvar2519 = (forvar2519 + (1'h1)))
            begin
              if (($signed((~reg2468)) ?
                  ((forvar2464 ?
                      $signed(reg2403) : $signed(reg2125)) <= reg2325[(2'h2):(1'h0)]) : $unsigned({reg1491[(3'h4):(2'h2)]})))
                begin
                  for (forvar2520 = (1'h0); (forvar2520 < (2'h3)); forvar2520 = (forvar2520 + (1'h1)))
                    begin
                      reg2521 <= $unsigned(reg1425);
                      reg2522 <= {(({reg2142} && forvar2492) == ((reg2507 != reg2393) ?
                              (~reg2046) : (reg2398 ? reg2510 : reg2347)))};
                      reg2523 <= $unsigned((($signed(reg2427) < $signed(reg2420)) <<< ({forvar2391} ?
                          (~forvar2506) : (-(8'haf)))));
                      reg2524 <= {(($signed(reg2154) >= (-reg2315)) >>> (reg2086 ?
                              (reg2059 > reg2504) : (forvar2488 > (8'hb9))))};
                    end
                  if ($signed($signed($unsigned($signed(forvar2361)))))
                    begin
                      reg2525 <= reg2293;
                      reg2526 <= forvar2488;
                      reg2527 <= $unsigned(({$signed((8'ha1))} >= ((8'hb0) ?
                          reg1443 : $unsigned(forvar2358))));
                      reg2528 <= {{($signed(reg2370) == $unsigned(reg2103))}};
                    end
                  else
                    begin
                      reg2525 <= (reg2498 || $signed(((~^reg1509) < ((8'hb1) < reg2470))));
                    end
                  reg2529 <= $signed(((~|(reg2180 && reg2268)) ?
                      reg2257[(1'h0):(1'h0)] : {((8'hb3) ?
                              reg2485 : reg2133)}));
                end
              else
                begin
                  if ((|$unsigned(($unsigned(forvar2441) ^~ ((8'ha1) ?
                      reg2156 : (8'hba))))))
                    begin
                      reg2520 <= ($signed((&$unsigned(reg2296))) <<< (~|$unsigned($signed(reg2127))));
                      reg2521 <= $unsigned(reg1442[(4'h9):(2'h2)]);
                      reg2522 <= $unsigned(reg1517);
                      reg2523 <= ((reg2333 ? reg2411[(4'hc):(2'h2)] : (8'hb5)) ?
                          $unsigned($signed({reg1476})) : (((8'ha6) ?
                                  (reg2212 ^ reg2037) : $unsigned(forvar2362)) ?
                              $signed($signed(reg2207)) : $signed($unsigned(reg2387))));
                    end
                  else
                    begin
                      reg2520 <= $signed({reg2471});
                      reg2521 <= (^~{((+reg2428) << (reg2413 ~^ reg1418))});
                      reg2522 <= ($unsigned((reg2459[(3'h4):(3'h4)] ?
                          reg2529[(2'h3):(1'h1)] : (reg2406 ?
                              reg1433 : reg1445))) >= ($signed($signed((8'haf))) + (reg2505 ?
                          ((8'hb7) ?
                              reg2135 : reg2302) : (reg2293 || reg2033))));
                      reg2523 <= reg2289[(3'h5):(2'h2)];
                    end
                  reg2524 <= $unsigned((reg2439 ?
                      reg2081[(2'h3):(1'h0)] : ((reg2063 ? reg2041 : reg2514) ?
                          $signed(reg2512) : $signed((8'h9c)))));
                  for (forvar2525 = (1'h0); (forvar2525 < (2'h3)); forvar2525 = (forvar2525 + (1'h1)))
                    begin
                      reg2526 <= (|((reg2357[(2'h3):(1'h0)] <<< ((8'ha7) ?
                          reg2257 : (8'ha3))) == (^((8'ha4) ?
                          wire1414 : reg1461))));
                      reg2527 <= (($unsigned($signed(reg1508)) > reg2409) ?
                          reg2449 : $unsigned((reg1535[(4'ha):(4'ha)] ?
                              reg1492[(4'hd):(3'h4)] : $signed(reg2244))));
                    end
                end
              for (forvar2530 = (1'h0); (forvar2530 < (2'h2)); forvar2530 = (forvar2530 + (1'h1)))
                begin
                  if (($signed($unsigned((reg2125 >= reg2371))) ?
                      reg2368[(2'h3):(2'h2)] : reg2343))
                    begin
                      reg2531 <= $unsigned($unsigned((reg2045[(1'h1):(1'h0)] ^ $signed(reg1519))));
                      reg2532 <= $signed(($unsigned(reg2133) < $unsigned(((8'ha0) ?
                          reg1450 : forvar2398))));
                      reg2533 <= {((reg1475 ?
                              $signed(reg2289) : (^reg2050)) >>> $signed(reg2112))};
                      reg2534 <= {reg2142};
                    end
                  else
                    begin
                      reg2531 <= $unsigned($unsigned((+$unsigned(reg1461))));
                      reg2532 <= (!((8'ha7) ?
                          ($unsigned(reg2531) ?
                              $unsigned(reg2400) : (forvar2350 >> (8'ha4))) : reg2136[(4'h8):(4'h8)]));
                      reg2533 <= reg2069[(4'h9):(1'h1)];
                    end
                  for (forvar2535 = (1'h0); (forvar2535 < (2'h2)); forvar2535 = (forvar2535 + (1'h1)))
                    begin
                      reg2536 <= $signed(forvar2380);
                      reg2537 <= reg2375;
                      reg2538 <= ((forvar2362 ~^ $unsigned((reg2369 ?
                          reg2111 : reg2212))) >>> $signed((&$signed(reg2335))));
                    end
                end
            end
        end
    end
  assign wire2539 = reg2155[(4'ha):(2'h2)];
  always
    @(posedge clk) begin
      if (reg2397)
        begin
          for (forvar2540 = (1'h0); (forvar2540 < (2'h2)); forvar2540 = (forvar2540 + (1'h1)))
            begin
              reg2541 <= $unsigned((reg2453 ?
                  (^~$unsigned(reg2469)) : (^$unsigned(reg2118))));
              for (forvar2542 = (1'h0); (forvar2542 < (2'h2)); forvar2542 = (forvar2542 + (1'h1)))
                begin
                  for (forvar2543 = (1'h0); (forvar2543 < (2'h3)); forvar2543 = (forvar2543 + (1'h1)))
                    begin
                      reg2544 <= (^~((reg2345 != $signed(reg2462)) ?
                          {(reg1494 ~^ wire1415)} : $signed($signed(reg2351))));
                    end
                  for (forvar2545 = (1'h0); (forvar2545 < (2'h2)); forvar2545 = (forvar2545 + (1'h1)))
                    begin
                      reg2546 <= $signed($signed(((reg2451 != reg2223) != {reg2170})));
                      reg2547 <= (~|(^($unsigned(reg2363) ?
                          (8'hac) : $signed(reg1435))));
                      reg2548 <= $unsigned(reg2302);
                      reg2549 <= $unsigned((~|$unsigned($unsigned(reg2349))));
                    end
                  for (forvar2550 = (1'h0); (forvar2550 < (1'h0)); forvar2550 = (forvar2550 + (1'h1)))
                    begin
                      reg2551 <= $unsigned((^~$unsigned(reg2515[(2'h2):(1'h1)])));
                    end
                  if (wire2251[(3'h6):(2'h3)])
                    begin
                      reg2552 <= (&(~(reg2163 ?
                          (reg2054 ? reg2306 : reg2129) : $unsigned(reg2082))));
                      reg2553 <= (^((8'ha2) ?
                          {$signed(reg1417)} : ($signed(reg2226) >= reg2234)));
                    end
                  else
                    begin
                      reg2552 <= (!(!((reg2344 ?
                          reg2233 : reg2245) >>> {reg1468})));
                      reg2553 <= reg2115;
                      reg2554 <= reg2086;
                      reg2555 <= {reg2266[(2'h2):(2'h2)]};
                    end
                end
              for (forvar2556 = (1'h0); (forvar2556 < (2'h3)); forvar2556 = (forvar2556 + (1'h1)))
                begin
                  reg2557 <= {(((reg1450 * reg2491) ~^ $unsigned(reg1459)) ?
                          $signed(reg2511[(4'hf):(4'hc)]) : reg2362)};
                  reg2558 <= {$signed(($signed(reg2416) && reg2135[(3'h4):(1'h1)]))};
                  for (forvar2559 = (1'h0); (forvar2559 < (1'h1)); forvar2559 = (forvar2559 + (1'h1)))
                    begin
                      reg2560 <= $unsigned((((8'ha1) > reg2142[(2'h2):(1'h1)]) ?
                          (-{reg2320}) : (!reg2269[(1'h0):(1'h0)])));
                      reg2561 <= (reg2122 + reg1509[(3'h5):(1'h1)]);
                      reg2562 <= (8'hac);
                      reg2563 <= $unsigned($unsigned($signed($signed(reg2130))));
                    end
                end
            end
          if (((8'ha1) >> reg2261))
            begin
              if (reg1517)
                begin
                  if ($unsigned({((reg2558 | forvar2559) ?
                          (^reg2282) : $signed(reg2041))}))
                    begin
                      reg2564 <= (~|{{$signed(reg1499)}});
                      reg2565 <= reg2414;
                      reg2566 <= (reg2343 ?
                          (({(8'hb4)} < (reg2121 ?
                              reg1507 : reg2278)) + (|(reg2231 < reg2110))) : ({(~&reg2307)} ?
                              $unsigned((reg1530 >> reg1420)) : $unsigned((reg2288 != reg2385))));
                      reg2567 <= {reg2388[(3'h4):(3'h4)]};
                    end
                  else
                    begin
                      reg2564 <= (~^{reg1436});
                      reg2565 <= reg2437;
                      reg2566 <= (({reg2120} ?
                          ($unsigned(reg2407) ~^ (reg2493 ?
                              reg2177 : reg2416)) : {(~&reg2341)}) >= (8'hb0));
                    end
                  if ((&reg2445[(4'h8):(3'h5)]))
                    begin
                      reg2568 <= (reg2072[(2'h3):(1'h0)] != ({$unsigned(reg2411)} ?
                          reg2464[(3'h6):(2'h2)] : reg2275[(3'h5):(3'h5)]));
                      reg2569 <= reg2227[(4'h8):(3'h4)];
                      reg2570 <= $signed($signed(((^(8'h9e)) >= {reg1444})));
                      reg2571 <= (reg2429[(4'hb):(1'h1)] != ($unsigned($signed(reg2330)) ?
                          $signed((8'haa)) : reg1531));
                    end
                  else
                    begin
                      reg2568 <= (reg2135 || reg2105);
                      reg2569 <= (8'hae);
                      reg2570 <= reg2335;
                      reg2571 <= $signed((~(|reg2086[(4'hc):(1'h1)])));
                    end
                  if ((~$signed((~|wire2030))))
                    begin
                      reg2572 <= ($unsigned($signed((reg1508 ?
                          reg1530 : reg2413))) <<< (((reg2408 ?
                              reg2190 : (8'hb0)) ?
                          $signed(reg2438) : reg1442[(3'h7):(3'h5)]) && reg2279));
                      reg2573 <= reg2226;
                      reg2574 <= wire1412;
                      reg2575 <= (|reg2459);
                    end
                  else
                    begin
                      reg2572 <= reg1539;
                      reg2573 <= $signed(reg2134[(1'h1):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar2564 = (1'h0); (forvar2564 < (1'h1)); forvar2564 = (forvar2564 + (1'h1)))
                    begin
                      reg2565 <= ((~|reg2330[(3'h6):(3'h4)]) ?
                          ($signed(reg1431) | $signed((&reg2368))) : (($signed(reg1532) ?
                                  $unsigned(reg2325) : (~reg1508)) ?
                              (reg2142[(2'h3):(2'h2)] ?
                                  $signed(reg2057) : reg1430[(2'h2):(1'h0)]) : ((forvar2540 ?
                                      reg2160 : reg2072) ?
                                  {reg2570} : {reg1492})));
                      reg2566 <= reg2136[(3'h7):(1'h0)];
                    end
                  for (forvar2567 = (1'h0); (forvar2567 < (2'h2)); forvar2567 = (forvar2567 + (1'h1)))
                    begin
                      reg2568 <= ({(reg2185 && $unsigned(reg2504))} ?
                          reg2290 : reg1481);
                      reg2569 <= (((^$signed(wire1412)) != $signed($signed(reg1438))) ?
                          $signed(reg2112) : ({(reg2479 ?
                                  reg2326 : reg1503)} >>> {$signed(reg2440)}));
                      reg2570 <= reg2558[(1'h1):(1'h0)];
                    end
                end
              reg2576 <= (reg2445[(1'h1):(1'h0)] ?
                  $unsigned(reg2357) : reg2403[(1'h0):(1'h0)]);
              for (forvar2577 = (1'h0); (forvar2577 < (1'h0)); forvar2577 = (forvar2577 + (1'h1)))
                begin
                  reg2578 <= (&(((reg2260 ?
                          reg2324 : reg2558) && $signed(reg2487)) ?
                      reg2258 : reg2137));
                end
              for (forvar2579 = (1'h0); (forvar2579 < (2'h3)); forvar2579 = (forvar2579 + (1'h1)))
                begin
                  for (forvar2580 = (1'h0); (forvar2580 < (1'h1)); forvar2580 = (forvar2580 + (1'h1)))
                    begin
                      reg2581 <= $signed((reg2047[(3'h7):(3'h7)] ?
                          $signed(reg2505) : reg1438[(4'h8):(1'h0)]));
                      reg2582 <= ({reg2059} * (~reg2362));
                      reg2583 <= $signed({reg2225[(1'h0):(1'h0)]});
                    end
                  for (forvar2584 = (1'h0); (forvar2584 < (2'h2)); forvar2584 = (forvar2584 + (1'h1)))
                    begin
                      reg2585 <= reg2274[(4'he):(4'h8)];
                    end
                end
            end
          else
            begin
              reg2564 <= $unsigned((((reg2499 * reg2110) ?
                  (reg2389 ?
                      (8'haf) : (8'ha3)) : reg1492) == $signed((reg2046 >= reg2222))));
              if ($unsigned($signed((+(reg2473 ? reg2076 : forvar2584)))))
                begin
                  for (forvar2565 = (1'h0); (forvar2565 < (1'h1)); forvar2565 = (forvar2565 + (1'h1)))
                    begin
                      reg2566 <= (+reg2103);
                    end
                  if ((($signed((|reg1492)) ?
                          $unsigned({reg1455}) : (reg2431[(2'h3):(1'h0)] > reg1525)) ?
                      $unsigned(((reg2182 ?
                          (8'haa) : (8'ha8)) - (!reg2112))) : reg2048))
                    begin
                      reg2567 <= reg2260[(1'h1):(1'h0)];
                      reg2568 <= reg2176;
                    end
                  else
                    begin
                      reg2567 <= (((~^$unsigned(reg2523)) < (~^(reg2226 ^~ reg2360))) ?
                          $signed(reg2389[(2'h3):(1'h0)]) : reg2203);
                      reg2568 <= {$unsigned({$unsigned(reg2221)})};
                      reg2569 <= $signed(($signed(((8'h9d) ?
                              reg1514 : reg2051)) ?
                          $signed($unsigned(reg2501)) : reg2232[(3'h5):(3'h4)]));
                      reg2570 <= reg2112[(4'ha):(1'h1)];
                    end
                  for (forvar2571 = (1'h0); (forvar2571 < (2'h3)); forvar2571 = (forvar2571 + (1'h1)))
                    begin
                      reg2572 <= ((reg1431 ?
                          (reg2183[(1'h1):(1'h1)] ?
                              (reg2110 ^ reg2453) : (forvar2584 ?
                                  reg2312 : (8'ha8))) : $signed($unsigned((8'ha1)))) & $unsigned((~{reg2471})));
                      reg2573 <= {(-reg2218[(3'h7):(2'h3)])};
                      reg2574 <= reg2328[(2'h2):(1'h1)];
                      reg2575 <= $unsigned((((reg1498 ?
                              reg2348 : (8'h9c)) || {reg2169}) ?
                          reg2151 : (~|$signed(reg1519))));
                    end
                end
              else
                begin
                  for (forvar2565 = (1'h0); (forvar2565 < (2'h2)); forvar2565 = (forvar2565 + (1'h1)))
                    begin
                      reg2566 <= ({$signed(reg1450)} < (^((8'ha5) ?
                          reg1539 : reg2449[(4'ha):(1'h0)])));
                      reg2567 <= {((reg1421[(1'h0):(1'h0)] + (reg2286 ?
                                  reg1485 : reg1524)) ?
                              $signed($signed(reg1484)) : (reg2147 ?
                                  reg2051 : $signed(reg2295)))};
                      reg2568 <= reg2493;
                      reg2569 <= reg2066;
                    end
                end
              for (forvar2576 = (1'h0); (forvar2576 < (1'h0)); forvar2576 = (forvar2576 + (1'h1)))
                begin
                  reg2577 <= {reg2214[(3'h4):(2'h2)]};
                  reg2578 <= $unsigned(($unsigned(reg2343) ?
                      $signed(reg1440[(3'h4):(2'h3)]) : reg2353[(4'h8):(3'h6)]));
                  for (forvar2579 = (1'h0); (forvar2579 < (2'h3)); forvar2579 = (forvar2579 + (1'h1)))
                    begin
                      reg2580 <= (^~(~&($signed(reg2296) ?
                          {(8'hb5)} : $unsigned((8'hb3)))));
                    end
                  if ({(reg2058 ?
                          (8'hb4) : ((reg1426 ^ reg2522) ?
                              (reg1526 ?
                                  reg2403 : reg1428) : (reg2335 - reg2450)))})
                    begin
                      reg2581 <= {reg2285};
                      reg2582 <= $unsigned(reg2122);
                      reg2583 <= (reg2341[(3'h5):(1'h1)] ?
                          {{wire1412}} : $signed($unsigned((~^(8'hb5)))));
                      reg2584 <= {reg2444};
                    end
                  else
                    begin
                      reg2581 <= (~&(|($signed((8'ha7)) ?
                          $signed((8'hab)) : (^~(8'ha1)))));
                      reg2582 <= $unsigned((reg1473[(4'hd):(4'ha)] ?
                          ((!reg2132) ?
                              (~reg2384) : reg2121[(2'h2):(2'h2)]) : ((wire2331 ?
                                  reg2417 : reg2292) ?
                              (reg2085 & reg2214) : (~^reg2273))));
                      reg2583 <= reg2437[(4'hc):(1'h0)];
                    end
                end
            end
        end
      else
        begin
          reg2540 <= reg2416[(1'h0):(1'h0)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1540  (y, clk, wire1545, wire1544, wire1543, wire1542, wire1541);
  output wire [(32'h15c5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire1545;
  input wire [(2'h3):(1'h0)] wire1544;
  input wire signed [(4'h9):(1'h0)] wire1543;
  input wire signed [(4'hc):(1'h0)] wire1542;
  input wire signed [(3'h7):(1'h0)] wire1541;
  wire [(4'he):(1'h0)] wire2026;
  wire signed [(4'hd):(1'h0)] wire2025;
  wire [(5'h10):(1'h0)] wire1887;
  wire [(4'hb):(1'h0)] wire1886;
  wire signed [(3'h7):(1'h0)] wire1816;
  wire [(4'ha):(1'h0)] wire1815;
  wire signed [(4'hf):(1'h0)] wire1814;
  wire [(4'h8):(1'h0)] wire1813;
  wire [(4'hb):(1'h0)] wire1812;
  wire [(3'h6):(1'h0)] wire1771;
  wire [(4'hc):(1'h0)] wire1770;
  wire [(3'h7):(1'h0)] wire1547;
  wire [(4'hd):(1'h0)] wire1546;
  reg signed [(3'h4):(1'h0)] reg2024 = (1'h0);
  reg [(2'h2):(1'h0)] reg2023 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2022 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2020 = (1'h0);
  reg [(4'hc):(1'h0)] reg2019 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2017 = (1'h0);
  reg [(4'hc):(1'h0)] reg2016 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2015 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2012 = (1'h0);
  reg [(4'ha):(1'h0)] reg2011 = (1'h0);
  reg [(4'ha):(1'h0)] reg2010 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2009 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2007 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2006 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2005 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2004 = (1'h0);
  reg [(4'h8):(1'h0)] reg2003 = (1'h0);
  reg [(4'hb):(1'h0)] reg2002 = (1'h0);
  reg [(2'h2):(1'h0)] reg2001 = (1'h0);
  reg [(5'h10):(1'h0)] reg2000 = (1'h0);
  reg [(4'h8):(1'h0)] reg1999 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1998 = (1'h0);
  reg [(4'hc):(1'h0)] reg1997 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1995 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1994 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1993 = (1'h0);
  reg [(4'he):(1'h0)] reg1992 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1990 = (1'h0);
  reg [(3'h4):(1'h0)] reg1989 = (1'h0);
  reg [(4'hf):(1'h0)] reg1988 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1987 = (1'h0);
  reg [(3'h6):(1'h0)] reg1985 = (1'h0);
  reg [(4'hf):(1'h0)] reg1984 = (1'h0);
  reg [(3'h4):(1'h0)] reg1983 = (1'h0);
  reg [(4'h9):(1'h0)] reg1981 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1980 = (1'h0);
  reg [(4'hc):(1'h0)] reg1982 = (1'h0);
  reg [(4'he):(1'h0)] reg1979 = (1'h0);
  reg [(2'h3):(1'h0)] reg1978 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1977 = (1'h0);
  reg [(4'h9):(1'h0)] reg1976 = (1'h0);
  reg [(3'h5):(1'h0)] reg1975 = (1'h0);
  reg [(4'he):(1'h0)] reg1974 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1972 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1971 = (1'h0);
  reg [(2'h3):(1'h0)] reg1968 = (1'h0);
  reg [(2'h2):(1'h0)] reg1970 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1969 = (1'h0);
  reg [(4'hf):(1'h0)] reg1967 = (1'h0);
  reg [(4'ha):(1'h0)] reg1966 = (1'h0);
  reg [(4'h9):(1'h0)] reg1965 = (1'h0);
  reg [(4'hf):(1'h0)] reg1958 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1946 = (1'h0);
  reg [(2'h2):(1'h0)] reg1964 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1963 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1961 = (1'h0);
  reg [(5'h10):(1'h0)] reg1960 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1959 = (1'h0);
  reg [(4'h9):(1'h0)] reg1957 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1956 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1955 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1954 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1953 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1952 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1951 = (1'h0);
  reg [(4'he):(1'h0)] reg1950 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1949 = (1'h0);
  reg [(4'hf):(1'h0)] reg1948 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1947 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1945 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1944 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1943 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1937 = (1'h0);
  reg [(4'he):(1'h0)] reg1942 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1933 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1941 = (1'h0);
  reg [(4'hc):(1'h0)] reg1940 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1939 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1938 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1936 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1935 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1934 = (1'h0);
  reg [(3'h7):(1'h0)] reg1932 = (1'h0);
  reg [(4'ha):(1'h0)] reg1931 = (1'h0);
  reg [(3'h4):(1'h0)] reg1930 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1929 = (1'h0);
  reg [(4'ha):(1'h0)] reg1927 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1923 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1926 = (1'h0);
  reg [(4'hc):(1'h0)] reg1925 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1924 = (1'h0);
  reg [(4'hb):(1'h0)] reg1922 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1921 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1920 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1919 = (1'h0);
  reg [(4'h8):(1'h0)] reg1918 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1917 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1916 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1915 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1914 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1912 = (1'h0);
  reg [(2'h2):(1'h0)] reg1911 = (1'h0);
  reg [(4'hb):(1'h0)] reg1910 = (1'h0);
  reg [(4'hf):(1'h0)] reg1909 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1908 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1907 = (1'h0);
  reg [(4'hc):(1'h0)] reg1904 = (1'h0);
  reg [(3'h7):(1'h0)] reg1903 = (1'h0);
  reg [(3'h6):(1'h0)] reg1902 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1901 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1900 = (1'h0);
  reg [(5'h10):(1'h0)] reg1899 = (1'h0);
  reg [(4'hc):(1'h0)] reg1898 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1897 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1896 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1894 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1893 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1892 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1891 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1888 = (1'h0);
  reg [(4'h8):(1'h0)] reg1885 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1879 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1875 = (1'h0);
  reg [(2'h2):(1'h0)] reg1865 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1884 = (1'h0);
  reg [(3'h6):(1'h0)] reg1883 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1882 = (1'h0);
  reg [(3'h5):(1'h0)] reg1881 = (1'h0);
  reg [(2'h2):(1'h0)] reg1880 = (1'h0);
  reg [(4'hb):(1'h0)] reg1878 = (1'h0);
  reg [(5'h10):(1'h0)] reg1877 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1876 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1874 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1873 = (1'h0);
  reg [(4'hf):(1'h0)] reg1872 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1871 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1870 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1869 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1868 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1867 = (1'h0);
  reg [(4'hd):(1'h0)] reg1866 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1864 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1860 = (1'h0);
  reg [(2'h3):(1'h0)] reg1855 = (1'h0);
  reg [(4'hb):(1'h0)] reg1852 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1863 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1862 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1861 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1859 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1858 = (1'h0);
  reg [(4'hf):(1'h0)] reg1857 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1856 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1854 = (1'h0);
  reg [(4'ha):(1'h0)] reg1853 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1851 = (1'h0);
  reg [(3'h4):(1'h0)] reg1850 = (1'h0);
  reg [(4'hf):(1'h0)] reg1849 = (1'h0);
  reg [(2'h2):(1'h0)] reg1848 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1819 = (1'h0);
  reg [(5'h10):(1'h0)] reg1817 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1842 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1839 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1832 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1831 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1823 = (1'h0);
  reg [(4'ha):(1'h0)] reg1821 = (1'h0);
  reg [(2'h3):(1'h0)] reg1847 = (1'h0);
  reg [(3'h7):(1'h0)] reg1837 = (1'h0);
  reg [(3'h5):(1'h0)] reg1846 = (1'h0);
  reg [(4'hb):(1'h0)] reg1844 = (1'h0);
  reg [(3'h7):(1'h0)] reg1843 = (1'h0);
  reg [(3'h6):(1'h0)] reg1841 = (1'h0);
  reg [(4'hc):(1'h0)] reg1840 = (1'h0);
  reg [(5'h10):(1'h0)] reg1838 = (1'h0);
  reg [(3'h7):(1'h0)] reg1836 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1835 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1834 = (1'h0);
  reg [(5'h10):(1'h0)] reg1833 = (1'h0);
  reg [(4'hd):(1'h0)] reg1830 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1829 = (1'h0);
  reg [(3'h6):(1'h0)] reg1828 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1827 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1826 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1825 = (1'h0);
  reg [(3'h5):(1'h0)] reg1824 = (1'h0);
  reg [(3'h5):(1'h0)] reg1822 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1820 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1818 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1811 = (1'h0);
  reg [(3'h7):(1'h0)] reg1809 = (1'h0);
  reg [(4'hb):(1'h0)] reg1793 = (1'h0);
  reg [(4'hb):(1'h0)] reg1791 = (1'h0);
  reg [(3'h6):(1'h0)] reg1790 = (1'h0);
  reg [(2'h2):(1'h0)] reg1784 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1778 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1810 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1794 = (1'h0);
  reg [(3'h5):(1'h0)] reg1808 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1807 = (1'h0);
  reg [(3'h5):(1'h0)] reg1806 = (1'h0);
  reg [(3'h6):(1'h0)] reg1805 = (1'h0);
  reg [(4'hb):(1'h0)] reg1804 = (1'h0);
  reg [(3'h7):(1'h0)] reg1803 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1802 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1801 = (1'h0);
  reg [(4'hb):(1'h0)] reg1800 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1799 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1798 = (1'h0);
  reg [(3'h7):(1'h0)] reg1797 = (1'h0);
  reg [(4'hf):(1'h0)] reg1796 = (1'h0);
  reg [(3'h6):(1'h0)] reg1795 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1792 = (1'h0);
  reg [(4'h9):(1'h0)] reg1789 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1788 = (1'h0);
  reg [(3'h6):(1'h0)] reg1787 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1786 = (1'h0);
  reg [(5'h10):(1'h0)] reg1785 = (1'h0);
  reg [(3'h4):(1'h0)] reg1783 = (1'h0);
  reg [(4'h8):(1'h0)] reg1782 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1781 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1780 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1779 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1773 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1777 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1776 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1775 = (1'h0);
  reg [(4'hb):(1'h0)] reg1774 = (1'h0);
  reg [(4'h8):(1'h0)] reg1769 = (1'h0);
  reg [(5'h10):(1'h0)] reg1768 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1767 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1766 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1764 = (1'h0);
  reg [(5'h10):(1'h0)] reg1763 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1762 = (1'h0);
  reg [(4'hb):(1'h0)] reg1761 = (1'h0);
  reg [(4'he):(1'h0)] reg1759 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1752 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1751 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1744 = (1'h0);
  reg [(4'hc):(1'h0)] reg1743 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1741 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1738 = (1'h0);
  reg [(4'he):(1'h0)] reg1758 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1757 = (1'h0);
  reg [(2'h3):(1'h0)] reg1756 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1755 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1754 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1753 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1750 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1749 = (1'h0);
  reg [(4'he):(1'h0)] reg1747 = (1'h0);
  reg [(2'h2):(1'h0)] reg1746 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1745 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1742 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1740 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1739 = (1'h0);
  reg [(4'h9):(1'h0)] reg1737 = (1'h0);
  reg [(3'h6):(1'h0)] reg1736 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1733 = (1'h0);
  reg [(4'hb):(1'h0)] reg1732 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1731 = (1'h0);
  reg [(4'h9):(1'h0)] reg1730 = (1'h0);
  reg [(4'h9):(1'h0)] reg1729 = (1'h0);
  reg [(3'h7):(1'h0)] reg1728 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1727 = (1'h0);
  reg [(4'he):(1'h0)] reg1721 = (1'h0);
  reg [(3'h4):(1'h0)] reg1716 = (1'h0);
  reg [(4'he):(1'h0)] reg1725 = (1'h0);
  reg [(5'h10):(1'h0)] reg1724 = (1'h0);
  reg [(2'h2):(1'h0)] reg1722 = (1'h0);
  reg [(4'h8):(1'h0)] reg1720 = (1'h0);
  reg [(3'h4):(1'h0)] reg1719 = (1'h0);
  reg [(4'h8):(1'h0)] reg1718 = (1'h0);
  reg [(5'h10):(1'h0)] reg1717 = (1'h0);
  reg [(4'he):(1'h0)] reg1714 = (1'h0);
  reg [(4'h8):(1'h0)] reg1713 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1712 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1711 = (1'h0);
  reg [(4'hf):(1'h0)] reg1701 = (1'h0);
  reg [(4'h9):(1'h0)] reg1710 = (1'h0);
  reg [(4'hf):(1'h0)] reg1709 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1707 = (1'h0);
  reg [(5'h10):(1'h0)] reg1706 = (1'h0);
  reg [(4'hb):(1'h0)] reg1705 = (1'h0);
  reg [(4'ha):(1'h0)] reg1704 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1703 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1702 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1700 = (1'h0);
  reg [(4'ha):(1'h0)] reg1699 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1698 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1696 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1695 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1694 = (1'h0);
  reg [(3'h6):(1'h0)] reg1693 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1680 = (1'h0);
  reg [(4'hd):(1'h0)] reg1678 = (1'h0);
  reg [(2'h3):(1'h0)] reg1691 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1690 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1689 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1688 = (1'h0);
  reg [(2'h2):(1'h0)] reg1686 = (1'h0);
  reg [(3'h5):(1'h0)] reg1685 = (1'h0);
  reg [(4'h9):(1'h0)] reg1683 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1682 = (1'h0);
  reg [(4'h9):(1'h0)] reg1681 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1679 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1675 = (1'h0);
  reg [(3'h7):(1'h0)] reg1674 = (1'h0);
  reg [(4'hd):(1'h0)] reg1673 = (1'h0);
  reg [(4'ha):(1'h0)] reg1671 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1670 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1669 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1668 = (1'h0);
  reg [(4'ha):(1'h0)] reg1667 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1665 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1664 = (1'h0);
  reg [(4'ha):(1'h0)] reg1663 = (1'h0);
  reg [(4'ha):(1'h0)] reg1662 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1661 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1659 = (1'h0);
  reg [(2'h3):(1'h0)] reg1658 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1657 = (1'h0);
  reg [(4'hf):(1'h0)] reg1653 = (1'h0);
  reg [(4'he):(1'h0)] reg1629 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1627 = (1'h0);
  reg [(2'h3):(1'h0)] reg1622 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1619 = (1'h0);
  reg [(4'hd):(1'h0)] reg1617 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1613 = (1'h0);
  reg [(3'h7):(1'h0)] reg1611 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1654 = (1'h0);
  reg [(4'hd):(1'h0)] reg1652 = (1'h0);
  reg [(2'h3):(1'h0)] reg1651 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1650 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1649 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1648 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1641 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1647 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1646 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1645 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1644 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1643 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1642 = (1'h0);
  reg [(4'h8):(1'h0)] reg1640 = (1'h0);
  reg [(4'hb):(1'h0)] reg1639 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1633 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1636 = (1'h0);
  reg [(5'h10):(1'h0)] reg1635 = (1'h0);
  reg [(2'h2):(1'h0)] reg1634 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1632 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1631 = (1'h0);
  reg [(3'h6):(1'h0)] reg1630 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1628 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1626 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1625 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1624 = (1'h0);
  reg [(3'h4):(1'h0)] reg1623 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1621 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1620 = (1'h0);
  reg [(4'h9):(1'h0)] reg1616 = (1'h0);
  reg [(5'h10):(1'h0)] reg1615 = (1'h0);
  reg [(4'hb):(1'h0)] reg1614 = (1'h0);
  reg [(2'h2):(1'h0)] reg1612 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1610 = (1'h0);
  reg [(3'h6):(1'h0)] reg1609 = (1'h0);
  reg [(4'hd):(1'h0)] reg1608 = (1'h0);
  reg [(4'he):(1'h0)] reg1607 = (1'h0);
  reg [(4'hf):(1'h0)] reg1606 = (1'h0);
  reg [(4'hd):(1'h0)] reg1591 = (1'h0);
  reg [(3'h5):(1'h0)] reg1590 = (1'h0);
  reg [(5'h10):(1'h0)] reg1588 = (1'h0);
  reg [(5'h10):(1'h0)] reg1584 = (1'h0);
  reg [(3'h7):(1'h0)] reg1603 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1602 = (1'h0);
  reg [(4'hf):(1'h0)] reg1601 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1600 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1599 = (1'h0);
  reg [(4'hb):(1'h0)] reg1598 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1597 = (1'h0);
  reg [(2'h2):(1'h0)] reg1596 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1595 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1594 = (1'h0);
  reg [(4'h8):(1'h0)] reg1593 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1592 = (1'h0);
  reg [(2'h3):(1'h0)] reg1589 = (1'h0);
  reg [(4'h9):(1'h0)] reg1587 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1586 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1585 = (1'h0);
  reg [(4'h9):(1'h0)] reg1583 = (1'h0);
  reg [(4'ha):(1'h0)] reg1582 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1581 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1580 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1579 = (1'h0);
  reg [(3'h4):(1'h0)] reg1577 = (1'h0);
  reg [(4'h9):(1'h0)] reg1556 = (1'h0);
  reg [(4'hd):(1'h0)] reg1576 = (1'h0);
  reg [(3'h5):(1'h0)] reg1575 = (1'h0);
  reg [(3'h6):(1'h0)] reg1574 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1573 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1572 = (1'h0);
  reg [(4'h8):(1'h0)] reg1571 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1570 = (1'h0);
  reg [(4'hf):(1'h0)] reg1568 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1567 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1566 = (1'h0);
  reg [(3'h4):(1'h0)] reg1563 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1562 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1561 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1549 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1558 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1557 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1555 = (1'h0);
  reg [(4'hf):(1'h0)] reg1554 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1553 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1552 = (1'h0);
  reg [(2'h2):(1'h0)] reg1551 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1550 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2021 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2018 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2014 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2013 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2008 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2003 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1996 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1991 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1986 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1982 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1979 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1978 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1981 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1980 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1973 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1964 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1968 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1957 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1951 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1950 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1962 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1954 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1958 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1946 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1942 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1941 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1931 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1916 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1920 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1907 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1932 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1937 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1933 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1928 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1926 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1922 = (1'h0);
  reg [(4'he):(1'h0)] forvar1924 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1921 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1918 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1923 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1913 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1906 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1905 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1895 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1890 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1889 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1876 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1870 = (1'h0);
  reg [(4'he):(1'h0)] forvar1872 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1866 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1879 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1875 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1865 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1861 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1859 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1860 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1855 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1852 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1846 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1834 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1826 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1818 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1840 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1828 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1824 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1820 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1845 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1842 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1839 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1837 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1832 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1831 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1823 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1821 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1819 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1817 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1806 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1803 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1799 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1797 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1788 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1782 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1775 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1809 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1795 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1794 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1793 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1791 = (1'h0);
  reg [(4'he):(1'h0)] forvar1790 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1784 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1778 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1773 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1772 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1765 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1760 = (1'h0);
  reg [(4'he):(1'h0)] forvar1756 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1754 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1745 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1752 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1751 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1748 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1744 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1743 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1741 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1738 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1735 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1734 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1727 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1726 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1719 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1723 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1721 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1716 = (1'h0);
  reg [(4'he):(1'h0)] forvar1715 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1708 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1701 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1694 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1697 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1692 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1679 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1687 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1684 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1680 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1678 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1677 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1676 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1672 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1666 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1660 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1656 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1655 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1643 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1628 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1623 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1610 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1608 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1653 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1640 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1641 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1638 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1637 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1633 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1629 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1627 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1622 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1619 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1618 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1617 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1613 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1611 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1605 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1604 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1598 = (1'h0);
  reg [(4'he):(1'h0)] forvar1594 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1589 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1585 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1591 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1590 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1588 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1584 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1578 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1557 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1550 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1569 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1565 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1564 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1560 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1559 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1556 = (1'h0);
  reg [(4'he):(1'h0)] forvar1549 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1548 = (1'h0);
  assign y = {wire2026,
                 wire2025,
                 wire1887,
                 wire1886,
                 wire1816,
                 wire1815,
                 wire1814,
                 wire1813,
                 wire1812,
                 wire1771,
                 wire1770,
                 wire1547,
                 wire1546,
                 reg2024,
                 reg2023,
                 reg2022,
                 reg2020,
                 reg2019,
                 reg2017,
                 reg2016,
                 reg2015,
                 reg2012,
                 reg2011,
                 reg2010,
                 reg2009,
                 reg2007,
                 reg2006,
                 reg2005,
                 reg2004,
                 reg2003,
                 reg2002,
                 reg2001,
                 reg2000,
                 reg1999,
                 reg1998,
                 reg1997,
                 reg1995,
                 reg1994,
                 reg1993,
                 reg1992,
                 reg1990,
                 reg1989,
                 reg1988,
                 reg1987,
                 reg1985,
                 reg1984,
                 reg1983,
                 reg1981,
                 reg1980,
                 reg1982,
                 reg1979,
                 reg1978,
                 reg1977,
                 reg1976,
                 reg1975,
                 reg1974,
                 reg1972,
                 reg1971,
                 reg1968,
                 reg1970,
                 reg1969,
                 reg1967,
                 reg1966,
                 reg1965,
                 reg1958,
                 reg1946,
                 reg1964,
                 reg1963,
                 reg1961,
                 reg1960,
                 reg1959,
                 reg1957,
                 reg1956,
                 reg1955,
                 reg1954,
                 reg1953,
                 reg1952,
                 reg1951,
                 reg1950,
                 reg1949,
                 reg1948,
                 reg1947,
                 reg1945,
                 reg1944,
                 reg1943,
                 reg1937,
                 reg1942,
                 reg1933,
                 reg1941,
                 reg1940,
                 reg1939,
                 reg1938,
                 reg1936,
                 reg1935,
                 reg1934,
                 reg1932,
                 reg1931,
                 reg1930,
                 reg1929,
                 reg1927,
                 reg1923,
                 reg1926,
                 reg1925,
                 reg1924,
                 reg1922,
                 reg1921,
                 reg1920,
                 reg1919,
                 reg1918,
                 reg1917,
                 reg1916,
                 reg1915,
                 reg1914,
                 reg1912,
                 reg1911,
                 reg1910,
                 reg1909,
                 reg1908,
                 reg1907,
                 reg1904,
                 reg1903,
                 reg1902,
                 reg1901,
                 reg1900,
                 reg1899,
                 reg1898,
                 reg1897,
                 reg1896,
                 reg1894,
                 reg1893,
                 reg1892,
                 reg1891,
                 reg1888,
                 reg1885,
                 reg1879,
                 reg1875,
                 reg1865,
                 reg1884,
                 reg1883,
                 reg1882,
                 reg1881,
                 reg1880,
                 reg1878,
                 reg1877,
                 reg1876,
                 reg1874,
                 reg1873,
                 reg1872,
                 reg1871,
                 reg1870,
                 reg1869,
                 reg1868,
                 reg1867,
                 reg1866,
                 reg1864,
                 reg1860,
                 reg1855,
                 reg1852,
                 reg1863,
                 reg1862,
                 reg1861,
                 reg1859,
                 reg1858,
                 reg1857,
                 reg1856,
                 reg1854,
                 reg1853,
                 reg1851,
                 reg1850,
                 reg1849,
                 reg1848,
                 reg1819,
                 reg1817,
                 reg1842,
                 reg1839,
                 reg1832,
                 reg1831,
                 reg1823,
                 reg1821,
                 reg1847,
                 reg1837,
                 reg1846,
                 reg1844,
                 reg1843,
                 reg1841,
                 reg1840,
                 reg1838,
                 reg1836,
                 reg1835,
                 reg1834,
                 reg1833,
                 reg1830,
                 reg1829,
                 reg1828,
                 reg1827,
                 reg1826,
                 reg1825,
                 reg1824,
                 reg1822,
                 reg1820,
                 reg1818,
                 reg1811,
                 reg1809,
                 reg1793,
                 reg1791,
                 reg1790,
                 reg1784,
                 reg1778,
                 reg1810,
                 reg1794,
                 reg1808,
                 reg1807,
                 reg1806,
                 reg1805,
                 reg1804,
                 reg1803,
                 reg1802,
                 reg1801,
                 reg1800,
                 reg1799,
                 reg1798,
                 reg1797,
                 reg1796,
                 reg1795,
                 reg1792,
                 reg1789,
                 reg1788,
                 reg1787,
                 reg1786,
                 reg1785,
                 reg1783,
                 reg1782,
                 reg1781,
                 reg1780,
                 reg1779,
                 reg1773,
                 reg1777,
                 reg1776,
                 reg1775,
                 reg1774,
                 reg1769,
                 reg1768,
                 reg1767,
                 reg1766,
                 reg1764,
                 reg1763,
                 reg1762,
                 reg1761,
                 reg1759,
                 reg1752,
                 reg1751,
                 reg1744,
                 reg1743,
                 reg1741,
                 reg1738,
                 reg1758,
                 reg1757,
                 reg1756,
                 reg1755,
                 reg1754,
                 reg1753,
                 reg1750,
                 reg1749,
                 reg1747,
                 reg1746,
                 reg1745,
                 reg1742,
                 reg1740,
                 reg1739,
                 reg1737,
                 reg1736,
                 reg1733,
                 reg1732,
                 reg1731,
                 reg1730,
                 reg1729,
                 reg1728,
                 reg1727,
                 reg1721,
                 reg1716,
                 reg1725,
                 reg1724,
                 reg1722,
                 reg1720,
                 reg1719,
                 reg1718,
                 reg1717,
                 reg1714,
                 reg1713,
                 reg1712,
                 reg1711,
                 reg1701,
                 reg1710,
                 reg1709,
                 reg1707,
                 reg1706,
                 reg1705,
                 reg1704,
                 reg1703,
                 reg1702,
                 reg1700,
                 reg1699,
                 reg1698,
                 reg1696,
                 reg1695,
                 reg1694,
                 reg1693,
                 reg1680,
                 reg1678,
                 reg1691,
                 reg1690,
                 reg1689,
                 reg1688,
                 reg1686,
                 reg1685,
                 reg1683,
                 reg1682,
                 reg1681,
                 reg1679,
                 reg1675,
                 reg1674,
                 reg1673,
                 reg1671,
                 reg1670,
                 reg1669,
                 reg1668,
                 reg1667,
                 reg1665,
                 reg1664,
                 reg1663,
                 reg1662,
                 reg1661,
                 reg1659,
                 reg1658,
                 reg1657,
                 reg1653,
                 reg1629,
                 reg1627,
                 reg1622,
                 reg1619,
                 reg1617,
                 reg1613,
                 reg1611,
                 reg1654,
                 reg1652,
                 reg1651,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1641,
                 reg1647,
                 reg1646,
                 reg1645,
                 reg1644,
                 reg1643,
                 reg1642,
                 reg1640,
                 reg1639,
                 reg1633,
                 reg1636,
                 reg1635,
                 reg1634,
                 reg1632,
                 reg1631,
                 reg1630,
                 reg1628,
                 reg1626,
                 reg1625,
                 reg1624,
                 reg1623,
                 reg1621,
                 reg1620,
                 reg1616,
                 reg1615,
                 reg1614,
                 reg1612,
                 reg1610,
                 reg1609,
                 reg1608,
                 reg1607,
                 reg1606,
                 reg1591,
                 reg1590,
                 reg1588,
                 reg1584,
                 reg1603,
                 reg1602,
                 reg1601,
                 reg1600,
                 reg1599,
                 reg1598,
                 reg1597,
                 reg1596,
                 reg1595,
                 reg1594,
                 reg1593,
                 reg1592,
                 reg1589,
                 reg1587,
                 reg1586,
                 reg1585,
                 reg1583,
                 reg1582,
                 reg1581,
                 reg1580,
                 reg1579,
                 reg1577,
                 reg1556,
                 reg1576,
                 reg1575,
                 reg1574,
                 reg1573,
                 reg1572,
                 reg1571,
                 reg1570,
                 reg1568,
                 reg1567,
                 reg1566,
                 reg1563,
                 reg1562,
                 reg1561,
                 reg1549,
                 reg1558,
                 reg1557,
                 reg1555,
                 reg1554,
                 reg1553,
                 reg1552,
                 reg1551,
                 reg1550,
                 forvar2021,
                 forvar2018,
                 forvar2014,
                 forvar2013,
                 forvar2008,
                 forvar2003,
                 forvar1996,
                 forvar1991,
                 forvar1986,
                 forvar1982,
                 forvar1979,
                 forvar1978,
                 forvar1981,
                 forvar1980,
                 forvar1973,
                 forvar1964,
                 forvar1968,
                 forvar1957,
                 forvar1951,
                 forvar1950,
                 forvar1962,
                 forvar1954,
                 forvar1958,
                 forvar1946,
                 forvar1942,
                 forvar1941,
                 forvar1931,
                 forvar1916,
                 forvar1920,
                 forvar1907,
                 forvar1932,
                 forvar1937,
                 forvar1933,
                 forvar1928,
                 forvar1926,
                 forvar1922,
                 forvar1924,
                 forvar1921,
                 forvar1918,
                 forvar1923,
                 forvar1913,
                 forvar1906,
                 forvar1905,
                 forvar1895,
                 forvar1890,
                 forvar1889,
                 forvar1876,
                 forvar1870,
                 forvar1872,
                 forvar1866,
                 forvar1879,
                 forvar1875,
                 forvar1865,
                 forvar1861,
                 forvar1859,
                 forvar1860,
                 forvar1855,
                 forvar1852,
                 forvar1846,
                 forvar1834,
                 forvar1826,
                 forvar1818,
                 forvar1840,
                 forvar1828,
                 forvar1824,
                 forvar1820,
                 forvar1845,
                 forvar1842,
                 forvar1839,
                 forvar1837,
                 forvar1832,
                 forvar1831,
                 forvar1823,
                 forvar1821,
                 forvar1819,
                 forvar1817,
                 forvar1806,
                 forvar1803,
                 forvar1799,
                 forvar1797,
                 forvar1788,
                 forvar1782,
                 forvar1775,
                 forvar1809,
                 forvar1795,
                 forvar1794,
                 forvar1793,
                 forvar1791,
                 forvar1790,
                 forvar1784,
                 forvar1778,
                 forvar1773,
                 forvar1772,
                 forvar1765,
                 forvar1760,
                 forvar1756,
                 forvar1754,
                 forvar1745,
                 forvar1752,
                 forvar1751,
                 forvar1748,
                 forvar1744,
                 forvar1743,
                 forvar1741,
                 forvar1738,
                 forvar1735,
                 forvar1734,
                 forvar1727,
                 forvar1726,
                 forvar1719,
                 forvar1723,
                 forvar1721,
                 forvar1716,
                 forvar1715,
                 forvar1708,
                 forvar1701,
                 forvar1694,
                 forvar1697,
                 forvar1692,
                 forvar1679,
                 forvar1687,
                 forvar1684,
                 forvar1680,
                 forvar1678,
                 forvar1677,
                 forvar1676,
                 forvar1672,
                 forvar1666,
                 forvar1660,
                 forvar1656,
                 forvar1655,
                 forvar1643,
                 forvar1628,
                 forvar1623,
                 forvar1610,
                 forvar1608,
                 forvar1653,
                 forvar1640,
                 forvar1641,
                 forvar1638,
                 forvar1637,
                 forvar1633,
                 forvar1629,
                 forvar1627,
                 forvar1622,
                 forvar1619,
                 forvar1618,
                 forvar1617,
                 forvar1613,
                 forvar1611,
                 forvar1605,
                 forvar1604,
                 forvar1598,
                 forvar1594,
                 forvar1589,
                 forvar1585,
                 forvar1591,
                 forvar1590,
                 forvar1588,
                 forvar1584,
                 forvar1578,
                 forvar1557,
                 forvar1550,
                 forvar1569,
                 forvar1565,
                 forvar1564,
                 forvar1560,
                 forvar1559,
                 forvar1556,
                 forvar1549,
                 forvar1548,
                 (1'h0)};
  assign wire1546 = ($signed(wire1544[(2'h2):(1'h0)]) >>> ({$unsigned(wire1542)} || ((!wire1544) << {wire1541})));
  assign wire1547 = ($unsigned($unsigned((~wire1542))) ?
                        {$unsigned($unsigned(wire1545))} : $unsigned(wire1546[(3'h5):(3'h4)]));
  always
    @(posedge clk) begin
      for (forvar1548 = (1'h0); (forvar1548 < (1'h0)); forvar1548 = (forvar1548 + (1'h1)))
        begin
          if ($unsigned({(wire1544[(1'h0):(1'h0)] * $unsigned(wire1545))}))
            begin
              if (wire1542)
                begin
                  for (forvar1549 = (1'h0); (forvar1549 < (2'h3)); forvar1549 = (forvar1549 + (1'h1)))
                    begin
                      reg1550 <= {wire1545[(2'h3):(1'h1)]};
                      reg1551 <= $signed($unsigned((+(wire1547 ?
                          wire1541 : wire1546))));
                      reg1552 <= (((8'h9f) ?
                              {(forvar1548 ?
                                      forvar1548 : wire1541)} : (8'ha9)) ?
                          $signed(((wire1543 ? wire1541 : wire1547) ?
                              (reg1550 ^ reg1550) : (wire1546 != reg1551))) : $signed(wire1546[(1'h1):(1'h0)]));
                      reg1553 <= (reg1552 ?
                          (^wire1545[(2'h2):(1'h0)]) : reg1550[(1'h1):(1'h1)]);
                    end
                  reg1554 <= {$unsigned(wire1547)};
                  if ($unsigned((forvar1549[(4'h9):(2'h3)] ?
                      (forvar1549 > {wire1543}) : $signed((reg1550 ?
                          wire1544 : forvar1549)))))
                    begin
                      reg1555 <= (^~{($signed(reg1554) >= (!reg1552))});
                    end
                  else
                    begin
                      reg1555 <= {$unsigned((reg1554[(4'h8):(3'h7)] >>> (reg1554 <= (8'h9c))))};
                    end
                  for (forvar1556 = (1'h0); (forvar1556 < (1'h1)); forvar1556 = (forvar1556 + (1'h1)))
                    begin
                      reg1557 <= $signed((~^wire1545));
                      reg1558 <= {(reg1553 ?
                              reg1551 : $signed($unsigned(wire1546)))};
                    end
                end
              else
                begin
                  if (forvar1549)
                    begin
                      reg1549 <= reg1552;
                      reg1550 <= $signed($signed(wire1543[(3'h6):(3'h6)]));
                      reg1551 <= (-($unsigned((|reg1553)) ^~ forvar1548[(3'h6):(1'h1)]));
                    end
                  else
                    begin
                      reg1549 <= (&$signed(wire1546[(2'h2):(1'h0)]));
                      reg1550 <= (($unsigned($signed(reg1554)) ~^ reg1557) ?
                          (($unsigned((8'ha9)) != {wire1547}) ?
                              reg1558 : ($signed(reg1549) << forvar1549[(4'h9):(3'h6)])) : forvar1549[(4'hb):(2'h3)]);
                      reg1551 <= (8'h9f);
                    end
                end
              for (forvar1559 = (1'h0); (forvar1559 < (2'h2)); forvar1559 = (forvar1559 + (1'h1)))
                begin
                  for (forvar1560 = (1'h0); (forvar1560 < (1'h0)); forvar1560 = (forvar1560 + (1'h1)))
                    begin
                      reg1561 <= $unsigned(forvar1559[(2'h3):(1'h1)]);
                      reg1562 <= forvar1549;
                      reg1563 <= (forvar1556 ?
                          $unsigned({wire1541[(3'h6):(3'h6)]}) : $unsigned($unsigned((~wire1547))));
                    end
                end
              for (forvar1564 = (1'h0); (forvar1564 < (1'h1)); forvar1564 = (forvar1564 + (1'h1)))
                begin
                  for (forvar1565 = (1'h0); (forvar1565 < (2'h2)); forvar1565 = (forvar1565 + (1'h1)))
                    begin
                      reg1566 <= $unsigned((((reg1550 > (8'hae)) < reg1553[(4'hd):(4'hc)]) <= {(reg1561 ?
                              (8'hb4) : forvar1559)}));
                      reg1567 <= (^$unsigned($signed((reg1561 && reg1562))));
                      reg1568 <= reg1558;
                    end
                  for (forvar1569 = (1'h0); (forvar1569 < (1'h1)); forvar1569 = (forvar1569 + (1'h1)))
                    begin
                      reg1570 <= (($signed((reg1568 >> (8'hb7))) >> $unsigned($unsigned(reg1554))) != ($signed((^wire1547)) && $unsigned((reg1563 ?
                          (8'hb1) : (8'ha3)))));
                      reg1571 <= forvar1549;
                      reg1572 <= (+forvar1569[(1'h0):(1'h0)]);
                      reg1573 <= ((reg1566[(3'h4):(2'h2)] ^ (~wire1545)) ?
                          $unsigned(wire1542[(3'h4):(2'h3)]) : reg1563[(3'h4):(1'h1)]);
                    end
                  if ($unsigned((($unsigned(wire1541) ?
                          $unsigned((8'ha6)) : $signed((8'hb8))) ?
                      ($signed((8'hb2)) >= $signed((8'haa))) : ($signed(wire1545) ?
                          (wire1546 || wire1542) : {(8'hae)}))))
                    begin
                      reg1574 <= (reg1561[(4'h8):(3'h6)] ?
                          forvar1565[(1'h0):(1'h0)] : reg1570);
                      reg1575 <= {(((8'hb2) ?
                                  forvar1549 : (reg1558 ? reg1553 : reg1573)) ?
                              wire1543[(1'h1):(1'h1)] : (reg1551[(1'h0):(1'h0)] ?
                                  $unsigned(forvar1556) : wire1545[(1'h1):(1'h0)]))};
                      reg1576 <= reg1566[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1574 <= $unsigned((8'ha1));
                    end
                end
            end
          else
            begin
              for (forvar1549 = (1'h0); (forvar1549 < (1'h0)); forvar1549 = (forvar1549 + (1'h1)))
                begin
                  for (forvar1550 = (1'h0); (forvar1550 < (2'h2)); forvar1550 = (forvar1550 + (1'h1)))
                    begin
                      reg1551 <= reg1568;
                      reg1552 <= (8'hb8);
                    end
                  if ($unsigned(wire1544[(1'h1):(1'h1)]))
                    begin
                      reg1553 <= {forvar1564[(3'h5):(2'h3)]};
                      reg1554 <= $signed((-{$signed(reg1550)}));
                      reg1555 <= wire1541[(1'h0):(1'h0)];
                      reg1556 <= {wire1544};
                    end
                  else
                    begin
                      reg1553 <= reg1556;
                    end
                  for (forvar1557 = (1'h0); (forvar1557 < (2'h2)); forvar1557 = (forvar1557 + (1'h1)))
                    begin
                      reg1558 <= {(reg1568 ?
                              reg1572[(4'h8):(3'h4)] : reg1558[(3'h6):(3'h5)])};
                    end
                end
            end
          reg1577 <= (|reg1563[(2'h2):(1'h1)]);
          for (forvar1578 = (1'h0); (forvar1578 < (1'h1)); forvar1578 = (forvar1578 + (1'h1)))
            begin
              reg1579 <= (forvar1549[(4'hc):(2'h3)] < $signed($signed((-wire1543))));
            end
          if ((&($signed(reg1566) ? (8'ha3) : $signed($unsigned(reg1558)))))
            begin
              if ($signed(reg1573[(4'hb):(3'h5)]))
                begin
                  if ($signed(reg1579[(3'h6):(2'h2)]))
                    begin
                      reg1580 <= $unsigned((^(!reg1549)));
                      reg1581 <= (|(8'hab));
                      reg1582 <= reg1574;
                    end
                  else
                    begin
                      reg1580 <= wire1547[(1'h0):(1'h0)];
                      reg1581 <= (!forvar1564[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  if ($signed(wire1546[(4'h8):(1'h0)]))
                    begin
                      reg1580 <= reg1562;
                      reg1581 <= forvar1578;
                      reg1582 <= reg1582;
                      reg1583 <= forvar1560[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg1580 <= reg1572[(3'h5):(1'h1)];
                      reg1581 <= (^~wire1544[(2'h3):(1'h0)]);
                      reg1582 <= reg1570[(4'h8):(1'h1)];
                      reg1583 <= ({$signed(((8'hae) | forvar1556))} ?
                          $unsigned(((reg1552 + wire1545) ?
                              reg1558 : (~reg1550))) : {({forvar1560} == (|forvar1565))});
                    end
                  for (forvar1584 = (1'h0); (forvar1584 < (1'h0)); forvar1584 = (forvar1584 + (1'h1)))
                    begin
                      reg1585 <= ($signed(reg1567) ^ reg1582[(4'h9):(2'h3)]);
                      reg1586 <= ($unsigned(({(8'ha2)} ?
                          reg1572[(4'ha):(3'h7)] : (~|wire1543))) || $unsigned((~^reg1574[(3'h4):(1'h0)])));
                      reg1587 <= ((!(-$unsigned(reg1561))) > ($signed(forvar1569) ^~ wire1545[(1'h0):(1'h0)]));
                    end
                end
              for (forvar1588 = (1'h0); (forvar1588 < (2'h2)); forvar1588 = (forvar1588 + (1'h1)))
                begin
                  reg1589 <= $unsigned(reg1556);
                end
              for (forvar1590 = (1'h0); (forvar1590 < (2'h2)); forvar1590 = (forvar1590 + (1'h1)))
                begin
                  for (forvar1591 = (1'h0); (forvar1591 < (1'h1)); forvar1591 = (forvar1591 + (1'h1)))
                    begin
                      reg1592 <= forvar1557[(2'h2):(1'h1)];
                    end
                  if ((8'hb4))
                    begin
                      reg1593 <= ((forvar1565 ?
                              forvar1565[(1'h0):(1'h0)] : ($unsigned(forvar1557) || reg1585[(1'h0):(1'h0)])) ?
                          $unsigned(({wire1544} ?
                              $unsigned((8'hac)) : $signed(forvar1590))) : reg1576);
                    end
                  else
                    begin
                      reg1593 <= (forvar1591[(1'h0):(1'h0)] ?
                          forvar1550 : $signed($signed((^~forvar1584))));
                      reg1594 <= ($unsigned(({(8'ha2)} ?
                              (forvar1560 || wire1541) : $signed(wire1546))) ?
                          (^$signed($unsigned(reg1576))) : (((reg1589 ~^ wire1541) ?
                                  reg1571[(1'h0):(1'h0)] : (8'ha6)) ?
                              (reg1586 ?
                                  $unsigned(reg1572) : wire1545) : {forvar1588}));
                      reg1595 <= $unsigned((!$unsigned($signed(reg1585))));
                      reg1596 <= reg1557[(3'h5):(1'h0)];
                    end
                  if ($signed($unsigned(reg1557[(1'h1):(1'h0)])))
                    begin
                      reg1597 <= $signed($signed(reg1579[(3'h7):(1'h0)]));
                      reg1598 <= (((~&$unsigned(reg1554)) ?
                          (forvar1557 ?
                              (reg1580 != reg1567) : $unsigned(reg1558)) : forvar1591[(1'h1):(1'h1)]) & $signed((8'haa)));
                      reg1599 <= $signed(((8'hab) + $unsigned({forvar1557})));
                      reg1600 <= {$unsigned(((reg1561 ?
                              wire1543 : reg1574) == reg1566))};
                    end
                  else
                    begin
                      reg1597 <= ((((forvar1584 ? reg1586 : (8'h9c)) ?
                                  $unsigned(reg1582) : $unsigned(wire1544)) ?
                              $unsigned((+reg1580)) : reg1597) ?
                          forvar1578 : $signed(reg1567[(4'hb):(2'h2)]));
                      reg1598 <= $signed(wire1546[(3'h6):(3'h4)]);
                      reg1599 <= forvar1591[(2'h2):(1'h0)];
                      reg1600 <= ($signed((reg1587[(1'h1):(1'h1)] ?
                          $unsigned(reg1587) : forvar1549)) < (~^(~$unsigned(reg1563))));
                    end
                  if (reg1553[(4'hf):(1'h1)])
                    begin
                      reg1601 <= {($signed(reg1554) | reg1585[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg1601 <= {{($signed(reg1555) ?
                                  $unsigned(wire1547) : $signed(forvar1569))}};
                      reg1602 <= forvar1556;
                      reg1603 <= ((((reg1602 >>> forvar1578) ~^ (!forvar1557)) ?
                              forvar1565[(1'h0):(1'h0)] : $unsigned(reg1566)) ?
                          (((reg1561 * reg1594) ?
                                  (reg1592 ? reg1595 : forvar1569) : reg1585) ?
                              reg1572[(1'h1):(1'h0)] : (&$signed(reg1577))) : forvar1549);
                    end
                end
            end
          else
            begin
              if ($signed($signed(((forvar1591 ? forvar1557 : reg1580) ?
                  (reg1601 ? forvar1556 : forvar1578) : $signed(forvar1569)))))
                begin
                  if ($signed(reg1575[(3'h5):(3'h5)]))
                    begin
                      reg1580 <= (forvar1588 ?
                          reg1592[(1'h1):(1'h1)] : wire1546[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg1580 <= $unsigned((~$unsigned((forvar1590 >= reg1555))));
                      reg1581 <= forvar1591[(1'h1):(1'h0)];
                      reg1582 <= $unsigned(wire1546);
                      reg1583 <= (forvar1569 <<< {reg1571});
                    end
                  for (forvar1584 = (1'h0); (forvar1584 < (1'h1)); forvar1584 = (forvar1584 + (1'h1)))
                    begin
                      reg1585 <= $unsigned((($signed(reg1562) ?
                          (&forvar1588) : (reg1562 && forvar1560)) >= reg1552[(3'h5):(2'h3)]));
                    end
                end
              else
                begin
                  if ((8'hb8))
                    begin
                      reg1580 <= ($unsigned((~&(reg1562 && (8'ha7)))) != {((8'ha5) ?
                              $unsigned(forvar1557) : (forvar1578 ?
                                  reg1553 : reg1567))});
                    end
                  else
                    begin
                      reg1580 <= (({(+wire1542)} ?
                              $signed(forvar1556) : wire1542[(3'h4):(1'h1)]) ?
                          (~^reg1582) : reg1600);
                      reg1581 <= $signed($unsigned(reg1550));
                    end
                  if ((!(^~($signed((8'ha8)) ^~ $unsigned(reg1598)))))
                    begin
                      reg1582 <= (8'h9c);
                      reg1583 <= reg1568;
                    end
                  else
                    begin
                      reg1582 <= $signed(((&(~reg1576)) <<< {reg1573}));
                      reg1583 <= {(8'hb3)};
                      reg1584 <= reg1563;
                    end
                  for (forvar1585 = (1'h0); (forvar1585 < (1'h1)); forvar1585 = (forvar1585 + (1'h1)))
                    begin
                      reg1586 <= $signed((forvar1550[(1'h1):(1'h0)] > {forvar1585[(1'h0):(1'h0)]}));
                      reg1587 <= $signed({($unsigned(reg1551) ?
                              $signed(reg1592) : (reg1580 ?
                                  forvar1556 : reg1602))});
                      reg1588 <= (($unsigned({reg1595}) ?
                          ((8'hac) ?
                              ((8'hb6) ?
                                  reg1556 : (8'ha6)) : $unsigned(reg1572)) : $unsigned({reg1570})) >= forvar1585[(1'h1):(1'h1)]);
                    end
                  for (forvar1589 = (1'h0); (forvar1589 < (2'h3)); forvar1589 = (forvar1589 + (1'h1)))
                    begin
                      reg1590 <= wire1543;
                      reg1591 <= $unsigned(reg1596);
                      reg1592 <= (($signed(wire1546) | $unsigned($signed(reg1591))) ?
                          $signed(($signed(reg1562) ^~ forvar1557)) : $unsigned($signed($signed(reg1555))));
                    end
                end
              if (((|(^reg1572)) & ({(wire1544 ?
                      reg1586 : reg1555)} & $signed(reg1593))))
                begin
                  if ((-$signed(($signed(forvar1560) <= reg1551))))
                    begin
                      reg1593 <= $unsigned($signed((&$signed(reg1584))));
                    end
                  else
                    begin
                      reg1593 <= reg1550[(1'h1):(1'h1)];
                    end
                  reg1594 <= $signed(($signed($signed(forvar1590)) ?
                      reg1601 : $signed((+reg1576))));
                  if (reg1566[(1'h1):(1'h0)])
                    begin
                      reg1595 <= (|(((wire1547 * (8'hb5)) ?
                          reg1603[(3'h6):(3'h4)] : (|forvar1569)) >> ($unsigned((8'h9d)) & (forvar1564 ?
                          forvar1564 : (8'haa)))));
                    end
                  else
                    begin
                      reg1595 <= reg1601[(4'hd):(2'h2)];
                      reg1596 <= ($unsigned(reg1586[(4'hf):(2'h2)]) ~^ (~|((^reg1570) ?
                          $signed(reg1550) : forvar1591)));
                    end
                  reg1597 <= $signed((reg1601 << $signed($unsigned(forvar1556))));
                end
              else
                begin
                  reg1593 <= ((~|{((8'hb5) & forvar1589)}) >>> reg1567);
                  for (forvar1594 = (1'h0); (forvar1594 < (2'h2)); forvar1594 = (forvar1594 + (1'h1)))
                    begin
                      reg1595 <= $signed((({reg1592} ?
                              $signed(reg1563) : (8'h9c)) ?
                          (^$signed(reg1589)) : (&(8'haf))));
                      reg1596 <= (($signed((^~forvar1557)) ?
                              reg1549[(1'h1):(1'h1)] : ((reg1566 ^ reg1580) << $unsigned(reg1555))) ?
                          reg1550[(2'h2):(1'h0)] : reg1577[(2'h3):(1'h1)]);
                      reg1597 <= reg1563;
                    end
                end
              for (forvar1598 = (1'h0); (forvar1598 < (1'h1)); forvar1598 = (forvar1598 + (1'h1)))
                begin
                  if ($signed(reg1573[(4'h9):(3'h6)]))
                    begin
                      reg1599 <= wire1545[(1'h1):(1'h1)];
                      reg1600 <= $signed((forvar1564 < reg1589[(2'h3):(2'h2)]));
                      reg1601 <= ($signed(($signed(reg1555) >>> $unsigned((8'ha5)))) != (reg1561 ?
                          ((reg1602 ?
                              (8'h9d) : reg1587) >>> {(8'hba)}) : (|(reg1585 <= reg1570))));
                    end
                  else
                    begin
                      reg1599 <= $unsigned(reg1598[(4'h8):(3'h4)]);
                      reg1600 <= $unsigned((!reg1592));
                    end
                end
            end
        end
      if ($unsigned($signed((&(forvar1588 > forvar1556)))))
        begin
          for (forvar1604 = (1'h0); (forvar1604 < (2'h3)); forvar1604 = (forvar1604 + (1'h1)))
            begin
              if ((($unsigned(reg1575[(3'h5):(1'h0)]) ?
                      ((8'ha5) ?
                          forvar1604[(4'hb):(1'h1)] : (-reg1582)) : (reg1567[(4'hc):(3'h7)] ?
                          forvar1549[(3'h4):(1'h1)] : $unsigned(reg1571))) ?
                  ({reg1570[(4'h8):(1'h0)]} + $signed((8'hab))) : $unsigned((!forvar1569[(2'h2):(1'h1)]))))
                begin
                  for (forvar1605 = (1'h0); (forvar1605 < (2'h2)); forvar1605 = (forvar1605 + (1'h1)))
                    begin
                      reg1606 <= (reg1598[(1'h1):(1'h1)] ?
                          {($signed(forvar1590) ?
                                  wire1547 : (wire1546 + reg1602))} : ({((8'h9f) ?
                                  reg1593 : forvar1589)} >>> $signed(reg1555)));
                      reg1607 <= forvar1556;
                    end
                  if ((reg1598[(3'h7):(3'h4)] ?
                      {$signed($signed(reg1561))} : forvar1588))
                    begin
                      reg1608 <= reg1596;
                      reg1609 <= $unsigned(((^reg1586) ?
                          (^((8'hb0) > reg1554)) : $signed((forvar1569 ?
                              reg1580 : reg1593))));
                    end
                  else
                    begin
                      reg1608 <= (^~(~^(&{reg1579})));
                      reg1609 <= $signed((+$signed((~wire1547))));
                      reg1610 <= (+(^(-$signed(reg1567))));
                    end
                  for (forvar1611 = (1'h0); (forvar1611 < (2'h2)); forvar1611 = (forvar1611 + (1'h1)))
                    begin
                      reg1612 <= forvar1598[(4'ha):(2'h3)];
                    end
                  for (forvar1613 = (1'h0); (forvar1613 < (1'h1)); forvar1613 = (forvar1613 + (1'h1)))
                    begin
                      reg1614 <= (~|$unsigned(forvar1613));
                      reg1615 <= reg1599[(3'h4):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar1605 = (1'h0); (forvar1605 < (2'h3)); forvar1605 = (forvar1605 + (1'h1)))
                    begin
                      reg1606 <= forvar1569;
                      reg1607 <= $unsigned((reg1608[(3'h6):(1'h0)] <= (!(^(8'haa)))));
                    end
                end
              reg1616 <= ((~|forvar1605[(3'h5):(2'h2)]) - $unsigned((+(wire1546 << forvar1557))));
            end
          for (forvar1617 = (1'h0); (forvar1617 < (1'h0)); forvar1617 = (forvar1617 + (1'h1)))
            begin
              for (forvar1618 = (1'h0); (forvar1618 < (2'h2)); forvar1618 = (forvar1618 + (1'h1)))
                begin
                  for (forvar1619 = (1'h0); (forvar1619 < (2'h2)); forvar1619 = (forvar1619 + (1'h1)))
                    begin
                      reg1620 <= {$unsigned((^(|reg1575)))};
                      reg1621 <= $signed($signed(wire1547[(2'h2):(1'h1)]));
                    end
                  for (forvar1622 = (1'h0); (forvar1622 < (1'h1)); forvar1622 = (forvar1622 + (1'h1)))
                    begin
                      reg1623 <= $signed(((^~$signed(reg1602)) ?
                          {reg1584} : (|wire1546)));
                      reg1624 <= reg1582[(3'h7):(3'h4)];
                      reg1625 <= $unsigned((forvar1559 > $unsigned($unsigned(forvar1564))));
                      reg1626 <= reg1598;
                    end
                end
              for (forvar1627 = (1'h0); (forvar1627 < (1'h0)); forvar1627 = (forvar1627 + (1'h1)))
                begin
                  reg1628 <= $unsigned($signed($signed($unsigned(forvar1617))));
                end
              if (reg1582[(1'h0):(1'h0)])
                begin
                  for (forvar1629 = (1'h0); (forvar1629 < (2'h2)); forvar1629 = (forvar1629 + (1'h1)))
                    begin
                      reg1630 <= (!(reg1592 <= reg1589));
                      reg1631 <= ({($unsigned(reg1599) >= (forvar1598 ?
                              reg1623 : (8'h9d)))} != ($signed($signed((8'hb2))) != {(^forvar1618)}));
                      reg1632 <= $signed(reg1590[(3'h4):(3'h4)]);
                    end
                  for (forvar1633 = (1'h0); (forvar1633 < (1'h0)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= (&reg1555[(2'h3):(1'h1)]);
                      reg1635 <= reg1616;
                    end
                  reg1636 <= reg1584;
                end
              else
                begin
                  for (forvar1629 = (1'h0); (forvar1629 < (2'h3)); forvar1629 = (forvar1629 + (1'h1)))
                    begin
                      reg1630 <= ($signed(reg1608[(4'h8):(4'h8)]) ?
                          (forvar1604 ?
                              reg1621 : $signed(reg1636[(2'h3):(1'h1)])) : (((reg1582 ?
                              forvar1590 : reg1563) >= reg1572) <<< ($signed(reg1550) ?
                              reg1635[(3'h6):(3'h5)] : $unsigned(reg1625))));
                      reg1631 <= ({{(wire1542 ?
                                  reg1570 : (8'ha6))}} || ((reg1561[(3'h5):(3'h5)] < reg1566) >>> $signed(reg1563[(2'h3):(2'h2)])));
                      reg1632 <= (^~((reg1587 - (~|reg1626)) != $signed($unsigned(reg1616))));
                      reg1633 <= $signed(forvar1611[(2'h2):(2'h2)]);
                    end
                  reg1634 <= (-(reg1602 ?
                      (!(~^(8'ha8))) : (+(reg1612 ~^ reg1570))));
                end
            end
          for (forvar1637 = (1'h0); (forvar1637 < (1'h0)); forvar1637 = (forvar1637 + (1'h1)))
            begin
              if ($unsigned(forvar1589[(3'h5):(1'h1)]))
                begin
                  for (forvar1638 = (1'h0); (forvar1638 < (1'h1)); forvar1638 = (forvar1638 + (1'h1)))
                    begin
                      reg1639 <= $unsigned($unsigned((8'hab)));
                      reg1640 <= ((forvar1556 ?
                          ((&forvar1550) << reg1561[(4'ha):(3'h7)]) : {$signed((8'hb7))}) >>> (~(reg1570 & (reg1571 && reg1551))));
                    end
                  for (forvar1641 = (1'h0); (forvar1641 < (1'h1)); forvar1641 = (forvar1641 + (1'h1)))
                    begin
                      reg1642 <= (($unsigned((~&(8'hae))) && $unsigned($unsigned((8'h9c)))) ^ reg1582);
                      reg1643 <= $unsigned(reg1626);
                    end
                  if (((-wire1544[(2'h2):(1'h0)]) ?
                      ((-$unsigned(reg1566)) ?
                          $unsigned((reg1557 ? reg1572 : reg1614)) : {(reg1607 ?
                                  reg1628 : reg1581)}) : ($unsigned({reg1579}) >> forvar1604)))
                    begin
                      reg1644 <= $signed(reg1602[(2'h3):(2'h2)]);
                      reg1645 <= (^~{$unsigned((~&forvar1605))});
                      reg1646 <= ((^~$unsigned($signed(reg1644))) * $unsigned(forvar1564[(1'h0):(1'h0)]));
                      reg1647 <= reg1561[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg1644 <= (~forvar1589[(3'h7):(3'h7)]);
                      reg1645 <= ((~&({reg1563} ?
                              forvar1590[(4'h9):(3'h7)] : $signed(reg1597))) ?
                          (($signed(reg1551) > reg1608[(1'h0):(1'h0)]) >> $signed((8'hae))) : (((reg1630 ?
                                  reg1639 : forvar1618) ?
                              $unsigned(reg1595) : (reg1593 ?
                                  reg1582 : (8'ha1))) || $unsigned(((8'hae) | wire1544))));
                      reg1646 <= $signed({$unsigned((&reg1550))});
                    end
                end
              else
                begin
                  for (forvar1638 = (1'h0); (forvar1638 < (2'h2)); forvar1638 = (forvar1638 + (1'h1)))
                    begin
                      reg1639 <= reg1595[(2'h2):(1'h0)];
                    end
                  for (forvar1640 = (1'h0); (forvar1640 < (1'h0)); forvar1640 = (forvar1640 + (1'h1)))
                    begin
                      reg1641 <= reg1574;
                      reg1642 <= reg1574;
                    end
                end
              reg1648 <= $signed({({wire1541} < forvar1548)});
              if ($unsigned({$unsigned(reg1644)}))
                begin
                  if ($unsigned((~^reg1573[(4'hc):(3'h5)])))
                    begin
                      reg1649 <= ({((reg1566 || forvar1559) <<< $unsigned(reg1631))} ?
                          (|$unsigned(wire1542[(2'h3):(2'h3)])) : $unsigned(reg1636));
                      reg1650 <= $signed((reg1610 ^~ (reg1588[(4'hc):(2'h3)] && $signed(reg1582))));
                    end
                  else
                    begin
                      reg1649 <= ((|(reg1609 >>> wire1543)) ?
                          {forvar1560} : (8'hb9));
                      reg1650 <= {reg1566};
                      reg1651 <= $unsigned((reg1634[(1'h0):(1'h0)] ?
                          (8'had) : ((!reg1599) ?
                              ((8'hb7) ?
                                  reg1628 : (8'hb9)) : (forvar1611 * reg1616))));
                    end
                  reg1652 <= (8'h9d);
                end
              else
                begin
                  if ($signed(($signed((~&reg1562)) <= ({(8'h9e)} | (-forvar1556)))))
                    begin
                      reg1649 <= $signed(forvar1578[(4'ha):(2'h2)]);
                    end
                  else
                    begin
                      reg1649 <= ($unsigned(reg1563) ^ (8'ha5));
                      reg1650 <= $signed(reg1586);
                      reg1651 <= forvar1560;
                    end
                end
              for (forvar1653 = (1'h0); (forvar1653 < (1'h0)); forvar1653 = (forvar1653 + (1'h1)))
                begin
                  reg1654 <= ($unsigned((+(forvar1637 ?
                          (8'hb5) : forvar1653))) ?
                      (~((wire1543 > reg1612) != (~^(8'hae)))) : ($unsigned(forvar1578) * $signed(forvar1591[(2'h2):(1'h0)])));
                end
            end
        end
      else
        begin
          for (forvar1604 = (1'h0); (forvar1604 < (2'h2)); forvar1604 = (forvar1604 + (1'h1)))
            begin
              if ({((~^{reg1557}) == $unsigned(((8'hb1) ?
                      reg1654 : forvar1637)))})
                begin
                  for (forvar1605 = (1'h0); (forvar1605 < (1'h1)); forvar1605 = (forvar1605 + (1'h1)))
                    begin
                      reg1606 <= reg1648[(4'h8):(3'h7)];
                      reg1607 <= reg1572;
                    end
                  for (forvar1608 = (1'h0); (forvar1608 < (2'h3)); forvar1608 = (forvar1608 + (1'h1)))
                    begin
                      reg1609 <= forvar1641[(2'h3):(2'h3)];
                      reg1610 <= $unsigned(((!((8'hb8) >= (8'hb0))) * ((reg1612 ^ reg1640) ?
                          (^~reg1612) : ((8'hb0) + reg1591))));
                      reg1611 <= ({reg1590[(3'h5):(2'h2)]} ?
                          {((!reg1553) & reg1600)} : forvar1627[(2'h3):(2'h2)]);
                    end
                  if (({(^(+reg1550))} ?
                      (8'hb0) : (((^~forvar1556) | (forvar1633 ?
                              reg1648 : forvar1611)) ?
                          ((~^reg1641) ?
                              (!reg1607) : (forvar1550 ?
                                  (8'hb9) : forvar1590)) : $signed((~forvar1588)))))
                    begin
                      reg1612 <= (~^(^~({wire1545} > forvar1564)));
                      reg1613 <= (^(~&(~&((8'hb5) ? reg1601 : reg1593))));
                      reg1614 <= ($unsigned((+(~forvar1590))) ~^ wire1547);
                    end
                  else
                    begin
                      reg1612 <= $signed((+(!$unsigned(forvar1559))));
                      reg1613 <= {(^reg1552)};
                    end
                end
              else
                begin
                  for (forvar1605 = (1'h0); (forvar1605 < (1'h1)); forvar1605 = (forvar1605 + (1'h1)))
                    begin
                      reg1606 <= reg1642;
                      reg1607 <= $unsigned(forvar1633[(1'h1):(1'h0)]);
                      reg1608 <= (($unsigned((^~forvar1638)) ?
                              reg1631 : $unsigned({reg1602})) ?
                          {$unsigned((+wire1542))} : (~{{forvar1594}}));
                      reg1609 <= (reg1592 > (-forvar1633));
                    end
                  for (forvar1610 = (1'h0); (forvar1610 < (1'h0)); forvar1610 = (forvar1610 + (1'h1)))
                    begin
                      reg1611 <= $unsigned((-(~|reg1646[(4'hb):(2'h2)])));
                    end
                end
              if ($unsigned($unsigned(reg1576)))
                begin
                  reg1615 <= (&$signed(({reg1585} >= $signed(reg1647))));
                end
              else
                begin
                  if ($unsigned(forvar1610[(1'h1):(1'h0)]))
                    begin
                      reg1615 <= $signed((~^$signed({(8'hb5)})));
                    end
                  else
                    begin
                      reg1615 <= (!reg1556[(2'h2):(2'h2)]);
                      reg1616 <= (|$signed($unsigned((reg1601 <<< reg1635))));
                      reg1617 <= $signed((forvar1611[(1'h0):(1'h0)] | (~&(reg1635 ?
                          reg1551 : reg1577))));
                    end
                  for (forvar1618 = (1'h0); (forvar1618 < (1'h1)); forvar1618 = (forvar1618 + (1'h1)))
                    begin
                      reg1619 <= forvar1610;
                      reg1620 <= $signed(forvar1588);
                    end
                  if ((forvar1629[(2'h2):(1'h0)] ?
                      (8'hab) : reg1582[(4'ha):(3'h5)]))
                    begin
                      reg1621 <= reg1580;
                      reg1622 <= $unsigned(forvar1569[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg1621 <= $signed(forvar1640[(1'h0):(1'h0)]);
                    end
                  for (forvar1623 = (1'h0); (forvar1623 < (1'h1)); forvar1623 = (forvar1623 + (1'h1)))
                    begin
                      reg1624 <= (forvar1590 - (!$unsigned((reg1647 ^~ forvar1629))));
                      reg1625 <= reg1599;
                      reg1626 <= $unsigned(((^~$signed(reg1587)) ?
                          forvar1638[(3'h7):(1'h1)] : $unsigned($signed(reg1648))));
                      reg1627 <= $signed($signed(reg1586));
                    end
                end
              if (forvar1550)
                begin
                  for (forvar1628 = (1'h0); (forvar1628 < (1'h1)); forvar1628 = (forvar1628 + (1'h1)))
                    begin
                      reg1629 <= forvar1653;
                      reg1630 <= $unsigned($unsigned({(reg1558 ?
                              reg1579 : forvar1622)}));
                    end
                  if (reg1584)
                    begin
                      reg1631 <= ((8'hb9) | reg1654);
                      reg1632 <= ((~^({reg1582} ?
                          forvar1619[(2'h3):(2'h2)] : $unsigned(reg1577))) * $signed(($unsigned(forvar1578) ?
                          reg1586[(4'hb):(1'h1)] : $unsigned((8'ha8)))));
                      reg1633 <= (($signed(reg1598[(4'ha):(1'h0)]) ?
                              reg1594 : {reg1614[(3'h5):(2'h3)]}) ?
                          $signed($signed({reg1609})) : wire1546[(3'h5):(2'h2)]);
                    end
                  else
                    begin
                      reg1631 <= $signed(((forvar1618 >>> $unsigned((8'hb3))) ?
                          (~$signed(forvar1556)) : reg1600[(2'h2):(1'h0)]));
                      reg1632 <= reg1615;
                      reg1633 <= reg1603;
                    end
                end
              else
                begin
                  reg1628 <= (^~({reg1617} < $unsigned({reg1583})));
                  if ((reg1611 << reg1582))
                    begin
                      reg1629 <= (reg1581[(4'h8):(3'h5)] ?
                          (((~^forvar1591) <= $unsigned(forvar1641)) ?
                              reg1644 : {(reg1608 - reg1642)}) : $unsigned($signed(forvar1627[(2'h2):(1'h1)])));
                      reg1630 <= reg1610[(4'he):(4'hb)];
                      reg1631 <= $unsigned(forvar1569[(2'h2):(1'h1)]);
                      reg1632 <= reg1567;
                    end
                  else
                    begin
                      reg1629 <= $unsigned(($signed((reg1631 ?
                          reg1570 : reg1583)) >= (reg1639[(4'ha):(4'ha)] || $signed(reg1580))));
                      reg1630 <= $signed(((-(~^wire1547)) >> (reg1573[(4'ha):(4'h8)] >>> forvar1637)));
                      reg1631 <= $signed(forvar1564[(1'h0):(1'h0)]);
                      reg1632 <= ($signed($unsigned($unsigned(reg1626))) != $unsigned(reg1558));
                    end
                  if ((|$unsigned(reg1626[(2'h3):(2'h2)])))
                    begin
                      reg1633 <= forvar1618;
                      reg1634 <= (($signed((forvar1550 ?
                              reg1576 : forvar1637)) ?
                          reg1652 : ((reg1647 ?
                              (8'ha6) : reg1576) >>> {reg1625})) >>> $unsigned(reg1652[(3'h4):(3'h4)]));
                      reg1635 <= {($unsigned({reg1639}) ?
                              reg1583 : ($signed(reg1646) ?
                                  $unsigned(forvar1641) : $unsigned(forvar1578)))};
                      reg1636 <= (reg1643 ?
                          reg1644 : (&(~$signed(forvar1589))));
                    end
                  else
                    begin
                      reg1633 <= forvar1638;
                      reg1634 <= $unsigned($signed(($unsigned(reg1616) - $unsigned(reg1607))));
                    end
                end
              for (forvar1637 = (1'h0); (forvar1637 < (1'h1)); forvar1637 = (forvar1637 + (1'h1)))
                begin
                  for (forvar1638 = (1'h0); (forvar1638 < (1'h1)); forvar1638 = (forvar1638 + (1'h1)))
                    begin
                      reg1639 <= $signed(((!reg1606[(4'hb):(3'h4)]) ?
                          ($unsigned(reg1587) << forvar1578) : (reg1652[(1'h0):(1'h0)] ^ $unsigned(reg1586))));
                      reg1640 <= forvar1564;
                      reg1641 <= (reg1597 ?
                          ($unsigned((!reg1612)) ^ reg1571[(4'h8):(2'h3)]) : $signed(((reg1549 & forvar1653) | (forvar1611 ?
                              forvar1548 : reg1646))));
                      reg1642 <= reg1610;
                    end
                  for (forvar1643 = (1'h0); (forvar1643 < (1'h1)); forvar1643 = (forvar1643 + (1'h1)))
                    begin
                      reg1644 <= forvar1598;
                      reg1645 <= $signed({(reg1630 ?
                              $signed(reg1571) : {reg1654})});
                      reg1646 <= (~($signed($signed(reg1608)) <= ({forvar1629} ?
                          (~|forvar1613) : $unsigned(forvar1611))));
                      reg1647 <= forvar1613[(1'h0):(1'h0)];
                    end
                  if ({forvar1590[(2'h3):(1'h0)]})
                    begin
                      reg1648 <= $unsigned(reg1612[(1'h1):(1'h0)]);
                      reg1649 <= wire1544[(2'h3):(1'h0)];
                      reg1650 <= (reg1609 >= ((8'haa) >> forvar1640[(3'h4):(1'h1)]));
                    end
                  else
                    begin
                      reg1648 <= $unsigned((reg1652 ^~ $unsigned({reg1624})));
                      reg1649 <= $signed((~^((~^reg1581) * reg1594)));
                      reg1650 <= reg1648;
                      reg1651 <= reg1567[(4'ha):(3'h6)];
                    end
                  if ($unsigned($signed((!(forvar1611 == forvar1619)))))
                    begin
                      reg1652 <= reg1585[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1652 <= forvar1613;
                      reg1653 <= ((8'hb2) ?
                          reg1635[(4'ha):(4'ha)] : ($unsigned((reg1645 ?
                                  reg1635 : (8'hb9))) ?
                              reg1576 : ($unsigned(reg1646) ?
                                  reg1599 : ((8'ha9) ? (8'ha0) : (8'haa)))));
                      reg1654 <= $unsigned($signed((+(^forvar1585))));
                    end
                end
            end
          for (forvar1655 = (1'h0); (forvar1655 < (2'h2)); forvar1655 = (forvar1655 + (1'h1)))
            begin
              if (({(8'ha7)} ?
                  ($unsigned(reg1610) ?
                      (8'ha6) : {$signed(reg1628)}) : {$signed((~reg1555))}))
                begin
                  for (forvar1656 = (1'h0); (forvar1656 < (2'h3)); forvar1656 = (forvar1656 + (1'h1)))
                    begin
                      reg1657 <= $signed($unsigned($unsigned((&forvar1569))));
                      reg1658 <= (reg1657 >= (~{(reg1613 || reg1649)}));
                      reg1659 <= (reg1645[(4'h8):(4'h8)] | forvar1656[(4'ha):(2'h3)]);
                    end
                end
              else
                begin
                  for (forvar1656 = (1'h0); (forvar1656 < (2'h3)); forvar1656 = (forvar1656 + (1'h1)))
                    begin
                      reg1657 <= reg1558[(4'h9):(2'h2)];
                      reg1658 <= (reg1621[(3'h7):(3'h7)] << $unsigned($signed((reg1551 ?
                          reg1580 : reg1623))));
                    end
                end
              for (forvar1660 = (1'h0); (forvar1660 < (1'h1)); forvar1660 = (forvar1660 + (1'h1)))
                begin
                  if ((reg1648 >>> reg1570))
                    begin
                      reg1661 <= (^~reg1611[(3'h6):(1'h0)]);
                    end
                  else
                    begin
                      reg1661 <= $signed(((reg1639 || forvar1598[(1'h1):(1'h1)]) && (8'hae)));
                      reg1662 <= (~(^((^~(8'ha7)) ?
                          forvar1604[(4'hc):(1'h0)] : {forvar1629})));
                      reg1663 <= $unsigned(($unsigned({forvar1591}) ^~ forvar1589[(3'h5):(3'h4)]));
                      reg1664 <= reg1654;
                    end
                  reg1665 <= ($signed(reg1592[(2'h3):(2'h3)]) ?
                      (reg1580 ^~ $signed((~forvar1608))) : (~^reg1610));
                end
              for (forvar1666 = (1'h0); (forvar1666 < (1'h1)); forvar1666 = (forvar1666 + (1'h1)))
                begin
                  reg1667 <= (8'ha4);
                  if (($signed((~^reg1625)) | (($unsigned(reg1553) - $signed(reg1599)) != (((8'hb8) && reg1635) <= reg1663))))
                    begin
                      reg1668 <= reg1620[(2'h2):(1'h0)];
                      reg1669 <= reg1602;
                      reg1670 <= reg1549;
                      reg1671 <= ($unsigned(((forvar1594 * reg1581) < $unsigned(reg1566))) ?
                          $signed(forvar1559) : forvar1557[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg1668 <= forvar1548;
                      reg1669 <= (reg1627[(3'h4):(2'h3)] ?
                          (&(-$unsigned((8'hb0)))) : forvar1549);
                      reg1670 <= reg1641[(2'h2):(1'h1)];
                      reg1671 <= $signed((8'hb5));
                    end
                  for (forvar1672 = (1'h0); (forvar1672 < (2'h2)); forvar1672 = (forvar1672 + (1'h1)))
                    begin
                      reg1673 <= reg1601;
                      reg1674 <= ($signed(reg1609) <<< (!$signed($unsigned(reg1615))));
                      reg1675 <= $signed((reg1667[(2'h2):(2'h2)] == reg1591[(4'h8):(3'h4)]));
                    end
                end
            end
        end
      for (forvar1676 = (1'h0); (forvar1676 < (2'h3)); forvar1676 = (forvar1676 + (1'h1)))
        begin
          for (forvar1677 = (1'h0); (forvar1677 < (1'h0)); forvar1677 = (forvar1677 + (1'h1)))
            begin
              if (forvar1672[(4'h8):(3'h5)])
                begin
                  for (forvar1678 = (1'h0); (forvar1678 < (1'h1)); forvar1678 = (forvar1678 + (1'h1)))
                    begin
                      reg1679 <= reg1563;
                    end
                  for (forvar1680 = (1'h0); (forvar1680 < (1'h0)); forvar1680 = (forvar1680 + (1'h1)))
                    begin
                      reg1681 <= $unsigned($unsigned((|(reg1651 ?
                          reg1595 : reg1552))));
                      reg1682 <= forvar1590[(4'hc):(2'h3)];
                      reg1683 <= (~^reg1584[(4'hb):(3'h5)]);
                    end
                  for (forvar1684 = (1'h0); (forvar1684 < (1'h0)); forvar1684 = (forvar1684 + (1'h1)))
                    begin
                      reg1685 <= (({forvar1556[(3'h5):(1'h0)]} ?
                              (^(~reg1663)) : ((reg1590 << forvar1643) ?
                                  $signed(forvar1560) : (reg1651 ?
                                      reg1679 : forvar1585))) ?
                          $unsigned($signed(reg1609)) : (+(reg1601 <= forvar1656)));
                      reg1686 <= reg1659;
                    end
                  for (forvar1687 = (1'h0); (forvar1687 < (1'h1)); forvar1687 = (forvar1687 + (1'h1)))
                    begin
                      reg1688 <= (-($signed($signed(forvar1672)) >= ((^~reg1659) ?
                          (~&reg1623) : $unsigned(forvar1618))));
                      reg1689 <= ($signed($unsigned($signed(reg1602))) || forvar1565);
                      reg1690 <= $unsigned($unsigned((~forvar1641[(4'he):(1'h0)])));
                      reg1691 <= reg1619[(3'h4):(3'h4)];
                    end
                end
              else
                begin
                  reg1678 <= forvar1564;
                  for (forvar1679 = (1'h0); (forvar1679 < (1'h1)); forvar1679 = (forvar1679 + (1'h1)))
                    begin
                      reg1680 <= (~&forvar1588);
                      reg1681 <= (~reg1634);
                      reg1682 <= (($signed((^~forvar1559)) ?
                          (reg1689 != reg1580[(4'hb):(3'h7)]) : ((reg1617 ?
                              reg1623 : reg1679) == $signed(reg1576))) ^~ $unsigned($signed($signed(reg1561))));
                      reg1683 <= (reg1577[(2'h3):(2'h2)] ?
                          {reg1581} : $signed({(~|reg1556)}));
                    end
                end
            end
        end
      for (forvar1692 = (1'h0); (forvar1692 < (1'h1)); forvar1692 = (forvar1692 + (1'h1)))
        begin
          if ($unsigned($unsigned($signed($signed((8'hac))))))
            begin
              reg1693 <= $unsigned({((reg1644 & reg1587) ?
                      $unsigned(reg1674) : $unsigned((8'ha7)))});
              if ({(reg1603 ?
                      ((reg1582 ? forvar1633 : (8'ha0)) ?
                          {(8'ha4)} : forvar1679[(3'h6):(3'h4)]) : {$signed(reg1617)})})
                begin
                  if (($unsigned($signed((~^forvar1622))) ?
                      $unsigned(($signed((8'hb6)) ?
                          (8'ha7) : (~|forvar1578))) : (8'ha9)))
                    begin
                      reg1694 <= $signed((reg1556 >>> $signed((reg1554 > (8'hb8)))));
                      reg1695 <= wire1546;
                    end
                  else
                    begin
                      reg1694 <= (-{($signed(reg1575) ^~ (reg1598 == forvar1638))});
                      reg1695 <= reg1562;
                      reg1696 <= reg1667[(4'h8):(1'h1)];
                    end
                  for (forvar1697 = (1'h0); (forvar1697 < (1'h0)); forvar1697 = (forvar1697 + (1'h1)))
                    begin
                      reg1698 <= (!reg1587[(3'h7):(1'h1)]);
                      reg1699 <= {(reg1583 && reg1585)};
                      reg1700 <= ((~|((&reg1622) ?
                          $unsigned(reg1597) : ((8'hb9) ?
                              reg1650 : forvar1613))) | (~&(&$signed(reg1633))));
                    end
                end
              else
                begin
                  for (forvar1694 = (1'h0); (forvar1694 < (1'h0)); forvar1694 = (forvar1694 + (1'h1)))
                    begin
                      reg1695 <= ((~^$unsigned(reg1671)) ?
                          $signed(({reg1607} ?
                              forvar1623 : (|(8'hb4)))) : $signed(forvar1585));
                    end
                end
              if ($signed(reg1576))
                begin
                  for (forvar1701 = (1'h0); (forvar1701 < (2'h2)); forvar1701 = (forvar1701 + (1'h1)))
                    begin
                      reg1702 <= $signed((^~(wire1545[(3'h6):(1'h0)] - (~^reg1654))));
                      reg1703 <= (8'hb7);
                      reg1704 <= ($unsigned($unsigned($unsigned((8'hae)))) ?
                          {forvar1588} : $unsigned((~&{reg1662})));
                    end
                  if (((~$signed({reg1570})) ?
                      ($signed({wire1544}) >>> $unsigned({reg1587})) : (-(^(wire1542 < reg1680)))))
                    begin
                      reg1705 <= (~({{reg1699}} != (~^(8'h9d))));
                      reg1706 <= $signed((~|$unsigned({reg1640})));
                      reg1707 <= (|forvar1619[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1705 <= ($signed({forvar1637[(4'ha):(3'h7)]}) & {(~&$signed(reg1556))});
                    end
                  for (forvar1708 = (1'h0); (forvar1708 < (1'h0)); forvar1708 = (forvar1708 + (1'h1)))
                    begin
                      reg1709 <= $signed((|$unsigned(reg1619)));
                      reg1710 <= reg1695[(4'he):(4'ha)];
                    end
                end
              else
                begin
                  if (reg1665)
                    begin
                      reg1701 <= {$unsigned(reg1645[(3'h7):(2'h2)])};
                      reg1702 <= ((|{(reg1624 ?
                              (8'hb6) : (8'ha7))}) | (~|(8'hb7)));
                      reg1703 <= $signed((8'had));
                    end
                  else
                    begin
                      reg1701 <= $unsigned(forvar1564);
                      reg1702 <= ($signed({(~|forvar1672)}) ?
                          ((8'h9d) || ((8'haa) ^~ reg1688[(2'h3):(1'h0)])) : reg1698[(4'hd):(2'h3)]);
                      reg1703 <= forvar1560;
                    end
                  if ($unsigned($unsigned($signed(((8'hb1) >= forvar1622)))))
                    begin
                      reg1704 <= reg1651;
                      reg1705 <= (($unsigned($signed((8'hb6))) <<< reg1555) ?
                          (reg1681 >>> $signed($unsigned(reg1603))) : ({(reg1678 && reg1593)} + $unsigned((reg1682 ?
                              forvar1708 : (8'hb1)))));
                      reg1706 <= $signed((&reg1611));
                      reg1707 <= reg1596;
                    end
                  else
                    begin
                      reg1704 <= ($unsigned(((&(8'ha7)) <= reg1651[(2'h2):(2'h2)])) << reg1587[(3'h7):(3'h4)]);
                      reg1705 <= (($unsigned(reg1593[(2'h2):(1'h1)]) ?
                              reg1640[(2'h2):(2'h2)] : (8'hb5)) ?
                          $unsigned($signed($unsigned((8'ha5)))) : {($signed((8'ha7)) ?
                                  ((8'h9f) ^~ reg1580) : (reg1675 ?
                                      reg1673 : (8'hb6)))});
                      reg1706 <= reg1580;
                      reg1707 <= (^(^{$unsigned(forvar1610)}));
                    end
                  for (forvar1708 = (1'h0); (forvar1708 < (2'h3)); forvar1708 = (forvar1708 + (1'h1)))
                    begin
                      reg1709 <= (($unsigned((8'h9f)) ?
                          reg1583 : ($unsigned(reg1617) + {(8'ha0)})) >> $unsigned((forvar1590[(3'h7):(2'h3)] ?
                          (reg1696 ? forvar1641 : reg1550) : forvar1585)));
                      reg1710 <= reg1688[(1'h0):(1'h0)];
                      reg1711 <= $unsigned((({forvar1611} ?
                              (&forvar1694) : reg1586[(4'hd):(3'h5)]) ?
                          $signed($unsigned(forvar1655)) : ((reg1576 ?
                                  forvar1627 : reg1568) ?
                              forvar1622 : {reg1690})));
                      reg1712 <= (+forvar1594);
                    end
                  if (forvar1655[(4'h8):(2'h2)])
                    begin
                      reg1713 <= reg1619[(2'h3):(1'h0)];
                      reg1714 <= $signed((8'hac));
                    end
                  else
                    begin
                      reg1713 <= $unsigned(reg1667);
                    end
                end
            end
          else
            begin
              reg1693 <= $unsigned((((reg1615 == reg1685) << (forvar1677 && reg1674)) ?
                  reg1703 : $signed((~&reg1663))));
            end
          if ($signed((+(reg1631 | forvar1619[(1'h1):(1'h0)]))))
            begin
              for (forvar1715 = (1'h0); (forvar1715 < (1'h0)); forvar1715 = (forvar1715 + (1'h1)))
                begin
                  for (forvar1716 = (1'h0); (forvar1716 < (1'h0)); forvar1716 = (forvar1716 + (1'h1)))
                    begin
                      reg1717 <= {$signed((&forvar1638))};
                    end
                end
              if ((-(&(8'hb1))))
                begin
                  reg1718 <= $signed((reg1631[(2'h3):(2'h2)] ?
                      forvar1613 : (~^$signed(reg1675))));
                  reg1719 <= ($unsigned({(reg1700 + (8'hb2))}) ?
                      reg1598 : (8'ha9));
                  if ({$signed($unsigned($unsigned(forvar1708)))})
                    begin
                      reg1720 <= forvar1605;
                    end
                  else
                    begin
                      reg1720 <= ({((|reg1590) ?
                                  forvar1643 : $signed((8'haf)))} ?
                          reg1599 : $unsigned(({forvar1660} ?
                              ((8'ha7) != reg1639) : reg1663)));
                    end
                end
              else
                begin
                  if ((|(~&$signed((&(8'ha6))))))
                    begin
                      reg1718 <= $signed(forvar1564[(3'h6):(2'h2)]);
                      reg1719 <= forvar1677;
                      reg1720 <= reg1658;
                    end
                  else
                    begin
                      reg1718 <= reg1597;
                      reg1719 <= (reg1591[(2'h2):(1'h0)] ^ (-$signed($signed((8'had)))));
                      reg1720 <= reg1643;
                    end
                end
              if (($signed($signed($unsigned(reg1641))) << ({((8'ha0) ?
                          (8'hac) : reg1661)} ?
                  $unsigned($signed(forvar1680)) : $signed(reg1688[(2'h2):(1'h0)]))))
                begin
                  for (forvar1721 = (1'h0); (forvar1721 < (1'h0)); forvar1721 = (forvar1721 + (1'h1)))
                    begin
                      reg1722 <= ({reg1590[(3'h5):(3'h5)]} != $unsigned($unsigned({reg1567})));
                    end
                end
              else
                begin
                  for (forvar1721 = (1'h0); (forvar1721 < (2'h3)); forvar1721 = (forvar1721 + (1'h1)))
                    begin
                      reg1722 <= ($unsigned(($unsigned(reg1563) ?
                          ((8'ha5) ? reg1595 : reg1589) : (reg1688 ?
                              reg1608 : reg1549))) ^ reg1671[(3'h7):(1'h0)]);
                    end
                  for (forvar1723 = (1'h0); (forvar1723 < (1'h1)); forvar1723 = (forvar1723 + (1'h1)))
                    begin
                      reg1724 <= (|reg1571);
                    end
                  reg1725 <= (forvar1629 ?
                      forvar1697 : ((&(~reg1626)) >>> $signed($unsigned((8'hb2)))));
                end
            end
          else
            begin
              for (forvar1715 = (1'h0); (forvar1715 < (1'h1)); forvar1715 = (forvar1715 + (1'h1)))
                begin
                  reg1716 <= ($unsigned(((|reg1558) < $unsigned(forvar1676))) ?
                      ($unsigned(reg1600[(1'h1):(1'h0)]) ?
                          $unsigned((!reg1682)) : $signed($unsigned(reg1597))) : $signed((+(wire1545 ~^ reg1717))));
                  if (reg1649[(3'h5):(3'h4)])
                    begin
                      reg1717 <= $unsigned($unsigned((8'hba)));
                      reg1718 <= (!reg1659);
                    end
                  else
                    begin
                      reg1717 <= $unsigned((~&$unsigned(((8'ha5) ?
                          forvar1666 : reg1592))));
                    end
                  for (forvar1719 = (1'h0); (forvar1719 < (1'h1)); forvar1719 = (forvar1719 + (1'h1)))
                    begin
                      reg1720 <= {(8'ha0)};
                      reg1721 <= $unsigned((~|(^~$unsigned(reg1669))));
                    end
                end
            end
          for (forvar1726 = (1'h0); (forvar1726 < (2'h3)); forvar1726 = (forvar1726 + (1'h1)))
            begin
              if (({(forvar1692 < $signed(reg1646))} ?
                  (($unsigned(wire1543) ?
                          {reg1681} : (reg1586 ? reg1615 : reg1679)) ?
                      ({reg1582} == (~forvar1618)) : reg1695) : (($unsigned(reg1558) ?
                          (reg1612 ?
                              reg1719 : reg1563) : forvar1653[(2'h3):(1'h0)]) ?
                      {$unsigned(forvar1588)} : $signed(reg1717))))
                begin
                  reg1727 <= (^$unsigned(((forvar1708 ?
                      reg1639 : forvar1627) <= $signed(forvar1641))));
                  if (($unsigned($signed((|reg1644))) ?
                      forvar1679[(2'h2):(1'h0)] : reg1649))
                    begin
                      reg1728 <= forvar1550[(4'ha):(1'h1)];
                      reg1729 <= {($unsigned((+forvar1578)) ?
                              reg1648 : ($signed(reg1593) ?
                                  (forvar1594 < reg1595) : (&reg1716)))};
                    end
                  else
                    begin
                      reg1728 <= $signed($signed({{forvar1672}}));
                      reg1729 <= forvar1617;
                    end
                end
              else
                begin
                  for (forvar1727 = (1'h0); (forvar1727 < (2'h3)); forvar1727 = (forvar1727 + (1'h1)))
                    begin
                      reg1728 <= reg1555[(3'h4):(1'h1)];
                      reg1729 <= reg1624[(3'h5):(3'h5)];
                    end
                  reg1730 <= (reg1635 ?
                      (+(+$signed(wire1546))) : $signed((~&(~&(8'hb8)))));
                  if ($signed(reg1549))
                    begin
                      reg1731 <= reg1603;
                      reg1732 <= (|$signed($unsigned({reg1710})));
                    end
                  else
                    begin
                      reg1731 <= (({(reg1667 >>> (8'hb7))} ?
                          ((reg1648 ? forvar1727 : reg1596) ?
                              {reg1556} : reg1561[(4'hc):(3'h5)]) : (~$signed(forvar1629))) > (reg1630 << {$signed(forvar1692)}));
                      reg1732 <= forvar1716[(2'h3):(1'h0)];
                      reg1733 <= forvar1727;
                    end
                end
              for (forvar1734 = (1'h0); (forvar1734 < (2'h2)); forvar1734 = (forvar1734 + (1'h1)))
                begin
                  for (forvar1735 = (1'h0); (forvar1735 < (1'h1)); forvar1735 = (forvar1735 + (1'h1)))
                    begin
                      reg1736 <= {$signed($unsigned(((8'ha3) ?
                              forvar1605 : reg1713)))};
                    end
                end
              reg1737 <= ($signed(((forvar1697 > reg1729) | (~^forvar1735))) >> forvar1622);
            end
          if (reg1579[(1'h0):(1'h0)])
            begin
              for (forvar1738 = (1'h0); (forvar1738 < (1'h1)); forvar1738 = (forvar1738 + (1'h1)))
                begin
                  if (($unsigned(($signed(reg1700) ?
                          reg1553[(4'hb):(4'h9)] : (~forvar1719))) ?
                      wire1543[(4'h8):(1'h1)] : ((reg1636[(3'h7):(3'h4)] == (reg1642 & reg1664)) && {reg1647})))
                    begin
                      reg1739 <= reg1732[(1'h1):(1'h0)];
                      reg1740 <= forvar1655;
                    end
                  else
                    begin
                      reg1739 <= $unsigned((reg1615[(4'hc):(1'h1)] - reg1730[(3'h6):(1'h1)]));
                      reg1740 <= ((reg1703[(4'ha):(2'h3)] ?
                          $unsigned($signed(reg1675)) : (~(reg1719 + reg1591))) <<< ($unsigned(reg1624) || $unsigned($signed((8'hb6)))));
                    end
                  for (forvar1741 = (1'h0); (forvar1741 < (1'h1)); forvar1741 = (forvar1741 + (1'h1)))
                    begin
                      reg1742 <= $unsigned($signed((8'hb0)));
                    end
                end
              for (forvar1743 = (1'h0); (forvar1743 < (1'h1)); forvar1743 = (forvar1743 + (1'h1)))
                begin
                  for (forvar1744 = (1'h0); (forvar1744 < (2'h2)); forvar1744 = (forvar1744 + (1'h1)))
                    begin
                      reg1745 <= (8'hae);
                      reg1746 <= (+forvar1622[(1'h1):(1'h0)]);
                      reg1747 <= ($signed($signed($unsigned((8'haa)))) ?
                          reg1602[(2'h3):(2'h3)] : (~^$unsigned(((8'ha8) ?
                              forvar1676 : reg1711))));
                    end
                  for (forvar1748 = (1'h0); (forvar1748 < (2'h2)); forvar1748 = (forvar1748 + (1'h1)))
                    begin
                      reg1749 <= $unsigned($signed((|(~|forvar1680))));
                      reg1750 <= (reg1640[(1'h1):(1'h1)] && ((&(8'h9e)) ?
                          ((reg1587 ? (8'hb5) : reg1584) ?
                              reg1552[(3'h4):(2'h3)] : reg1651) : ((^~reg1563) != (reg1592 || reg1573))));
                    end
                end
              for (forvar1751 = (1'h0); (forvar1751 < (2'h2)); forvar1751 = (forvar1751 + (1'h1)))
                begin
                  for (forvar1752 = (1'h0); (forvar1752 < (2'h3)); forvar1752 = (forvar1752 + (1'h1)))
                    begin
                      reg1753 <= (~|reg1713);
                      reg1754 <= ($signed((forvar1680[(2'h2):(2'h2)] ?
                              (~^(8'hac)) : (-reg1725))) ?
                          (8'hae) : reg1749);
                    end
                  if (forvar1564)
                    begin
                      reg1755 <= (($unsigned($unsigned(reg1601)) ?
                              $unsigned((reg1581 ?
                                  reg1702 : reg1644)) : reg1695[(3'h5):(3'h5)]) ?
                          $signed(forvar1672) : ({(~^reg1615)} ?
                              $signed($unsigned(forvar1677)) : (!forvar1628[(3'h5):(2'h3)])));
                      reg1756 <= reg1582;
                      reg1757 <= $unsigned(forvar1716[(1'h0):(1'h0)]);
                      reg1758 <= $unsigned(((+reg1714) + forvar1640[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1755 <= (wire1545[(2'h2):(1'h1)] ?
                          ({reg1554} ?
                              reg1549[(2'h2):(2'h2)] : reg1722[(2'h2):(1'h1)]) : $unsigned((~|$signed((8'hb5)))));
                      reg1756 <= forvar1751[(4'h9):(1'h1)];
                      reg1757 <= $signed($signed($signed($unsigned(reg1705))));
                    end
                end
            end
          else
            begin
              if ((((reg1705 ? {forvar1618} : forvar1585) ?
                      ((8'ha7) + reg1696[(3'h7):(1'h0)]) : (!(forvar1727 != reg1756))) ?
                  (((reg1649 <= reg1606) ?
                          reg1705[(1'h0):(1'h0)] : $unsigned(reg1678)) ?
                      $unsigned((reg1551 << reg1675)) : (^(reg1640 ?
                          reg1552 : (8'hb2)))) : reg1626[(2'h3):(2'h3)]))
                begin
                  reg1738 <= (~^reg1714[(3'h6):(3'h4)]);
                  if ($unsigned(reg1678[(4'hb):(1'h1)]))
                    begin
                      reg1739 <= $unsigned($unsigned(((forvar1565 && reg1740) ?
                          (forvar1653 >>> forvar1578) : $signed(reg1664))));
                      reg1740 <= (($unsigned({forvar1565}) | forvar1613[(2'h2):(1'h1)]) ?
                          $signed($unsigned((forvar1738 ?
                              (8'ha4) : reg1594))) : {((forvar1687 ?
                                      reg1653 : forvar1748) ?
                                  {forvar1738} : (reg1563 ?
                                      forvar1588 : reg1727))});
                      reg1741 <= {$unsigned($unsigned(reg1664))};
                    end
                  else
                    begin
                      reg1739 <= reg1556[(4'h8):(3'h7)];
                      reg1740 <= $signed(reg1550[(1'h0):(1'h0)]);
                      reg1741 <= ($unsigned(reg1608[(4'hd):(4'ha)]) ?
                          ((~&(reg1709 ? (8'hb1) : reg1717)) ?
                              (~^$signed(reg1594)) : reg1588) : ((~(reg1561 ?
                                  reg1574 : reg1641)) ?
                              $signed((reg1598 ?
                                  reg1701 : reg1685)) : $signed((reg1566 ?
                                  reg1756 : forvar1627))));
                    end
                end
              else
                begin
                  for (forvar1738 = (1'h0); (forvar1738 < (1'h1)); forvar1738 = (forvar1738 + (1'h1)))
                    begin
                      reg1739 <= (forvar1751[(4'h8):(4'h8)] ?
                          reg1693 : $signed(((reg1671 & reg1631) ^~ reg1659)));
                      reg1740 <= (((-(^forvar1618)) <= $unsigned(forvar1672)) & (~^$unsigned((forvar1622 ~^ reg1731))));
                    end
                  for (forvar1741 = (1'h0); (forvar1741 < (2'h3)); forvar1741 = (forvar1741 + (1'h1)))
                    begin
                      reg1742 <= reg1595[(1'h0):(1'h0)];
                      reg1743 <= (!(+$unsigned($unsigned((8'h9d)))));
                      reg1744 <= $unsigned((reg1745[(3'h4):(1'h0)] ?
                          $signed((~|reg1685)) : ((&reg1682) ?
                              (reg1665 <<< forvar1748) : reg1651)));
                    end
                  for (forvar1745 = (1'h0); (forvar1745 < (2'h3)); forvar1745 = (forvar1745 + (1'h1)))
                    begin
                      reg1746 <= forvar1617;
                      reg1747 <= ({($signed(reg1727) <<< (~&forvar1708))} - $signed($signed(forvar1752)));
                    end
                end
              for (forvar1748 = (1'h0); (forvar1748 < (1'h1)); forvar1748 = (forvar1748 + (1'h1)))
                begin
                  if (({(~^reg1572[(5'h10):(3'h4)])} < {$unsigned(forvar1623[(3'h4):(2'h2)])}))
                    begin
                      reg1749 <= ((reg1754 ?
                              $unsigned((forvar1643 ?
                                  wire1547 : forvar1627)) : $signed($unsigned(reg1625))) ?
                          forvar1619[(2'h3):(1'h0)] : ($signed({reg1703}) << $unsigned((forvar1697 ?
                              forvar1641 : wire1541))));
                      reg1750 <= (&reg1657);
                      reg1751 <= $unsigned((((~|reg1690) < (reg1551 || forvar1679)) ?
                          (reg1720[(4'h8):(3'h6)] ?
                              (reg1671 ?
                                  reg1728 : reg1581) : (+(8'hb8))) : $unsigned((^~reg1661))));
                    end
                  else
                    begin
                      reg1749 <= (reg1688[(3'h4):(3'h4)] >> reg1673);
                      reg1750 <= (8'hba);
                    end
                  if ((($unsigned($signed(forvar1627)) + {forvar1557[(2'h2):(1'h1)]}) | forvar1687))
                    begin
                      reg1752 <= reg1675[(3'h4):(1'h1)];
                      reg1753 <= ($unsigned(((reg1639 ?
                          (8'hb5) : (8'ha8)) <<< $signed(reg1585))) >> reg1724[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg1752 <= (forvar1598 ?
                          (!forvar1640) : reg1568[(4'h9):(4'h9)]);
                    end
                end
              for (forvar1754 = (1'h0); (forvar1754 < (2'h3)); forvar1754 = (forvar1754 + (1'h1)))
                begin
                  reg1755 <= (|$signed(reg1709[(4'hc):(4'hc)]));
                  for (forvar1756 = (1'h0); (forvar1756 < (1'h0)); forvar1756 = (forvar1756 + (1'h1)))
                    begin
                      reg1757 <= (forvar1727 && reg1629[(4'hd):(4'ha)]);
                      reg1758 <= forvar1716[(2'h3):(2'h2)];
                      reg1759 <= (8'haa);
                    end
                  for (forvar1760 = (1'h0); (forvar1760 < (2'h2)); forvar1760 = (forvar1760 + (1'h1)))
                    begin
                      reg1761 <= ({(reg1758 << wire1547)} ?
                          {reg1592} : $unsigned(forvar1550[(4'h8):(3'h6)]));
                      reg1762 <= forvar1613[(2'h3):(1'h1)];
                      reg1763 <= reg1589[(2'h3):(1'h0)];
                    end
                  reg1764 <= (~^$unsigned($signed(reg1698)));
                end
              for (forvar1765 = (1'h0); (forvar1765 < (2'h2)); forvar1765 = (forvar1765 + (1'h1)))
                begin
                  if ((~(reg1571 ?
                      ($signed(reg1706) || reg1630[(3'h4):(1'h1)]) : $unsigned((reg1745 - reg1614)))))
                    begin
                      reg1766 <= $unsigned($unsigned($unsigned(reg1711)));
                      reg1767 <= ($unsigned($unsigned((reg1577 >= (8'hb0)))) << $unsigned(($unsigned(reg1644) ^ (forvar1608 ?
                          reg1594 : reg1679))));
                      reg1768 <= (reg1730 ?
                          forvar1672[(4'hc):(4'h8)] : reg1610);
                    end
                  else
                    begin
                      reg1766 <= (|forvar1617);
                      reg1767 <= reg1588[(1'h1):(1'h0)];
                      reg1768 <= reg1588;
                      reg1769 <= $signed($unsigned(forvar1745));
                    end
                end
            end
        end
    end
  assign wire1770 = $unsigned(reg1752);
  assign wire1771 = ({reg1606} >>> {$unsigned((~|reg1670))});
  always
    @(posedge clk) begin
      if ((({((8'hba) ?
              reg1642 : reg1698)} * $unsigned((+reg1744))) != (reg1568[(4'h9):(3'h6)] ~^ $unsigned($unsigned(reg1630)))))
        begin
          for (forvar1772 = (1'h0); (forvar1772 < (2'h3)); forvar1772 = (forvar1772 + (1'h1)))
            begin
              if ($signed((8'hb3)))
                begin
                  for (forvar1773 = (1'h0); (forvar1773 < (2'h3)); forvar1773 = (forvar1773 + (1'h1)))
                    begin
                      reg1774 <= {$signed(((8'ha8) ?
                              (reg1552 != reg1552) : reg1651[(1'h1):(1'h1)]))};
                      reg1775 <= (^~$signed(reg1769[(1'h0):(1'h0)]));
                      reg1776 <= {$unsigned(forvar1772)};
                      reg1777 <= $unsigned(({$signed(reg1611)} ?
                          ((8'had) ?
                              $signed(reg1738) : $unsigned(reg1576)) : ((reg1718 >= reg1746) + $signed(reg1718))));
                    end
                end
              else
                begin
                  if (reg1639)
                    begin
                      reg1773 <= reg1682[(1'h1):(1'h0)];
                      reg1774 <= (-reg1642);
                      reg1775 <= ($unsigned((reg1640 != (reg1646 ?
                              reg1688 : (8'hb7)))) ?
                          reg1745[(2'h3):(2'h2)] : (8'ha7));
                      reg1776 <= $signed(($signed((^~(8'haf))) << (~|$signed((8'hb2)))));
                    end
                  else
                    begin
                      reg1773 <= (^~(~($signed(reg1661) + (~^reg1733))));
                      reg1774 <= $unsigned($unsigned(((|reg1761) ?
                          (~&reg1630) : reg1567)));
                      reg1775 <= $unsigned((-reg1607[(4'h8):(3'h7)]));
                      reg1776 <= $signed(((&reg1642) != (~&reg1590)));
                    end
                  reg1777 <= (~|(^reg1707[(3'h6):(1'h1)]));
                  for (forvar1778 = (1'h0); (forvar1778 < (2'h3)); forvar1778 = (forvar1778 + (1'h1)))
                    begin
                      reg1779 <= {reg1711};
                      reg1780 <= ($signed((~reg1742[(2'h3):(2'h3)])) ?
                          ((reg1747 == (reg1602 ? reg1707 : reg1600)) ?
                              ($unsigned(reg1762) >> (+reg1570)) : reg1586[(4'hc):(4'h9)]) : $signed(($signed(reg1758) <<< reg1625)));
                    end
                  if (reg1698[(3'h5):(3'h5)])
                    begin
                      reg1781 <= $signed((reg1623[(1'h1):(1'h1)] ?
                          ($unsigned((8'ha6)) ^ reg1739[(3'h4):(3'h4)]) : ({(8'ha1)} ?
                              $unsigned(wire1541) : (reg1673 | reg1663))));
                    end
                  else
                    begin
                      reg1781 <= $signed(reg1704);
                      reg1782 <= ((reg1563 - reg1571) ?
                          (|(reg1745[(2'h3):(1'h0)] ?
                              reg1582[(3'h5):(1'h0)] : $unsigned(reg1752))) : $signed(((reg1707 == reg1619) ?
                              reg1597 : reg1550)));
                      reg1783 <= $signed(((reg1766 ?
                              $signed(reg1675) : (reg1742 ?
                                  (8'ha2) : reg1682)) ?
                          $unsigned($signed(reg1598)) : reg1640));
                    end
                end
              for (forvar1784 = (1'h0); (forvar1784 < (2'h3)); forvar1784 = (forvar1784 + (1'h1)))
                begin
                  reg1785 <= $unsigned(($unsigned((~^reg1574)) ?
                      $signed(reg1624[(1'h0):(1'h0)]) : $signed($unsigned(reg1738))));
                  if ($signed((($signed(reg1664) == (wire1771 << reg1558)) ?
                      reg1724[(4'hc):(3'h7)] : $signed((^~reg1621)))))
                    begin
                      reg1786 <= $unsigned((reg1643 == reg1783));
                      reg1787 <= $signed($signed(reg1577));
                      reg1788 <= (&((reg1611 != {reg1775}) ?
                          $unsigned(reg1749) : reg1588));
                      reg1789 <= $unsigned(($signed(reg1582[(3'h5):(2'h3)]) ?
                          ((reg1683 == wire1545) & (wire1770 ?
                              reg1590 : reg1623)) : {$unsigned(reg1757)}));
                    end
                  else
                    begin
                      reg1786 <= (|(($unsigned(reg1785) >> reg1611) ?
                          (8'h9d) : $signed((reg1631 & reg1585))));
                      reg1787 <= $unsigned((reg1556 ?
                          ($unsigned(reg1661) ?
                              reg1650 : reg1623[(3'h4):(2'h3)]) : reg1570));
                      reg1788 <= (8'ha9);
                    end
                end
              for (forvar1790 = (1'h0); (forvar1790 < (1'h1)); forvar1790 = (forvar1790 + (1'h1)))
                begin
                  for (forvar1791 = (1'h0); (forvar1791 < (2'h3)); forvar1791 = (forvar1791 + (1'h1)))
                    begin
                      reg1792 <= (^$unsigned(($signed(reg1668) ~^ (reg1696 ?
                          reg1657 : reg1575))));
                    end
                end
            end
          for (forvar1793 = (1'h0); (forvar1793 < (1'h1)); forvar1793 = (forvar1793 + (1'h1)))
            begin
              if ($signed($unsigned($signed($unsigned((8'ha1))))))
                begin
                  for (forvar1794 = (1'h0); (forvar1794 < (2'h2)); forvar1794 = (forvar1794 + (1'h1)))
                    begin
                      reg1795 <= (~(^reg1591[(2'h3):(2'h2)]));
                      reg1796 <= (!(((8'h9d) ?
                          $unsigned(forvar1784) : (~reg1594)) << {{reg1673}}));
                    end
                  if (wire1544[(2'h3):(1'h1)])
                    begin
                      reg1797 <= (|$unsigned(reg1718[(3'h6):(3'h5)]));
                      reg1798 <= {$unsigned(reg1662[(4'h9):(3'h7)])};
                      reg1799 <= $unsigned({($signed(reg1786) + reg1730[(3'h5):(1'h1)])});
                      reg1800 <= ((8'hac) ?
                          (reg1707[(1'h1):(1'h0)] ?
                              {(reg1583 ?
                                      reg1681 : reg1737)} : $signed($signed(reg1581))) : (reg1646 ?
                              (8'hb3) : $signed((forvar1784 && reg1690))));
                    end
                  else
                    begin
                      reg1797 <= reg1624;
                      reg1798 <= $signed({((~^reg1690) | $signed(reg1590))});
                    end
                  if (((reg1594 ?
                          reg1674[(1'h1):(1'h0)] : reg1640[(3'h7):(2'h2)]) ?
                      (^$signed((forvar1773 ?
                          reg1636 : reg1568))) : (~|(reg1719[(2'h3):(2'h3)] + $signed(reg1619)))))
                    begin
                      reg1801 <= reg1567[(1'h0):(1'h0)];
                      reg1802 <= (((8'hb9) >>> (forvar1790 ?
                              (reg1557 < (8'hac)) : $signed((8'h9c)))) ?
                          {(~&reg1800[(2'h2):(1'h0)])} : (~&$signed((^reg1572))));
                    end
                  else
                    begin
                      reg1801 <= $unsigned(forvar1791[(2'h2):(1'h0)]);
                      reg1802 <= reg1657;
                      reg1803 <= reg1728;
                      reg1804 <= $unsigned((-reg1717));
                    end
                  if ((&$unsigned((-(reg1582 ? (8'hac) : reg1602)))))
                    begin
                      reg1805 <= (-($signed({reg1798}) ?
                          (8'hb3) : ({reg1711} >>> $unsigned(reg1743))));
                      reg1806 <= ((~&(~^reg1796)) == {(8'hae)});
                      reg1807 <= $signed({reg1689[(4'hb):(2'h3)]});
                      reg1808 <= (reg1712[(3'h5):(1'h1)] ?
                          forvar1773[(1'h1):(1'h1)] : $unsigned($unsigned((reg1712 ?
                              reg1686 : reg1640))));
                    end
                  else
                    begin
                      reg1805 <= (^reg1602[(1'h0):(1'h0)]);
                      reg1806 <= ((($unsigned((8'h9e)) ?
                          reg1756[(2'h2):(1'h1)] : (^reg1589)) + $unsigned($signed(forvar1790))) - {$signed((+reg1694))});
                      reg1807 <= ((&reg1683) & reg1751);
                      reg1808 <= $unsigned(reg1629);
                    end
                end
              else
                begin
                  reg1794 <= (((reg1776 ~^ reg1752[(1'h0):(1'h0)]) ^~ (8'hb7)) && ((8'haf) && {((8'had) <<< (8'hb1))}));
                  for (forvar1795 = (1'h0); (forvar1795 < (1'h0)); forvar1795 = (forvar1795 + (1'h1)))
                    begin
                      reg1796 <= (~^(8'hb9));
                      reg1797 <= ((reg1706 ?
                          (&(reg1702 ? reg1630 : reg1795)) : {(reg1764 ?
                                  reg1557 : reg1781)}) <= (8'hb8));
                      reg1798 <= $unsigned($signed($signed((reg1743 ?
                          reg1794 : reg1785))));
                      reg1799 <= (reg1719 ?
                          reg1700[(1'h1):(1'h1)] : reg1802[(3'h5):(2'h3)]);
                    end
                end
            end
          for (forvar1809 = (1'h0); (forvar1809 < (2'h2)); forvar1809 = (forvar1809 + (1'h1)))
            begin
              reg1810 <= $unsigned($unsigned((8'ha8)));
            end
        end
      else
        begin
          if (($signed($signed({reg1580})) & $unsigned(reg1806)))
            begin
              if (reg1744)
                begin
                  for (forvar1772 = (1'h0); (forvar1772 < (2'h3)); forvar1772 = (forvar1772 + (1'h1)))
                    begin
                      reg1773 <= (reg1701 << (($unsigned((8'ha6)) ?
                              (reg1633 ?
                                  (8'h9c) : reg1736) : $unsigned(reg1645)) ?
                          reg1663[(2'h3):(2'h3)] : (|reg1785)));
                      reg1774 <= $signed(reg1745);
                    end
                  for (forvar1775 = (1'h0); (forvar1775 < (2'h2)); forvar1775 = (forvar1775 + (1'h1)))
                    begin
                      reg1776 <= reg1675[(2'h3):(2'h2)];
                      reg1777 <= (8'ha0);
                      reg1778 <= $signed(reg1681);
                    end
                end
              else
                begin
                  for (forvar1772 = (1'h0); (forvar1772 < (1'h1)); forvar1772 = (forvar1772 + (1'h1)))
                    begin
                      reg1773 <= $signed(reg1591);
                      reg1774 <= {$unsigned((8'haa))};
                      reg1775 <= $unsigned(reg1694[(4'ha):(4'h9)]);
                    end
                  if ({reg1572[(4'hf):(4'hd)]})
                    begin
                      reg1776 <= (~|(8'ha6));
                      reg1777 <= {reg1554};
                      reg1778 <= (({$unsigned(reg1557)} - (^forvar1772[(2'h3):(2'h3)])) ?
                          (reg1616[(1'h0):(1'h0)] ?
                              {reg1759} : ((+forvar1791) ?
                                  $unsigned((8'hb6)) : {reg1608})) : reg1599[(3'h5):(3'h4)]);
                    end
                  else
                    begin
                      reg1776 <= reg1732;
                      reg1777 <= (~$signed({reg1645[(3'h5):(2'h3)]}));
                      reg1778 <= (reg1654[(3'h7):(3'h5)] ?
                          $unsigned((+reg1783)) : ($signed(reg1663) ?
                              $signed((|reg1622)) : (reg1648[(4'h9):(2'h3)] & reg1736[(3'h5):(2'h2)])));
                      reg1779 <= (reg1622[(1'h0):(1'h0)] ?
                          (-$unsigned((reg1742 ?
                              (8'hb9) : reg1700))) : ($unsigned((reg1613 ~^ reg1673)) << {(reg1802 & reg1755)}));
                    end
                end
            end
          else
            begin
              for (forvar1772 = (1'h0); (forvar1772 < (2'h3)); forvar1772 = (forvar1772 + (1'h1)))
                begin
                  for (forvar1773 = (1'h0); (forvar1773 < (2'h2)); forvar1773 = (forvar1773 + (1'h1)))
                    begin
                      reg1774 <= $unsigned($signed(reg1652));
                    end
                end
              if (reg1802[(1'h0):(1'h0)])
                begin
                  for (forvar1775 = (1'h0); (forvar1775 < (2'h3)); forvar1775 = (forvar1775 + (1'h1)))
                    begin
                      reg1776 <= reg1775;
                    end
                end
              else
                begin
                  if ($signed($unsigned($unsigned(reg1615))))
                    begin
                      reg1775 <= (|(+$signed(reg1556)));
                      reg1776 <= (-reg1732);
                      reg1777 <= $signed(($signed($signed(reg1665)) ?
                          (reg1768[(4'h8):(1'h1)] ?
                              reg1796 : reg1789[(1'h0):(1'h0)]) : reg1688[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg1775 <= (^($signed(((8'had) && reg1614)) == ($signed(reg1777) ?
                          {reg1592} : (reg1606 * (8'ha8)))));
                      reg1776 <= (^~reg1596[(1'h0):(1'h0)]);
                    end
                end
              for (forvar1778 = (1'h0); (forvar1778 < (1'h1)); forvar1778 = (forvar1778 + (1'h1)))
                begin
                  if ($signed($unsigned(reg1671[(4'h8):(4'h8)])))
                    begin
                      reg1779 <= reg1563[(1'h0):(1'h0)];
                      reg1780 <= $unsigned(reg1741);
                      reg1781 <= ($unsigned(reg1596) <= $unsigned(reg1615));
                    end
                  else
                    begin
                      reg1779 <= reg1728;
                      reg1780 <= (reg1732[(4'h8):(3'h5)] ?
                          $unsigned(((8'h9f) ?
                              $signed(reg1707) : {reg1778})) : {((reg1786 ^~ reg1798) ?
                                  (+reg1626) : (!reg1644))});
                    end
                  for (forvar1782 = (1'h0); (forvar1782 < (2'h2)); forvar1782 = (forvar1782 + (1'h1)))
                    begin
                      reg1783 <= reg1587[(2'h2):(1'h1)];
                    end
                  reg1784 <= wire1544;
                  if (reg1653[(4'h8):(3'h6)])
                    begin
                      reg1785 <= ((-reg1717[(4'hc):(3'h5)]) ?
                          (~&($unsigned(reg1582) ^ (reg1804 >= reg1806))) : (+reg1807));
                    end
                  else
                    begin
                      reg1785 <= $unsigned($unsigned(((reg1792 <<< reg1635) ?
                          (reg1797 ?
                              reg1781 : (8'hb8)) : reg1633[(1'h1):(1'h0)])));
                      reg1786 <= reg1649[(2'h2):(1'h0)];
                      reg1787 <= ({$unsigned({(8'ha5)})} ?
                          reg1779 : $signed(({reg1727} ?
                              $signed(reg1743) : (wire1543 | reg1615))));
                    end
                end
              for (forvar1788 = (1'h0); (forvar1788 < (1'h0)); forvar1788 = (forvar1788 + (1'h1)))
                begin
                  if (reg1568[(2'h2):(1'h1)])
                    begin
                      reg1789 <= ((^~reg1807) ^~ (forvar1795 ?
                          $signed((~|(8'ha1))) : reg1567));
                    end
                  else
                    begin
                      reg1789 <= $unsigned(($unsigned((8'hae)) ?
                          (8'hb0) : (((8'ha5) > reg1591) < $signed(wire1771))));
                    end
                  if ((~^(&$signed(((8'hb0) ? (8'ha5) : reg1795)))))
                    begin
                      reg1790 <= $unsigned((^$signed((^~reg1678))));
                      reg1791 <= $unsigned(($unsigned({reg1690}) ?
                          $signed($unsigned(forvar1773)) : ($unsigned(reg1653) ?
                              reg1620[(3'h4):(1'h0)] : ((8'hb4) * forvar1793))));
                      reg1792 <= $unsigned(((!((8'ha4) ^ forvar1778)) >>> {(-reg1643)}));
                    end
                  else
                    begin
                      reg1790 <= reg1706[(1'h0):(1'h0)];
                      reg1791 <= reg1787;
                    end
                end
            end
          if ((-((8'hab) >>> reg1721[(2'h2):(1'h0)])))
            begin
              if (({reg1568} ?
                  $signed($unsigned(((8'h9d) ?
                      (8'ha2) : wire1546))) : (reg1780[(4'h8):(1'h0)] * (^~(reg1802 ?
                      reg1613 : reg1746)))))
                begin
                  for (forvar1793 = (1'h0); (forvar1793 < (2'h2)); forvar1793 = (forvar1793 + (1'h1)))
                    begin
                      reg1794 <= reg1686;
                      reg1795 <= reg1664;
                      reg1796 <= {$signed(forvar1791)};
                      reg1797 <= reg1802[(3'h4):(1'h0)];
                    end
                end
              else
                begin
                  if (reg1623)
                    begin
                      reg1793 <= wire1547;
                      reg1794 <= (reg1806[(3'h5):(1'h1)] ?
                          $unsigned(reg1593[(2'h3):(2'h3)]) : $signed(((reg1722 ?
                              (8'hae) : (8'ha0)) < (reg1751 | reg1600))));
                      reg1795 <= (8'h9c);
                    end
                  else
                    begin
                      reg1793 <= (($signed(reg1620) && $signed(reg1691[(2'h3):(2'h3)])) > $unsigned($signed(reg1573[(4'hc):(3'h6)])));
                      reg1794 <= ((($unsigned(reg1668) * (+reg1719)) ?
                              $unsigned($unsigned(reg1663)) : reg1555[(3'h4):(1'h0)]) ?
                          (reg1658[(2'h2):(1'h1)] ~^ {(reg1646 ^ reg1600)}) : reg1761);
                      reg1795 <= {($signed(((8'h9f) ?
                              reg1764 : (8'haa))) || (8'ha4))};
                      reg1796 <= $signed($signed($unsigned(((8'hb1) ?
                          reg1641 : reg1704))));
                    end
                  for (forvar1797 = (1'h0); (forvar1797 < (1'h1)); forvar1797 = (forvar1797 + (1'h1)))
                    begin
                      reg1798 <= {($unsigned((~&reg1702)) * (!forvar1795[(4'hf):(2'h2)]))};
                    end
                  for (forvar1799 = (1'h0); (forvar1799 < (1'h1)); forvar1799 = (forvar1799 + (1'h1)))
                    begin
                      reg1800 <= reg1642[(4'h8):(3'h5)];
                      reg1801 <= reg1608[(4'ha):(3'h6)];
                    end
                  reg1802 <= reg1744;
                end
              for (forvar1803 = (1'h0); (forvar1803 < (2'h3)); forvar1803 = (forvar1803 + (1'h1)))
                begin
                  if (reg1729)
                    begin
                      reg1804 <= reg1802;
                      reg1805 <= reg1590;
                    end
                  else
                    begin
                      reg1804 <= reg1740;
                    end
                  for (forvar1806 = (1'h0); (forvar1806 < (1'h1)); forvar1806 = (forvar1806 + (1'h1)))
                    begin
                      reg1807 <= $signed((reg1686 >= $unsigned((reg1777 ^~ (8'ha7)))));
                    end
                  if ((~reg1588))
                    begin
                      reg1808 <= $signed(reg1789[(3'h4):(2'h3)]);
                      reg1809 <= (~(8'haa));
                      reg1810 <= ((8'ha9) >= (8'hb4));
                      reg1811 <= ((8'h9d) ^ {reg1629[(4'ha):(3'h6)]});
                    end
                  else
                    begin
                      reg1808 <= (reg1584[(2'h2):(2'h2)] ?
                          $unsigned((|reg1633)) : {reg1658});
                    end
                end
            end
          else
            begin
              if (((8'haa) ^ ($signed((reg1745 && reg1720)) ?
                  ($signed(reg1780) ?
                      {(8'hac)} : {reg1587}) : reg1608[(4'hc):(2'h3)])))
                begin
                  if ((!(!reg1724)))
                    begin
                      reg1793 <= reg1639[(1'h1):(1'h1)];
                      reg1794 <= reg1570[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg1793 <= (reg1742 ^~ (reg1773[(1'h0):(1'h0)] ?
                          $unsigned({reg1746}) : {$unsigned(reg1756)}));
                      reg1794 <= $signed($unsigned(reg1739));
                    end
                end
              else
                begin
                  reg1793 <= (((-$signed(reg1615)) + $unsigned((reg1556 << reg1689))) ?
                      ($unsigned({reg1574}) ?
                          $unsigned($signed(reg1752)) : $unsigned((reg1794 ^~ forvar1809))) : (~&(reg1782 ~^ reg1745[(1'h1):(1'h0)])));
                  for (forvar1794 = (1'h0); (forvar1794 < (1'h1)); forvar1794 = (forvar1794 + (1'h1)))
                    begin
                      reg1795 <= (((+reg1664) ^ (+(8'ha8))) ?
                          reg1787 : (~|(reg1613[(2'h3):(2'h3)] ?
                              (-reg1683) : (reg1801 ? reg1583 : reg1594))));
                      reg1796 <= (reg1661 <<< (|reg1698[(3'h6):(2'h3)]));
                    end
                  for (forvar1797 = (1'h0); (forvar1797 < (1'h0)); forvar1797 = (forvar1797 + (1'h1)))
                    begin
                      reg1798 <= $unsigned(reg1632);
                    end
                end
              for (forvar1799 = (1'h0); (forvar1799 < (2'h2)); forvar1799 = (forvar1799 + (1'h1)))
                begin
                  if ((8'ha5))
                    begin
                      reg1800 <= $signed((reg1784 << reg1596[(1'h0):(1'h0)]));
                      reg1801 <= forvar1794[(4'he):(4'ha)];
                    end
                  else
                    begin
                      reg1800 <= $signed(reg1710[(4'h9):(3'h6)]);
                    end
                end
            end
        end
    end
  assign wire1812 = reg1781[(1'h0):(1'h0)];
  assign wire1813 = $unsigned(((~&$signed(reg1599)) ?
                        ($unsigned(reg1661) ?
                            $unsigned(reg1591) : (reg1776 >= reg1757)) : $unsigned($signed(reg1743))));
  assign wire1814 = (($signed(reg1750[(4'h8):(3'h6)]) ?
                        {$unsigned(reg1608)} : wire1546) && $signed((-(reg1782 << reg1714))));
  assign wire1815 = reg1657;
  assign wire1816 = $signed((!reg1679[(2'h3):(1'h0)]));
  always
    @(posedge clk) begin
      if (reg1681[(4'h8):(4'h8)])
        begin
          for (forvar1817 = (1'h0); (forvar1817 < (1'h0)); forvar1817 = (forvar1817 + (1'h1)))
            begin
              reg1818 <= (($unsigned((&reg1693)) || {(reg1616 ?
                          reg1776 : reg1550)}) ?
                  ((-(reg1596 ? reg1746 : reg1597)) ?
                      (^~$unsigned(reg1627)) : reg1613[(1'h1):(1'h0)]) : reg1773[(3'h5):(3'h4)]);
            end
          if ({$signed(reg1572)})
            begin
              for (forvar1819 = (1'h0); (forvar1819 < (2'h2)); forvar1819 = (forvar1819 + (1'h1)))
                begin
                  if (($signed(($unsigned(reg1674) ?
                      reg1729 : $signed(reg1756))) != $unsigned((+(reg1549 || (8'ha4))))))
                    begin
                      reg1820 <= {reg1742[(4'ha):(1'h1)]};
                    end
                  else
                    begin
                      reg1820 <= reg1784;
                    end
                  for (forvar1821 = (1'h0); (forvar1821 < (2'h2)); forvar1821 = (forvar1821 + (1'h1)))
                    begin
                      reg1822 <= reg1776;
                    end
                  for (forvar1823 = (1'h0); (forvar1823 < (1'h1)); forvar1823 = (forvar1823 + (1'h1)))
                    begin
                      reg1824 <= $signed((reg1729[(2'h3):(1'h0)] ?
                          (^~(reg1749 * reg1751)) : $signed(reg1706[(4'hd):(3'h4)])));
                      reg1825 <= (~&(^(((8'hb1) ?
                          reg1629 : (8'ha6)) < {reg1804})));
                      reg1826 <= ($unsigned((|(~^reg1627))) == $unsigned((reg1803 ?
                          reg1681 : $unsigned((8'haf)))));
                    end
                  if ((~|(reg1729[(4'h8):(3'h6)] ^~ ($unsigned(reg1639) ?
                      (reg1759 ? reg1794 : reg1738) : (reg1556 ?
                          (8'hb2) : reg1608)))))
                    begin
                      reg1827 <= reg1623;
                      reg1828 <= $unsigned((&((reg1630 ? reg1783 : reg1634) ?
                          reg1680 : (^forvar1821))));
                      reg1829 <= reg1732;
                      reg1830 <= (($signed((reg1774 >>> reg1750)) ?
                          $signed((8'ha0)) : forvar1823[(4'h8):(3'h4)]) ~^ {reg1685[(3'h5):(1'h1)]});
                    end
                  else
                    begin
                      reg1827 <= reg1801;
                      reg1828 <= (reg1730 != (8'hb1));
                      reg1829 <= reg1550;
                      reg1830 <= $signed({$signed(reg1556)});
                    end
                end
              for (forvar1831 = (1'h0); (forvar1831 < (1'h0)); forvar1831 = (forvar1831 + (1'h1)))
                begin
                  for (forvar1832 = (1'h0); (forvar1832 < (2'h3)); forvar1832 = (forvar1832 + (1'h1)))
                    begin
                      reg1833 <= {(^~$signed(reg1674[(1'h1):(1'h0)]))};
                    end
                  if (((~&(~^$signed(reg1661))) ?
                      reg1725 : $unsigned(({reg1808} ?
                          $unsigned(reg1709) : $unsigned(reg1624)))))
                    begin
                      reg1834 <= reg1574[(3'h5):(1'h0)];
                      reg1835 <= $signed(reg1590);
                      reg1836 <= (reg1737[(2'h3):(1'h0)] ?
                          reg1563[(1'h1):(1'h0)] : $unsigned($unsigned((reg1608 ?
                              reg1611 : reg1768))));
                    end
                  else
                    begin
                      reg1834 <= $unsigned((!$signed((|reg1742))));
                    end
                end
              if (reg1822)
                begin
                  for (forvar1837 = (1'h0); (forvar1837 < (1'h0)); forvar1837 = (forvar1837 + (1'h1)))
                    begin
                      reg1838 <= (~|{reg1596[(1'h1):(1'h1)]});
                    end
                  for (forvar1839 = (1'h0); (forvar1839 < (2'h2)); forvar1839 = (forvar1839 + (1'h1)))
                    begin
                      reg1840 <= $signed(($signed($signed(reg1788)) & (|reg1777[(4'h9):(1'h1)])));
                      reg1841 <= {$signed(((reg1763 ? (8'h9d) : reg1627) ?
                              $signed(reg1719) : reg1778))};
                    end
                  for (forvar1842 = (1'h0); (forvar1842 < (2'h3)); forvar1842 = (forvar1842 + (1'h1)))
                    begin
                      reg1843 <= (-((&reg1791[(2'h2):(2'h2)]) >>> reg1753[(2'h3):(2'h2)]));
                      reg1844 <= $signed(reg1811[(4'ha):(4'h8)]);
                    end
                  for (forvar1845 = (1'h0); (forvar1845 < (1'h0)); forvar1845 = (forvar1845 + (1'h1)))
                    begin
                      reg1846 <= reg1644;
                    end
                end
              else
                begin
                  reg1837 <= reg1808[(3'h5):(2'h2)];
                end
              reg1847 <= ((reg1745[(3'h4):(1'h0)] ?
                      (reg1701[(2'h3):(1'h0)] ?
                          reg1555[(1'h1):(1'h1)] : $signed(wire1546)) : $signed(reg1659)) ?
                  reg1703 : $signed((reg1609[(2'h2):(1'h0)] ?
                      ((8'ha9) ? wire1544 : reg1786) : $unsigned(reg1668))));
            end
          else
            begin
              for (forvar1819 = (1'h0); (forvar1819 < (2'h2)); forvar1819 = (forvar1819 + (1'h1)))
                begin
                  for (forvar1820 = (1'h0); (forvar1820 < (1'h0)); forvar1820 = (forvar1820 + (1'h1)))
                    begin
                      reg1821 <= (({(reg1808 != reg1640)} >>> (|reg1700)) - (reg1590[(2'h2):(2'h2)] ?
                          (^~(8'hb7)) : reg1570[(3'h4):(1'h1)]));
                      reg1822 <= $signed((reg1843[(1'h1):(1'h0)] ?
                          {$signed(reg1628)} : (-(8'ha9))));
                      reg1823 <= reg1786[(1'h1):(1'h0)];
                    end
                end
              if ($unsigned({($signed(reg1788) ? (|(8'hac)) : reg1841)}))
                begin
                  for (forvar1824 = (1'h0); (forvar1824 < (1'h1)); forvar1824 = (forvar1824 + (1'h1)))
                    begin
                      reg1825 <= $signed(({(reg1835 ? reg1776 : reg1776)} ?
                          (reg1776[(3'h5):(2'h2)] ?
                              reg1614 : $unsigned((8'hba))) : (~&(reg1783 < reg1712))));
                      reg1826 <= $unsigned((~|(^(reg1601 ?
                          (8'ha4) : reg1651))));
                    end
                end
              else
                begin
                  if (forvar1823[(4'h8):(1'h0)])
                    begin
                      reg1824 <= ($signed(reg1716[(2'h3):(1'h0)]) ?
                          $signed({reg1596[(1'h0):(1'h0)]}) : ($signed($signed(reg1576)) << reg1603));
                      reg1825 <= wire1814;
                    end
                  else
                    begin
                      reg1824 <= {reg1809};
                      reg1825 <= reg1829[(3'h7):(2'h3)];
                      reg1826 <= (8'haf);
                      reg1827 <= (^~(~^(~reg1629)));
                    end
                  for (forvar1828 = (1'h0); (forvar1828 < (2'h3)); forvar1828 = (forvar1828 + (1'h1)))
                    begin
                      reg1829 <= $signed(reg1623[(1'h0):(1'h0)]);
                      reg1830 <= (reg1658[(2'h3):(1'h0)] ?
                          $unsigned({$unsigned(reg1581)}) : $signed(reg1745[(3'h5):(2'h3)]));
                      reg1831 <= ({{(-reg1757)}} ?
                          (($signed(reg1614) ^ $unsigned(reg1775)) < $signed(reg1826[(1'h0):(1'h0)])) : (!$unsigned((wire1541 ?
                              reg1615 : reg1802))));
                      reg1832 <= $signed(($unsigned(reg1711) ?
                          reg1749 : (~^reg1620)));
                    end
                  if (reg1670[(1'h1):(1'h1)])
                    begin
                      reg1833 <= $unsigned((^$unsigned($unsigned(reg1789))));
                      reg1834 <= reg1675[(3'h7):(1'h0)];
                      reg1835 <= (~$unsigned(reg1601));
                      reg1836 <= reg1635;
                    end
                  else
                    begin
                      reg1833 <= reg1667[(1'h0):(1'h0)];
                      reg1834 <= reg1745;
                      reg1835 <= reg1690[(1'h0):(1'h0)];
                    end
                end
              if (({$unsigned({reg1792})} ~^ (~^forvar1823)))
                begin
                  for (forvar1837 = (1'h0); (forvar1837 < (2'h2)); forvar1837 = (forvar1837 + (1'h1)))
                    begin
                      reg1838 <= $unsigned($unsigned((~|reg1678[(2'h2):(1'h0)])));
                      reg1839 <= (~^(^~((8'hb4) < $unsigned(reg1685))));
                    end
                  reg1840 <= reg1668;
                end
              else
                begin
                  if (reg1551[(2'h2):(1'h0)])
                    begin
                      reg1837 <= (-({{(8'ha1)}} ?
                          ({reg1742} && (reg1740 ?
                              reg1761 : reg1679)) : (((8'ha7) ?
                              reg1789 : reg1777) && (~^reg1606))));
                    end
                  else
                    begin
                      reg1837 <= $signed(reg1758);
                      reg1838 <= $unsigned((^reg1622[(2'h3):(1'h0)]));
                      reg1839 <= $unsigned((reg1710 & reg1606[(3'h4):(2'h3)]));
                    end
                  for (forvar1840 = (1'h0); (forvar1840 < (2'h2)); forvar1840 = (forvar1840 + (1'h1)))
                    begin
                      reg1841 <= reg1586;
                      reg1842 <= {(^reg1790)};
                      reg1843 <= (+$unsigned({reg1553[(4'h8):(3'h6)]}));
                    end
                end
            end
        end
      else
        begin
          reg1817 <= ($unsigned((~^$unsigned(reg1835))) ?
              ((~^(reg1594 ? reg1594 : wire1546)) ?
                  ($unsigned(reg1799) ?
                      ((8'ha8) ^~ reg1570) : (+reg1561)) : $unsigned(((8'ha4) ?
                      (8'hb2) : reg1678))) : (forvar1837[(1'h1):(1'h1)] ?
                  $signed(reg1639) : (~^(reg1786 ? reg1642 : reg1759))));
          for (forvar1818 = (1'h0); (forvar1818 < (1'h0)); forvar1818 = (forvar1818 + (1'h1)))
            begin
              if ((+((^(reg1704 ? reg1691 : wire1544)) ?
                  (&(|reg1667)) : ($unsigned(reg1644) & reg1587[(3'h5):(1'h0)]))))
                begin
                  if (((reg1587 ?
                      $signed((^reg1798)) : ($unsigned(reg1810) == (reg1561 <= reg1714))) >> $signed($unsigned($unsigned(reg1724)))))
                    begin
                      reg1819 <= (!(reg1646[(3'h5):(1'h1)] ?
                          ((!(8'ha6)) ?
                              reg1843[(1'h1):(1'h0)] : (reg1659 ?
                                  reg1731 : reg1594)) : wire1545));
                      reg1820 <= reg1551[(1'h1):(1'h0)];
                      reg1821 <= ($unsigned(((~&(8'hac)) == $signed(reg1716))) ?
                          (reg1662[(2'h3):(1'h1)] ?
                              ($unsigned(reg1786) & $signed(reg1640)) : reg1773) : (^reg1701));
                      reg1822 <= {$signed(($unsigned(reg1759) == $unsigned(reg1575)))};
                    end
                  else
                    begin
                      reg1819 <= $unsigned((reg1602 ?
                          $signed((~^reg1792)) : reg1789));
                    end
                  if ((reg1789[(3'h5):(3'h4)] >>> $signed(reg1751[(4'h8):(2'h2)])))
                    begin
                      reg1823 <= (-$signed({reg1668}));
                      reg1824 <= (|($unsigned((reg1580 == (8'hae))) > reg1685[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1823 <= (reg1783[(3'h4):(1'h1)] ?
                          (~^reg1724[(4'h8):(3'h6)]) : $signed($signed(reg1804[(3'h7):(1'h1)])));
                    end
                  reg1825 <= {(reg1553 - (&$unsigned(reg1738)))};
                  for (forvar1826 = (1'h0); (forvar1826 < (2'h2)); forvar1826 = (forvar1826 + (1'h1)))
                    begin
                      reg1827 <= {$signed(reg1829)};
                      reg1828 <= {((^~$unsigned(wire1547)) ?
                              (-$signed(reg1602)) : {reg1810})};
                      reg1829 <= (+$signed((-$unsigned(reg1733))));
                      reg1830 <= $signed($unsigned((8'hb0)));
                    end
                end
              else
                begin
                  reg1819 <= reg1824[(2'h2):(1'h0)];
                  for (forvar1820 = (1'h0); (forvar1820 < (2'h2)); forvar1820 = (forvar1820 + (1'h1)))
                    begin
                      reg1821 <= {$signed(reg1801)};
                      reg1822 <= $unsigned((((~&reg1710) ?
                              $signed(reg1741) : reg1641[(1'h1):(1'h0)]) ?
                          {$unsigned(reg1838)} : (8'h9e)));
                      reg1823 <= $unsigned((8'hb6));
                    end
                  reg1824 <= $signed({$signed(reg1574)});
                end
              for (forvar1831 = (1'h0); (forvar1831 < (1'h0)); forvar1831 = (forvar1831 + (1'h1)))
                begin
                  if (((((reg1665 ?
                      reg1839 : reg1698) ^~ {(8'h9c)}) <= ((reg1653 ?
                          wire1815 : (8'h9f)) ?
                      (reg1792 ?
                          reg1563 : (8'hb8)) : $unsigned(reg1729))) >>> reg1713))
                    begin
                      reg1832 <= ($signed(($unsigned(reg1798) ?
                              reg1709[(3'h7):(3'h5)] : reg1837)) ?
                          reg1800 : (!(~^reg1836)));
                      reg1833 <= (~|(-(^$unsigned(reg1653))));
                    end
                  else
                    begin
                      reg1832 <= ((8'ha9) && $unsigned(({reg1555} - reg1636)));
                      reg1833 <= reg1727[(2'h3):(1'h0)];
                    end
                  for (forvar1834 = (1'h0); (forvar1834 < (2'h2)); forvar1834 = (forvar1834 + (1'h1)))
                    begin
                      reg1835 <= ((|(reg1696 && reg1827)) >= (^$unsigned((~|(8'h9f)))));
                      reg1836 <= {((!$signed(reg1631)) && (reg1693[(3'h5):(1'h1)] ?
                              (reg1575 ?
                                  reg1762 : reg1606) : reg1737[(4'h8):(3'h6)]))};
                      reg1837 <= $signed($unsigned($unsigned($unsigned(reg1711))));
                    end
                  reg1838 <= reg1834;
                  for (forvar1839 = (1'h0); (forvar1839 < (2'h3)); forvar1839 = (forvar1839 + (1'h1)))
                    begin
                      reg1840 <= ((8'ha0) >> ({(+reg1847)} != ($unsigned((8'hab)) ?
                          (forvar1840 || reg1614) : $signed(reg1713))));
                      reg1841 <= ((-$unsigned(((8'hae) ~^ reg1743))) ?
                          reg1721 : (^~reg1591[(4'hc):(3'h5)]));
                      reg1842 <= (reg1836 ?
                          $unsigned((~$signed(forvar1818))) : {reg1621});
                    end
                end
              reg1843 <= (^{($signed(reg1709) ?
                      $unsigned(reg1675) : (reg1554 * forvar1839))});
              reg1844 <= ((^reg1563[(2'h3):(2'h2)]) ?
                  ((reg1595 ? reg1624[(2'h3):(1'h0)] : $signed(reg1589)) ?
                      (forvar1828[(3'h4):(3'h4)] ?
                          (reg1725 || reg1704) : (^reg1831)) : reg1840) : ($signed($signed(reg1617)) ?
                      $signed(reg1675[(3'h4):(2'h3)]) : $signed((reg1636 ?
                          (8'h9d) : reg1619))));
            end
          for (forvar1845 = (1'h0); (forvar1845 < (2'h2)); forvar1845 = (forvar1845 + (1'h1)))
            begin
              if ((((~((8'hac) >= reg1627)) ^ $unsigned($unsigned(reg1738))) ?
                  reg1619 : reg1837))
                begin
                  for (forvar1846 = (1'h0); (forvar1846 < (2'h2)); forvar1846 = (forvar1846 + (1'h1)))
                    begin
                      reg1847 <= (+$signed(reg1581));
                    end
                  if (reg1665)
                    begin
                      reg1848 <= ($signed((reg1703[(4'ha):(2'h3)] ?
                          ((8'ha5) ^~ reg1733) : (^reg1668))) == $unsigned((+((8'hb8) <= (8'hba)))));
                      reg1849 <= reg1740[(3'h4):(2'h3)];
                      reg1850 <= ($signed(($signed(reg1651) < forvar1832[(1'h0):(1'h0)])) ?
                          (~^(+reg1582[(3'h5):(2'h3)])) : ($unsigned(reg1694) || (reg1635[(4'ha):(4'h9)] ?
                              reg1757[(1'h1):(1'h0)] : reg1586)));
                      reg1851 <= ((8'h9c) <= $unsigned(($unsigned(reg1808) << reg1573[(3'h6):(3'h5)])));
                    end
                  else
                    begin
                      reg1848 <= $signed(($unsigned((reg1570 ?
                          wire1542 : reg1795)) <<< reg1729));
                      reg1849 <= (8'ha1);
                    end
                end
              else
                begin
                  for (forvar1846 = (1'h0); (forvar1846 < (1'h0)); forvar1846 = (forvar1846 + (1'h1)))
                    begin
                      reg1847 <= $unsigned(reg1788);
                      reg1848 <= reg1834[(2'h2):(1'h1)];
                    end
                end
              if ((~|forvar1823[(4'h8):(3'h6)]))
                begin
                  for (forvar1852 = (1'h0); (forvar1852 < (1'h0)); forvar1852 = (forvar1852 + (1'h1)))
                    begin
                      reg1853 <= $unsigned((-{$unsigned(reg1838)}));
                      reg1854 <= (reg1831 ^ (reg1556[(2'h3):(1'h0)] != ($unsigned(reg1658) >= reg1647)));
                    end
                  for (forvar1855 = (1'h0); (forvar1855 < (2'h2)); forvar1855 = (forvar1855 + (1'h1)))
                    begin
                      reg1856 <= (|$signed(reg1844[(3'h7):(3'h5)]));
                      reg1857 <= ($signed(reg1840[(4'hb):(2'h3)]) || ((~&(reg1722 + reg1678)) | ({reg1657} <<< (reg1549 ?
                          wire1542 : reg1590))));
                      reg1858 <= {reg1716};
                      reg1859 <= (|(~&((reg1573 << forvar1832) != $unsigned(reg1829))));
                    end
                  for (forvar1860 = (1'h0); (forvar1860 < (1'h0)); forvar1860 = (forvar1860 + (1'h1)))
                    begin
                      reg1861 <= {(reg1717[(4'h9):(1'h1)] > reg1798[(1'h0):(1'h0)])};
                      reg1862 <= $signed($unsigned($signed($signed(reg1839))));
                      reg1863 <= reg1647;
                    end
                end
              else
                begin
                  if (reg1743)
                    begin
                      reg1852 <= (reg1749 ^ {($signed((8'h9e)) << $unsigned(reg1630))});
                      reg1853 <= $unsigned(reg1558);
                      reg1854 <= (~reg1786[(2'h3):(1'h0)]);
                    end
                  else
                    begin
                      reg1852 <= reg1778[(4'hb):(4'hb)];
                      reg1853 <= ((~&(reg1774 || {reg1794})) ?
                          (|((+reg1701) | $signed(reg1595))) : $signed(($signed(reg1607) ?
                              (&reg1590) : $unsigned(reg1648))));
                    end
                  if ($unsigned(reg1614))
                    begin
                      reg1855 <= (^~$unsigned($signed((!reg1755))));
                    end
                  else
                    begin
                      reg1855 <= $unsigned($unsigned((((8'haa) ^ (8'haa)) <= (|reg1590))));
                      reg1856 <= $unsigned((!(reg1781[(4'h8):(2'h2)] << $unsigned(wire1546))));
                      reg1857 <= reg1804;
                      reg1858 <= (reg1795 + $unsigned(reg1572));
                    end
                  for (forvar1859 = (1'h0); (forvar1859 < (1'h0)); forvar1859 = (forvar1859 + (1'h1)))
                    begin
                      reg1860 <= $signed(((!(!(8'hb4))) ?
                          (~(~reg1601)) : $signed($signed(reg1811))));
                    end
                  for (forvar1861 = (1'h0); (forvar1861 < (2'h2)); forvar1861 = (forvar1861 + (1'h1)))
                    begin
                      reg1862 <= ((8'h9c) >> ($signed((reg1829 > reg1820)) * reg1729[(4'h8):(3'h6)]));
                      reg1863 <= (reg1704 & forvar1855[(2'h3):(2'h2)]);
                      reg1864 <= reg1632[(1'h1):(1'h1)];
                    end
                end
            end
          if ((~|$signed(reg1667)))
            begin
              if ($unsigned($unsigned(((reg1825 ^ reg1558) ^~ (reg1750 ?
                  (8'hb7) : reg1701)))))
                begin
                  for (forvar1865 = (1'h0); (forvar1865 < (1'h0)); forvar1865 = (forvar1865 + (1'h1)))
                    begin
                      reg1866 <= ((~((^~(8'ha2)) ?
                              reg1601 : (forvar1820 ? reg1717 : reg1681))) ?
                          forvar1846[(3'h4):(1'h1)] : $unsigned((reg1861 ^~ (reg1750 ?
                              (8'had) : reg1782))));
                      reg1867 <= (~&(($unsigned(reg1553) ?
                              (reg1662 || reg1847) : (reg1602 ?
                                  reg1597 : reg1550)) ?
                          reg1586 : (reg1731[(1'h1):(1'h0)] ?
                              ((8'h9f) ?
                                  reg1632 : wire1545) : $signed(wire1812))));
                      reg1868 <= {($unsigned((reg1600 ?
                              reg1714 : reg1745)) || (8'h9c))};
                      reg1869 <= (|(reg1632[(1'h1):(1'h1)] && $unsigned($signed((8'ha1)))));
                    end
                end
              else
                begin
                  for (forvar1865 = (1'h0); (forvar1865 < (1'h1)); forvar1865 = (forvar1865 + (1'h1)))
                    begin
                      reg1866 <= forvar1820;
                      reg1867 <= reg1628;
                      reg1868 <= $unsigned({($unsigned(reg1669) ?
                              (!reg1861) : {reg1665})});
                    end
                  if (wire1544)
                    begin
                      reg1869 <= (({{reg1733}} ?
                              (!reg1832[(4'hc):(4'hb)]) : (~reg1663)) ?
                          (+$signed(((8'ha2) ?
                              (8'h9e) : reg1736))) : $signed(((-reg1702) ?
                              $unsigned(reg1634) : (reg1691 ?
                                  reg1832 : reg1785))));
                    end
                  else
                    begin
                      reg1869 <= reg1857[(2'h2):(2'h2)];
                      reg1870 <= reg1744[(4'h9):(1'h1)];
                    end
                  if ((8'hb1))
                    begin
                      reg1871 <= {reg1867};
                      reg1872 <= reg1836[(2'h2):(1'h1)];
                      reg1873 <= reg1864[(4'hb):(4'h9)];
                      reg1874 <= $unsigned((reg1861 || reg1654));
                    end
                  else
                    begin
                      reg1871 <= reg1761[(4'h9):(4'h8)];
                      reg1872 <= $signed(reg1713[(3'h6):(1'h1)]);
                      reg1873 <= ((reg1806[(3'h5):(2'h2)] & (~|((8'ha6) >= reg1744))) ?
                          (^reg1631) : $unsigned(reg1649[(2'h3):(2'h2)]));
                    end
                  for (forvar1875 = (1'h0); (forvar1875 < (1'h0)); forvar1875 = (forvar1875 + (1'h1)))
                    begin
                      reg1876 <= (8'ha4);
                      reg1877 <= reg1805;
                      reg1878 <= $unsigned((-$unsigned($unsigned(forvar1824))));
                    end
                end
              for (forvar1879 = (1'h0); (forvar1879 < (2'h2)); forvar1879 = (forvar1879 + (1'h1)))
                begin
                  if ($unsigned({$unsigned((~^reg1712))}))
                    begin
                      reg1880 <= $signed((((+reg1731) ^~ (reg1603 ?
                              (8'hb2) : reg1740)) ?
                          reg1607[(4'hb):(4'ha)] : $signed(forvar1846[(2'h2):(1'h0)])));
                      reg1881 <= (~&((+(forvar1828 ^~ reg1849)) ?
                          {(|reg1664)} : {$unsigned(reg1550)}));
                      reg1882 <= reg1866[(1'h1):(1'h0)];
                      reg1883 <= $unsigned((reg1671 ?
                          $unsigned((reg1838 & reg1721)) : $unsigned((!reg1796))));
                    end
                  else
                    begin
                      reg1880 <= (~^reg1757);
                      reg1881 <= $unsigned((((&forvar1823) ?
                              (&reg1830) : $unsigned((8'h9c))) ?
                          $signed($unsigned(reg1835)) : ((~&reg1801) ?
                              $signed(reg1596) : forvar1875[(1'h1):(1'h1)])));
                      reg1882 <= $signed($unsigned((reg1713[(3'h4):(3'h4)] ?
                          reg1791 : (reg1593 >>> forvar1821))));
                      reg1883 <= $unsigned(reg1743[(3'h4):(3'h4)]);
                    end
                end
              reg1884 <= (^~forvar1834[(2'h2):(1'h0)]);
            end
          else
            begin
              reg1865 <= ({$signed(((8'hab) ?
                      reg1762 : reg1774))} - ({(reg1784 >> reg1834)} ?
                  reg1657 : reg1570[(3'h5):(1'h1)]));
              if ((~&$signed(({reg1574} >>> {reg1720}))))
                begin
                  for (forvar1866 = (1'h0); (forvar1866 < (2'h3)); forvar1866 = (forvar1866 + (1'h1)))
                    begin
                      reg1867 <= reg1641[(1'h1):(1'h0)];
                      reg1868 <= $signed((-((~|reg1549) >>> $unsigned(reg1863))));
                      reg1869 <= reg1555;
                    end
                  reg1870 <= (~^$signed((~&$signed(reg1862))));
                  reg1871 <= {({$unsigned(reg1669)} ?
                          $signed(reg1644) : forvar1842[(4'h9):(2'h3)])};
                  for (forvar1872 = (1'h0); (forvar1872 < (1'h0)); forvar1872 = (forvar1872 + (1'h1)))
                    begin
                      reg1873 <= (-(!reg1876));
                      reg1874 <= reg1568[(4'hc):(1'h1)];
                      reg1875 <= ($signed(reg1794) ?
                          (reg1731 ~^ (^(^reg1665))) : {reg1741[(2'h3):(2'h2)]});
                    end
                end
              else
                begin
                  reg1866 <= $signed(((~^reg1563) ?
                      $signed((reg1658 < reg1756)) : $signed(reg1710)));
                  if ((+(-{(reg1839 ^ reg1827)})))
                    begin
                      reg1867 <= reg1586;
                      reg1868 <= (&$unsigned(($signed(reg1702) ?
                          (reg1580 ?
                              reg1654 : forvar1819) : reg1710[(3'h7):(1'h0)])));
                    end
                  else
                    begin
                      reg1867 <= (+$unsigned({reg1823[(4'he):(4'hc)]}));
                      reg1868 <= $signed(reg1764);
                    end
                  reg1869 <= $unsigned($unsigned(($signed(wire1812) ?
                      $unsigned(reg1738) : reg1868)));
                  for (forvar1870 = (1'h0); (forvar1870 < (1'h0)); forvar1870 = (forvar1870 + (1'h1)))
                    begin
                      reg1871 <= ((($unsigned((8'ha1)) ~^ $unsigned(reg1595)) > (&$unsigned(reg1587))) ?
                          {reg1702[(2'h2):(1'h0)]} : $signed((reg1881 >>> reg1688)));
                    end
                end
              if ({(8'hb0)})
                begin
                  if (reg1811)
                    begin
                      reg1876 <= $signed(((reg1549[(1'h1):(1'h1)] ?
                          $signed(reg1561) : reg1743[(3'h4):(1'h1)]) ^ $signed(reg1741[(2'h3):(1'h0)])));
                      reg1877 <= $signed($signed(reg1682));
                      reg1878 <= (-{($signed(reg1841) ?
                              (reg1727 ?
                                  reg1609 : reg1551) : $signed(reg1837))});
                    end
                  else
                    begin
                      reg1876 <= reg1844[(3'h6):(3'h6)];
                      reg1877 <= (((^~(-forvar1817)) >= ($signed(reg1662) << $unsigned(reg1860))) ?
                          reg1839[(1'h0):(1'h0)] : (^reg1683));
                      reg1878 <= $unsigned(forvar1852);
                    end
                  for (forvar1879 = (1'h0); (forvar1879 < (1'h1)); forvar1879 = (forvar1879 + (1'h1)))
                    begin
                      reg1880 <= $signed(($signed($signed((8'ha4))) ?
                          reg1595 : reg1597[(1'h1):(1'h1)]));
                      reg1881 <= ($signed($unsigned({(8'ha4)})) >>> $signed((&(|wire1542))));
                    end
                end
              else
                begin
                  for (forvar1876 = (1'h0); (forvar1876 < (2'h2)); forvar1876 = (forvar1876 + (1'h1)))
                    begin
                      reg1877 <= $unsigned($unsigned(reg1836[(3'h5):(2'h3)]));
                      reg1878 <= wire1541;
                    end
                  if (reg1764[(3'h5):(1'h0)])
                    begin
                      reg1879 <= $unsigned($signed({$signed(reg1602)}));
                      reg1880 <= $unsigned((^~((forvar1821 ^ reg1788) ?
                          (reg1589 <= (8'hab)) : wire1545)));
                      reg1881 <= (((^(reg1714 & reg1871)) ?
                          ($signed((8'hb3)) & (8'h9d)) : $unsigned($unsigned(reg1742))) + (reg1729[(1'h0):(1'h0)] ?
                          (forvar1842[(4'hb):(2'h2)] ?
                              ((8'h9d) | reg1875) : $unsigned(reg1884)) : (~&$unsigned(reg1619))));
                    end
                  else
                    begin
                      reg1879 <= ($signed(({reg1658} ?
                          (reg1757 < reg1792) : $unsigned(reg1623))) < reg1626[(3'h7):(3'h4)]);
                      reg1880 <= $unsigned((($signed(reg1648) ?
                              (reg1628 - reg1884) : reg1567) ?
                          (8'ha3) : $signed($signed(reg1700))));
                      reg1881 <= (reg1626 ?
                          reg1706 : ($unsigned((reg1862 ^ forvar1870)) ?
                              ($signed((8'ha6)) ?
                                  (!forvar1842) : (forvar1866 ?
                                      reg1609 : reg1633)) : $unsigned($unsigned(forvar1866))));
                    end
                end
              reg1882 <= reg1859[(2'h3):(2'h2)];
            end
        end
      reg1885 <= $unsigned((~reg1647[(2'h3):(2'h3)]));
    end
  assign wire1886 = ((+($unsigned((8'haf)) * reg1690[(4'hf):(4'he)])) ?
                        reg1712[(3'h4):(1'h1)] : reg1645[(1'h0):(1'h0)]);
  assign wire1887 = $unsigned((~($unsigned(reg1622) & (&reg1615))));
  always
    @(posedge clk) begin
      reg1888 <= reg1622[(2'h2):(2'h2)];
      for (forvar1889 = (1'h0); (forvar1889 < (1'h1)); forvar1889 = (forvar1889 + (1'h1)))
        begin
          if ((({{(8'ha7)}} ?
              {(~|reg1610)} : $unsigned($unsigned(reg1868))) | reg1792[(3'h4):(2'h2)]))
            begin
              for (forvar1890 = (1'h0); (forvar1890 < (2'h2)); forvar1890 = (forvar1890 + (1'h1)))
                begin
                  reg1891 <= (reg1867 ?
                      $signed($unsigned((reg1780 ~^ reg1680))) : reg1857[(4'h8):(3'h7)]);
                end
            end
          else
            begin
              if (reg1869[(4'h9):(4'h8)])
                begin
                  for (forvar1890 = (1'h0); (forvar1890 < (2'h2)); forvar1890 = (forvar1890 + (1'h1)))
                    begin
                      reg1891 <= $unsigned(((reg1673 << $signed((8'ha9))) ?
                          $signed($signed(reg1767)) : wire1543[(3'h7):(1'h0)]));
                      reg1892 <= $unsigned((8'h9c));
                      reg1893 <= ((reg1860[(1'h0):(1'h0)] + (8'ha8)) ?
                          reg1832[(4'hc):(3'h7)] : (((wire1543 ?
                              reg1609 : reg1641) >= $signed((8'hae))) < $unsigned((8'h9f))));
                      reg1894 <= ($unsigned({{reg1711}}) ~^ $unsigned({reg1623[(2'h2):(1'h0)]}));
                    end
                end
              else
                begin
                  for (forvar1890 = (1'h0); (forvar1890 < (2'h2)); forvar1890 = (forvar1890 + (1'h1)))
                    begin
                      reg1891 <= {reg1826};
                      reg1892 <= reg1737;
                      reg1893 <= (^~reg1621);
                      reg1894 <= $unsigned($unsigned($unsigned((reg1853 ?
                          reg1891 : reg1581))));
                    end
                  for (forvar1895 = (1'h0); (forvar1895 < (1'h1)); forvar1895 = (forvar1895 + (1'h1)))
                    begin
                      reg1896 <= reg1843[(2'h2):(1'h0)];
                      reg1897 <= $signed((((^~(8'hb5)) ~^ reg1834[(1'h1):(1'h1)]) + $signed({reg1801})));
                      reg1898 <= $unsigned($signed(($unsigned(reg1632) ^~ $unsigned(reg1591))));
                      reg1899 <= reg1853[(1'h1):(1'h1)];
                    end
                end
              reg1900 <= ((^reg1872) ? reg1826 : $unsigned($unsigned(reg1741)));
              reg1901 <= {reg1762[(1'h1):(1'h0)]};
            end
          reg1902 <= reg1617;
          reg1903 <= reg1800[(3'h6):(2'h3)];
          reg1904 <= (~($unsigned($signed(reg1876)) ?
              (8'hb5) : reg1589[(1'h1):(1'h1)]));
        end
    end
  always
    @(posedge clk) begin
      if ($signed(reg1636[(2'h2):(2'h2)]))
        begin
          for (forvar1905 = (1'h0); (forvar1905 < (2'h2)); forvar1905 = (forvar1905 + (1'h1)))
            begin
              for (forvar1906 = (1'h0); (forvar1906 < (1'h0)); forvar1906 = (forvar1906 + (1'h1)))
                begin
                  reg1907 <= (((^$signed(reg1825)) ?
                      (8'ha7) : {$unsigned((8'ha4))}) <= (($unsigned(reg1600) ?
                          wire1544 : (reg1872 ? reg1616 : wire1886)) ?
                      reg1616 : reg1893[(1'h0):(1'h0)]));
                  if (reg1709[(4'he):(3'h4)])
                    begin
                      reg1908 <= $unsigned($signed($unsigned(reg1701)));
                      reg1909 <= (reg1693 ? $signed(reg1894) : (8'hb9));
                      reg1910 <= (reg1642 >>> $unsigned($unsigned((8'h9d))));
                    end
                  else
                    begin
                      reg1908 <= reg1910[(3'h6):(1'h0)];
                    end
                  if (reg1761[(4'h8):(3'h7)])
                    begin
                      reg1911 <= $unsigned((reg1865 ?
                          (((8'hac) ?
                              reg1607 : reg1904) << $signed(reg1661)) : reg1727));
                      reg1912 <= reg1685;
                    end
                  else
                    begin
                      reg1911 <= reg1777[(3'h5):(2'h3)];
                    end
                end
              for (forvar1913 = (1'h0); (forvar1913 < (1'h0)); forvar1913 = (forvar1913 + (1'h1)))
                begin
                  if ({{($signed(reg1614) ? (8'hb6) : reg1873)}})
                    begin
                      reg1914 <= (^$unsigned((~^reg1707[(2'h3):(1'h0)])));
                      reg1915 <= reg1671[(3'h7):(1'h1)];
                      reg1916 <= ({reg1899} >> reg1840[(3'h6):(1'h1)]);
                      reg1917 <= {({(|reg1899)} ?
                              $signed(reg1746) : $signed(reg1875))};
                    end
                  else
                    begin
                      reg1914 <= (($signed((~|reg1674)) && (reg1747[(4'hd):(1'h1)] ^~ (reg1917 && reg1878))) <= {($unsigned(reg1739) <= $unsigned(wire1546))});
                    end
                end
            end
          if (({$signed(reg1583)} & reg1792))
            begin
              if ((8'haa))
                begin
                  reg1918 <= (reg1804[(3'h4):(1'h1)] ?
                      reg1673 : ((~&$unsigned(reg1763)) ?
                          $signed($unsigned((8'ha1))) : $signed((reg1811 ?
                              reg1583 : reg1670))));
                  if (reg1850)
                    begin
                      reg1919 <= {(8'hab)};
                      reg1920 <= {(~&(+(~|reg1891)))};
                      reg1921 <= (reg1668[(2'h3):(2'h2)] ?
                          reg1596[(1'h1):(1'h0)] : reg1702[(1'h1):(1'h1)]);
                      reg1922 <= ($unsigned((~^(~&(8'haa)))) ?
                          (^(~$unsigned(reg1704))) : (|((^~reg1688) ?
                              ((8'ha7) ?
                                  reg1603 : reg1826) : (reg1807 >= reg1798))));
                    end
                  else
                    begin
                      reg1919 <= ($signed($unsigned(reg1753[(3'h4):(3'h4)])) > ((reg1857 + $unsigned(reg1720)) ~^ $unsigned((~&reg1793))));
                    end
                  for (forvar1923 = (1'h0); (forvar1923 < (2'h3)); forvar1923 = (forvar1923 + (1'h1)))
                    begin
                      reg1924 <= $signed((reg1778[(3'h6):(3'h4)] != $signed($signed(reg1788))));
                      reg1925 <= $signed($unsigned(($signed(reg1619) ?
                          ((8'ha0) ? reg1714 : (8'h9d)) : (reg1800 ?
                              reg1856 : reg1884))));
                      reg1926 <= ($unsigned($signed(reg1719)) && reg1607[(4'hd):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar1918 = (1'h0); (forvar1918 < (2'h2)); forvar1918 = (forvar1918 + (1'h1)))
                    begin
                      reg1919 <= reg1811[(2'h2):(1'h0)];
                      reg1920 <= (!$signed((8'hb4)));
                    end
                  for (forvar1921 = (1'h0); (forvar1921 < (2'h2)); forvar1921 = (forvar1921 + (1'h1)))
                    begin
                      reg1922 <= $unsigned(reg1636[(3'h4):(1'h1)]);
                      reg1923 <= $unsigned((&$unsigned((8'hb7))));
                    end
                  for (forvar1924 = (1'h0); (forvar1924 < (1'h0)); forvar1924 = (forvar1924 + (1'h1)))
                    begin
                      reg1925 <= reg1852;
                    end
                end
            end
          else
            begin
              for (forvar1918 = (1'h0); (forvar1918 < (2'h3)); forvar1918 = (forvar1918 + (1'h1)))
                begin
                  if (((reg1694 ?
                          ({reg1626} ?
                              (reg1700 ?
                                  reg1891 : (8'ha3)) : reg1865) : $unsigned($signed(reg1668))) ?
                      (8'hb5) : ((!(-(8'hb0))) ~^ (~$signed(reg1884)))))
                    begin
                      reg1919 <= reg1721[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg1919 <= (~reg1623);
                      reg1920 <= (|((~^reg1635[(4'he):(4'ha)]) ?
                          ((+reg1695) ?
                              (reg1556 & reg1596) : $signed(wire1771)) : ({forvar1913} < (reg1689 ?
                              reg1821 : (8'ha6)))));
                    end
                end
              for (forvar1921 = (1'h0); (forvar1921 < (1'h1)); forvar1921 = (forvar1921 + (1'h1)))
                begin
                  for (forvar1922 = (1'h0); (forvar1922 < (2'h2)); forvar1922 = (forvar1922 + (1'h1)))
                    begin
                      reg1923 <= $unsigned($unsigned(reg1781[(1'h1):(1'h1)]));
                      reg1924 <= $unsigned((~({reg1680} ?
                          (reg1710 ^ reg1737) : reg1661[(2'h3):(2'h3)])));
                      reg1925 <= reg1797[(3'h7):(1'h1)];
                    end
                  for (forvar1926 = (1'h0); (forvar1926 < (2'h3)); forvar1926 = (forvar1926 + (1'h1)))
                    begin
                      reg1927 <= (forvar1906[(4'h8):(1'h1)] << $signed($signed($unsigned(reg1870))));
                    end
                  for (forvar1928 = (1'h0); (forvar1928 < (2'h2)); forvar1928 = (forvar1928 + (1'h1)))
                    begin
                      reg1929 <= $signed((^(~|(~reg1654))));
                    end
                end
              if ($signed(reg1861))
                begin
                  if (($unsigned(((reg1766 + reg1658) ?
                      $signed(reg1836) : $signed(reg1756))) >> $signed(reg1730[(3'h4):(1'h0)])))
                    begin
                      reg1930 <= $unsigned($unsigned((~&(~&reg1803))));
                    end
                  else
                    begin
                      reg1930 <= $signed((|(+reg1795[(3'h5):(2'h2)])));
                      reg1931 <= reg1555;
                      reg1932 <= ((reg1631[(3'h4):(2'h2)] ?
                          ((~|reg1791) << $unsigned(reg1784)) : reg1717[(3'h5):(2'h3)]) && (8'h9d));
                    end
                  for (forvar1933 = (1'h0); (forvar1933 < (1'h0)); forvar1933 = (forvar1933 + (1'h1)))
                    begin
                      reg1934 <= (~&$unsigned(reg1663));
                      reg1935 <= (($unsigned(((8'hba) > reg1861)) ?
                          (~&$signed(reg1599)) : reg1763) != reg1646[(1'h0):(1'h0)]);
                      reg1936 <= reg1654;
                    end
                  for (forvar1937 = (1'h0); (forvar1937 < (1'h0)); forvar1937 = (forvar1937 + (1'h1)))
                    begin
                      reg1938 <= $unsigned(reg1634);
                      reg1939 <= reg1633[(2'h2):(1'h0)];
                      reg1940 <= reg1602[(2'h2):(1'h0)];
                      reg1941 <= (reg1789[(2'h3):(1'h0)] ?
                          ($unsigned($signed(reg1649)) ?
                              ({reg1626} ?
                                  reg1678 : $signed((8'hb6))) : reg1752[(2'h3):(1'h0)]) : (reg1912[(2'h3):(1'h0)] ?
                              (&(reg1556 ?
                                  reg1634 : reg1732)) : $unsigned((reg1750 || reg1852))));
                    end
                end
              else
                begin
                  if ((!reg1878))
                    begin
                      reg1930 <= reg1830;
                      reg1931 <= (reg1639[(2'h2):(1'h0)] >= {$unsigned(reg1901[(2'h3):(2'h2)])});
                    end
                  else
                    begin
                      reg1930 <= (reg1902 > (|(|(~^reg1798))));
                      reg1931 <= (&($signed(((8'ha5) ?
                          reg1738 : reg1599)) || ($unsigned(wire1771) ?
                          $signed(reg1745) : (!reg1635))));
                    end
                  for (forvar1932 = (1'h0); (forvar1932 < (1'h1)); forvar1932 = (forvar1932 + (1'h1)))
                    begin
                      reg1933 <= (~^$signed((-(reg1935 <<< (8'h9f)))));
                      reg1934 <= (-$unsigned($unsigned((-forvar1913))));
                      reg1935 <= (~^$signed((^(reg1617 ? reg1881 : (8'h9d)))));
                    end
                end
            end
          reg1942 <= {{(^~reg1724)}};
        end
      else
        begin
          for (forvar1905 = (1'h0); (forvar1905 < (1'h0)); forvar1905 = (forvar1905 + (1'h1)))
            begin
              for (forvar1906 = (1'h0); (forvar1906 < (2'h2)); forvar1906 = (forvar1906 + (1'h1)))
                begin
                  for (forvar1907 = (1'h0); (forvar1907 < (2'h3)); forvar1907 = (forvar1907 + (1'h1)))
                    begin
                      reg1908 <= $unsigned((~&reg1892[(2'h3):(1'h1)]));
                      reg1909 <= $signed($signed($signed(reg1648)));
                    end
                  if (reg1822[(1'h0):(1'h0)])
                    begin
                      reg1910 <= $signed((^~reg1827));
                      reg1911 <= (!$signed((~&reg1927[(2'h3):(1'h1)])));
                      reg1912 <= $signed(reg1941);
                    end
                  else
                    begin
                      reg1910 <= ((~|reg1736) >= {reg1807[(3'h5):(2'h3)]});
                      reg1911 <= reg1817[(4'h9):(3'h7)];
                      reg1912 <= {$unsigned(reg1759)};
                    end
                  for (forvar1913 = (1'h0); (forvar1913 < (1'h1)); forvar1913 = (forvar1913 + (1'h1)))
                    begin
                      reg1914 <= $signed(($signed($unsigned(reg1843)) || $unsigned((reg1685 != reg1835))));
                      reg1915 <= reg1834;
                    end
                end
              if ($unsigned($signed($signed($unsigned(reg1862)))))
                begin
                  reg1916 <= $unsigned({($unsigned(reg1786) == (reg1614 ?
                          reg1874 : reg1829))});
                  if ((reg1838 ?
                      reg1780 : {($signed(reg1888) ? {reg1831} : (&reg1761))}))
                    begin
                      reg1917 <= $unsigned((((reg1919 < reg1852) ?
                              $unsigned(reg1820) : (reg1837 != reg1643)) ?
                          $signed($unsigned(reg1681)) : ((~&reg1556) + reg1908[(3'h5):(1'h0)])));
                      reg1918 <= (reg1885 & (&$unsigned((!reg1807))));
                      reg1919 <= reg1926;
                    end
                  else
                    begin
                      reg1917 <= (|((reg1790[(2'h3):(2'h2)] >>> (reg1596 ?
                              reg1577 : reg1658)) ?
                          {((8'ha1) ? reg1784 : (8'hb6))} : reg1807));
                      reg1918 <= $signed(reg1693);
                    end
                  for (forvar1920 = (1'h0); (forvar1920 < (1'h0)); forvar1920 = (forvar1920 + (1'h1)))
                    begin
                      reg1921 <= {$unsigned(reg1861)};
                    end
                  for (forvar1922 = (1'h0); (forvar1922 < (1'h0)); forvar1922 = (forvar1922 + (1'h1)))
                    begin
                      reg1923 <= ($signed((+reg1801)) != reg1769[(4'h8):(1'h0)]);
                      reg1924 <= (reg1918 - $unsigned(({reg1924} ?
                          ((8'hb4) ? (8'haf) : reg1631) : (!reg1740))));
                    end
                end
              else
                begin
                  for (forvar1916 = (1'h0); (forvar1916 < (2'h2)); forvar1916 = (forvar1916 + (1'h1)))
                    begin
                      reg1917 <= (reg1823[(4'h9):(1'h1)] ?
                          $unsigned((wire1543[(4'h9):(2'h2)] ?
                              (reg1764 ? reg1864 : reg1888) : (reg1811 ?
                                  reg1634 : (8'ha2)))) : {$signed($unsigned(reg1821))});
                      reg1918 <= reg1747;
                      reg1919 <= reg1833[(4'ha):(3'h4)];
                      reg1920 <= ((($unsigned(reg1695) ?
                                  $unsigned((8'ha8)) : (8'had)) ?
                              reg1659[(1'h1):(1'h0)] : $unsigned(reg1576[(4'h9):(2'h2)])) ?
                          $signed((reg1840 ?
                              (reg1891 ?
                                  (8'h9f) : reg1933) : reg1581[(4'h9):(1'h0)])) : reg1784);
                    end
                  for (forvar1921 = (1'h0); (forvar1921 < (1'h0)); forvar1921 = (forvar1921 + (1'h1)))
                    begin
                      reg1922 <= $unsigned(((~&(+reg1717)) ?
                          (^$unsigned(forvar1937)) : ({reg1769} ?
                              (reg1774 ? reg1658 : reg1738) : {reg1567})));
                    end
                  for (forvar1923 = (1'h0); (forvar1923 < (2'h3)); forvar1923 = (forvar1923 + (1'h1)))
                    begin
                      reg1924 <= reg1873;
                      reg1925 <= (~&(^(((8'hae) ?
                          reg1808 : (8'hac)) ^ (~&reg1552))));
                      reg1926 <= {$unsigned($unsigned(reg1782[(3'h5):(3'h4)]))};
                      reg1927 <= reg1841[(3'h5):(2'h3)];
                    end
                  for (forvar1928 = (1'h0); (forvar1928 < (2'h3)); forvar1928 = (forvar1928 + (1'h1)))
                    begin
                      reg1929 <= $signed(reg1557[(3'h5):(2'h2)]);
                      reg1930 <= ((($signed(reg1721) << $signed(reg1752)) ?
                              reg1661 : reg1902[(1'h1):(1'h0)]) ?
                          ($unsigned($unsigned(reg1610)) >>> reg1567[(3'h7):(2'h2)]) : (reg1657 ^~ (reg1791 != reg1590[(1'h1):(1'h1)])));
                    end
                end
              for (forvar1931 = (1'h0); (forvar1931 < (1'h1)); forvar1931 = (forvar1931 + (1'h1)))
                begin
                  if (($unsigned(wire1543[(3'h4):(3'h4)]) ?
                      ($signed(reg1938) >> reg1596[(1'h1):(1'h1)]) : ($unsigned((^~(8'hba))) || $signed((reg1756 ?
                          reg1625 : reg1791)))))
                    begin
                      reg1932 <= $signed(reg1769);
                      reg1933 <= $unsigned(reg1774);
                      reg1934 <= (+$unsigned(reg1704[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1932 <= ($unsigned($unsigned($unsigned(wire1771))) << {((reg1597 & reg1649) - $signed(reg1625))});
                      reg1933 <= (|(reg1552[(3'h4):(3'h4)] ?
                          $signed(reg1914[(1'h1):(1'h1)]) : ($signed((8'h9e)) ?
                              $unsigned((8'ha7)) : {reg1731})));
                    end
                  if ($signed({$unsigned((^reg1806))}))
                    begin
                      reg1935 <= ($unsigned((reg1629[(4'hc):(4'hb)] ?
                          {reg1591} : (~|reg1686))) != $signed($signed((reg1576 >> reg1571))));
                      reg1936 <= reg1617;
                    end
                  else
                    begin
                      reg1935 <= ($unsigned($unsigned($unsigned(reg1864))) & ($signed(((8'hb1) ?
                              forvar1918 : reg1894)) ?
                          $unsigned(reg1718[(4'h8):(3'h7)]) : {$unsigned(reg1803)}));
                      reg1936 <= $unsigned((reg1721[(4'hd):(4'h9)] > ((reg1784 == reg1941) ?
                          (reg1821 == (8'haf)) : {reg1552})));
                      reg1937 <= (&({(~&reg1841)} < (reg1793[(3'h6):(3'h4)] ?
                          $unsigned(reg1820) : (~|reg1832))));
                      reg1938 <= ($signed(reg1749[(3'h4):(1'h1)]) ?
                          $signed(reg1794[(1'h0):(1'h0)]) : reg1580);
                    end
                  reg1939 <= reg1844;
                end
              reg1940 <= (~|$signed(reg1598[(4'h8):(2'h3)]));
            end
          if ((~|$unsigned($signed(reg1922[(3'h7):(3'h4)]))))
            begin
              for (forvar1941 = (1'h0); (forvar1941 < (2'h3)); forvar1941 = (forvar1941 + (1'h1)))
                begin
                  for (forvar1942 = (1'h0); (forvar1942 < (1'h0)); forvar1942 = (forvar1942 + (1'h1)))
                    begin
                      reg1943 <= (-reg1822[(3'h5):(1'h1)]);
                      reg1944 <= forvar1916[(3'h6):(3'h4)];
                      reg1945 <= $unsigned($signed(reg1893[(4'h8):(2'h2)]));
                    end
                  for (forvar1946 = (1'h0); (forvar1946 < (2'h2)); forvar1946 = (forvar1946 + (1'h1)))
                    begin
                      reg1947 <= $signed((($unsigned(reg1619) ?
                          (~&reg1680) : reg1598[(3'h7):(1'h1)]) || (+((8'h9f) ?
                          reg1757 : reg1649))));
                      reg1948 <= reg1749[(3'h4):(3'h4)];
                      reg1949 <= ($signed({wire1812}) ?
                          (reg1821[(4'h8):(3'h6)] ?
                              reg1558[(3'h5):(2'h3)] : (!$unsigned(reg1774))) : $unsigned(reg1775[(1'h0):(1'h0)]));
                      reg1950 <= (reg1789[(1'h0):(1'h0)] ?
                          $signed((~$signed(forvar1905))) : (&(~|$signed(reg1727))));
                    end
                  if ($signed($signed((reg1747[(2'h3):(1'h0)] ?
                      ((8'ha5) & reg1581) : (reg1654 ? reg1740 : forvar1923)))))
                    begin
                      reg1951 <= ($signed({reg1835[(2'h3):(2'h2)]}) ?
                          reg1786 : (8'hb3));
                      reg1952 <= $unsigned(reg1873);
                    end
                  else
                    begin
                      reg1951 <= {(8'ha0)};
                      reg1952 <= reg1693[(1'h1):(1'h0)];
                      reg1953 <= $signed($signed((((8'hae) | reg1833) * (reg1756 ?
                          reg1904 : (8'hba)))));
                    end
                end
              if ((reg1879 >>> $signed(reg1674)))
                begin
                  reg1954 <= $signed({$unsigned(reg1871[(4'h8):(1'h1)])});
                  if (($signed((reg1835[(1'h0):(1'h0)] ?
                      (reg1925 & reg1874) : reg1668[(2'h2):(1'h0)])) && reg1938))
                    begin
                      reg1955 <= (&(^~(~|{forvar1923})));
                      reg1956 <= reg1603;
                      reg1957 <= (^~$signed((reg1591[(4'hc):(4'hb)] <= (reg1798 ?
                          reg1924 : reg1741))));
                    end
                  else
                    begin
                      reg1955 <= (wire1887 <<< reg1931);
                      reg1956 <= reg1790[(2'h2):(1'h0)];
                    end
                  for (forvar1958 = (1'h0); (forvar1958 < (1'h1)); forvar1958 = (forvar1958 + (1'h1)))
                    begin
                      reg1959 <= $unsigned(({(-reg1925)} ?
                          reg1957[(3'h5):(3'h5)] : {(reg1635 << reg1931)}));
                      reg1960 <= $signed((~&(&$signed(reg1808))));
                    end
                end
              else
                begin
                  for (forvar1954 = (1'h0); (forvar1954 < (2'h3)); forvar1954 = (forvar1954 + (1'h1)))
                    begin
                      reg1955 <= (&$signed($unsigned((reg1657 - reg1591))));
                      reg1956 <= reg1622[(1'h1):(1'h1)];
                    end
                  reg1957 <= $unsigned(($unsigned((~(8'haa))) <<< ({reg1607} || reg1904[(3'h4):(2'h2)])));
                  for (forvar1958 = (1'h0); (forvar1958 < (1'h0)); forvar1958 = (forvar1958 + (1'h1)))
                    begin
                      reg1959 <= (^~($unsigned({reg1614}) <<< reg1644[(2'h2):(1'h0)]));
                      reg1960 <= reg1773[(3'h4):(2'h3)];
                      reg1961 <= reg1862[(2'h3):(1'h0)];
                    end
                  for (forvar1962 = (1'h0); (forvar1962 < (1'h0)); forvar1962 = (forvar1962 + (1'h1)))
                    begin
                      reg1963 <= (8'h9d);
                      reg1964 <= reg1714[(3'h6):(1'h0)];
                    end
                end
            end
          else
            begin
              if ((reg1932[(3'h5):(3'h4)] ?
                  (!reg1922[(2'h2):(1'h0)]) : $signed({(reg1830 >> reg1617)})))
                begin
                  for (forvar1941 = (1'h0); (forvar1941 < (1'h1)); forvar1941 = (forvar1941 + (1'h1)))
                    begin
                      reg1942 <= (!wire1815);
                      reg1943 <= (reg1662 > reg1804);
                      reg1944 <= ($unsigned(((reg1757 ? reg1930 : reg1788) ?
                              $unsigned(reg1617) : reg1557)) ?
                          ((reg1855[(1'h1):(1'h1)] < reg1937[(1'h1):(1'h1)]) ?
                              reg1571[(2'h3):(2'h2)] : reg1891[(3'h6):(2'h2)]) : (reg1710 ?
                              {$signed(reg1956)} : ((reg1849 ?
                                  reg1700 : (8'hb8)) << $unsigned(reg1747))));
                      reg1945 <= {(({reg1934} ? reg1707 : reg1783) ?
                              ($unsigned(reg1599) ?
                                  {reg1947} : (reg1576 != reg1563)) : wire1813[(3'h6):(3'h6)])};
                    end
                  if ((8'hb3))
                    begin
                      reg1946 <= {({$signed(reg1918)} >>> (~^$unsigned((8'hb6))))};
                      reg1947 <= (~((forvar1937[(1'h0):(1'h0)] ?
                          reg1549[(1'h0):(1'h0)] : $signed(reg1869)) > $signed(reg1877)));
                      reg1948 <= ((8'hac) ?
                          {$unsigned(reg1549[(2'h2):(1'h0)])} : reg1803);
                      reg1949 <= reg1841;
                    end
                  else
                    begin
                      reg1946 <= (^~$unsigned(reg1615));
                      reg1947 <= $unsigned($unsigned(reg1783[(2'h3):(2'h3)]));
                      reg1948 <= (+(8'hba));
                    end
                end
              else
                begin
                  for (forvar1941 = (1'h0); (forvar1941 < (1'h0)); forvar1941 = (forvar1941 + (1'h1)))
                    begin
                      reg1942 <= reg1791[(1'h0):(1'h0)];
                    end
                end
              for (forvar1950 = (1'h0); (forvar1950 < (2'h2)); forvar1950 = (forvar1950 + (1'h1)))
                begin
                  for (forvar1951 = (1'h0); (forvar1951 < (2'h2)); forvar1951 = (forvar1951 + (1'h1)))
                    begin
                      reg1952 <= forvar1913;
                    end
                  if ((((+(reg1912 ? forvar1926 : reg1949)) ?
                          reg1790[(2'h3):(2'h3)] : reg1830[(3'h4):(2'h2)]) ?
                      reg1563 : $signed(($unsigned(reg1876) || {reg1846}))))
                    begin
                      reg1953 <= $unsigned($signed(reg1909));
                      reg1954 <= reg1914;
                      reg1955 <= $unsigned({((wire1814 ?
                              reg1673 : (8'hac)) || (reg1912 | reg1685))});
                      reg1956 <= wire1814[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg1953 <= $signed($signed(((+reg1851) || (reg1854 ?
                          reg1841 : reg1862))));
                      reg1954 <= {(8'hb2)};
                      reg1955 <= (reg1570 ?
                          reg1922[(3'h7):(1'h1)] : ($unsigned((~^(8'ha6))) ^ (~&((8'ha4) ?
                              reg1753 : reg1628))));
                    end
                  for (forvar1957 = (1'h0); (forvar1957 < (2'h2)); forvar1957 = (forvar1957 + (1'h1)))
                    begin
                      reg1958 <= $unsigned(reg1911);
                      reg1959 <= (reg1668 * $unsigned(reg1764[(4'hb):(3'h5)]));
                      reg1960 <= reg1924;
                      reg1961 <= (+(~((reg1686 ?
                          reg1831 : reg1784) && reg1711[(3'h4):(2'h3)])));
                    end
                  for (forvar1962 = (1'h0); (forvar1962 < (2'h2)); forvar1962 = (forvar1962 + (1'h1)))
                    begin
                      reg1963 <= (reg1957[(1'h0):(1'h0)] ^ $signed({$unsigned((8'hb7))}));
                    end
                end
              if (((reg1774 ?
                  ($signed(reg1773) ?
                      wire1541[(1'h0):(1'h0)] : (reg1857 ?
                          (8'ha1) : reg1951)) : $unsigned($unsigned(reg1925))) ^ {(~(reg1591 ?
                      reg1651 : reg1854))}))
                begin
                  if ($signed({$unsigned({reg1785})}))
                    begin
                      reg1964 <= $unsigned($signed(reg1803[(1'h0):(1'h0)]));
                      reg1965 <= reg1625;
                      reg1966 <= $signed((8'haa));
                      reg1967 <= {$signed(reg1780)};
                    end
                  else
                    begin
                      reg1964 <= reg1670;
                      reg1965 <= ((forvar1962 ^ ($signed(reg1904) || {reg1868})) ?
                          $signed($signed((reg1779 ?
                              wire1541 : reg1670))) : reg1818[(4'hb):(1'h0)]);
                      reg1966 <= $unsigned((((reg1717 ? reg1791 : (8'hab)) ?
                              ((8'had) ? reg1802 : (8'ha0)) : reg1868) ?
                          {(8'hb9)} : (~^((8'ha3) >= reg1958))));
                    end
                  for (forvar1968 = (1'h0); (forvar1968 < (1'h0)); forvar1968 = (forvar1968 + (1'h1)))
                    begin
                      reg1969 <= (forvar1931 <= (reg1766[(1'h0):(1'h0)] ?
                          reg1593 : reg1600));
                      reg1970 <= reg1635[(4'h9):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar1964 = (1'h0); (forvar1964 < (2'h3)); forvar1964 = (forvar1964 + (1'h1)))
                    begin
                      reg1965 <= $unsigned($unsigned((8'ha6)));
                      reg1966 <= reg1834[(2'h2):(2'h2)];
                      reg1967 <= (reg1634 ?
                          $unsigned({$unsigned(wire1541)}) : forvar1942);
                      reg1968 <= ((8'hb6) ~^ reg1786[(1'h0):(1'h0)]);
                    end
                  if ($unsigned($unsigned($signed(reg1587))))
                    begin
                      reg1969 <= reg1673;
                      reg1970 <= reg1882[(3'h7):(3'h5)];
                      reg1971 <= reg1759;
                      reg1972 <= reg1801[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1969 <= ((&reg1806[(3'h5):(2'h2)]) && ($signed(reg1642) & {{(8'h9c)}}));
                      reg1970 <= $signed($unsigned($unsigned({(8'hb4)})));
                      reg1971 <= reg1931[(1'h1):(1'h0)];
                    end
                  for (forvar1973 = (1'h0); (forvar1973 < (1'h0)); forvar1973 = (forvar1973 + (1'h1)))
                    begin
                      reg1974 <= $signed((+reg1597[(3'h7):(3'h6)]));
                      reg1975 <= {$signed($signed(reg1750[(2'h2):(1'h1)]))};
                    end
                  reg1976 <= reg1738[(2'h2):(1'h0)];
                end
            end
          reg1977 <= {$signed((8'hb2))};
          if ($unsigned(reg1623))
            begin
              reg1978 <= (($signed(reg1831) ^ (reg1801 ?
                  $unsigned(reg1829) : (reg1581 == (8'ha8)))) >>> reg1837[(2'h2):(1'h0)]);
              reg1979 <= reg1768;
              for (forvar1980 = (1'h0); (forvar1980 < (2'h3)); forvar1980 = (forvar1980 + (1'h1)))
                begin
                  for (forvar1981 = (1'h0); (forvar1981 < (1'h0)); forvar1981 = (forvar1981 + (1'h1)))
                    begin
                      reg1982 <= (+$unsigned(((reg1732 ^ reg1916) == $unsigned(reg1606))));
                    end
                end
            end
          else
            begin
              for (forvar1978 = (1'h0); (forvar1978 < (2'h3)); forvar1978 = (forvar1978 + (1'h1)))
                begin
                  for (forvar1979 = (1'h0); (forvar1979 < (2'h3)); forvar1979 = (forvar1979 + (1'h1)))
                    begin
                      reg1980 <= reg1907;
                      reg1981 <= $unsigned(reg1601);
                    end
                  for (forvar1982 = (1'h0); (forvar1982 < (2'h3)); forvar1982 = (forvar1982 + (1'h1)))
                    begin
                      reg1983 <= $signed(reg1555[(2'h3):(2'h2)]);
                      reg1984 <= reg1840[(4'ha):(3'h6)];
                      reg1985 <= reg1917[(1'h0):(1'h0)];
                    end
                  for (forvar1986 = (1'h0); (forvar1986 < (1'h0)); forvar1986 = (forvar1986 + (1'h1)))
                    begin
                      reg1987 <= (+reg1631[(1'h0):(1'h0)]);
                      reg1988 <= reg1573[(4'h9):(3'h6)];
                      reg1989 <= $unsigned($signed($signed(reg1980[(3'h6):(3'h4)])));
                      reg1990 <= (^($signed((reg1894 ?
                          reg1871 : forvar1922)) > $signed($unsigned((8'had)))));
                    end
                  for (forvar1991 = (1'h0); (forvar1991 < (1'h1)); forvar1991 = (forvar1991 + (1'h1)))
                    begin
                      reg1992 <= ($unsigned(reg1908) ?
                          ($unsigned((reg1828 >= reg1924)) ~^ $signed((~|reg1574))) : $unsigned((~&(wire1541 ?
                              (8'hab) : (8'hb2)))));
                      reg1993 <= ($unsigned($unsigned(reg1982[(4'h8):(2'h3)])) ?
                          {{$signed(reg1591)}} : reg1822);
                      reg1994 <= (~^{$signed($unsigned(forvar1941))});
                      reg1995 <= $signed((|(~^$unsigned(reg1866))));
                    end
                end
              for (forvar1996 = (1'h0); (forvar1996 < (1'h0)); forvar1996 = (forvar1996 + (1'h1)))
                begin
                  reg1997 <= $signed((($signed(reg1762) ?
                          {reg1716} : (reg1584 ~^ reg1942)) ?
                      (!(~reg1582)) : {$signed(reg1745)}));
                  reg1998 <= $signed(($signed($signed(reg1779)) ?
                      reg1980[(1'h0):(1'h0)] : (~|reg1865)));
                end
              if (reg1696[(3'h4):(1'h1)])
                begin
                  if ($signed(reg1799))
                    begin
                      reg1999 <= reg1746[(1'h0):(1'h0)];
                      reg2000 <= (!($unsigned((8'ha4)) ?
                          (((8'ha0) ?
                              reg1883 : reg1617) >> $unsigned((8'h9f))) : {(+wire1815)}));
                    end
                  else
                    begin
                      reg1999 <= {(^$signed($signed(reg1669)))};
                      reg2000 <= $signed(reg1691[(1'h0):(1'h0)]);
                      reg2001 <= reg1653[(3'h5):(2'h3)];
                      reg2002 <= reg1758[(4'h8):(3'h7)];
                    end
                  reg2003 <= ($signed(reg1678[(4'h8):(2'h2)]) ?
                      reg1975[(1'h1):(1'h0)] : (((~reg1612) ?
                          $unsigned((8'hb7)) : $unsigned((8'h9f))) << reg1551[(1'h1):(1'h1)]));
                end
              else
                begin
                  if ($unsigned($signed($signed(wire1815[(4'ha):(2'h2)]))))
                    begin
                      reg1999 <= (~|{(~|reg1881)});
                      reg2000 <= reg1640[(2'h2):(2'h2)];
                      reg2001 <= {forvar1951[(2'h2):(2'h2)]};
                      reg2002 <= $signed((^~(|(reg1990 ? (8'ha2) : reg1879))));
                    end
                  else
                    begin
                      reg1999 <= ($signed(($unsigned(reg1971) >> forvar1957[(3'h6):(2'h2)])) ?
                          {(reg1689 ?
                                  (8'hb8) : (&reg1938))} : {({reg1767} ~^ $unsigned(reg1736))});
                      reg2000 <= reg1963;
                    end
                  for (forvar2003 = (1'h0); (forvar2003 < (1'h1)); forvar2003 = (forvar2003 + (1'h1)))
                    begin
                      reg2004 <= (({$signed(reg1610)} ?
                          $signed(reg1643) : (8'h9d)) ~^ (&(reg1800[(2'h3):(1'h0)] ?
                          (-forvar1931) : forvar1946)));
                    end
                  if ({$signed((((8'hb5) ? reg1879 : reg1804) || ((8'hb1) ?
                          reg1948 : reg1874)))})
                    begin
                      reg2005 <= $unsigned(reg1780[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2005 <= reg1699;
                      reg2006 <= $unsigned({$signed((^reg1634))});
                      reg2007 <= reg1712;
                    end
                  for (forvar2008 = (1'h0); (forvar2008 < (1'h1)); forvar2008 = (forvar2008 + (1'h1)))
                    begin
                      reg2009 <= ((+forvar1964) ?
                          ($unsigned({reg1554}) != forvar1981) : ((forvar1928[(4'h9):(2'h3)] < reg1883[(3'h4):(1'h0)]) ?
                              reg1840 : $unsigned({reg1577})));
                      reg2010 <= $unsigned($unsigned(reg1882));
                      reg2011 <= ({$signed(reg1792)} ?
                          $signed($unsigned($signed(reg1908))) : reg1554[(4'h8):(4'h8)]);
                      reg2012 <= (^(~$unsigned(reg1963[(2'h2):(2'h2)])));
                    end
                end
              for (forvar2013 = (1'h0); (forvar2013 < (2'h2)); forvar2013 = (forvar2013 + (1'h1)))
                begin
                  for (forvar2014 = (1'h0); (forvar2014 < (2'h2)); forvar2014 = (forvar2014 + (1'h1)))
                    begin
                      reg2015 <= reg1652;
                      reg2016 <= (!reg1597);
                      reg2017 <= $unsigned(($unsigned(reg1673[(3'h7):(2'h3)]) << (-{reg1615})));
                    end
                  for (forvar2018 = (1'h0); (forvar2018 < (1'h1)); forvar2018 = (forvar2018 + (1'h1)))
                    begin
                      reg2019 <= ((&($signed(reg1561) ?
                          ((8'ha7) ?
                              forvar1958 : reg1737) : reg1938)) & (!$signed(((8'ha2) ?
                          reg1853 : reg1821))));
                      reg2020 <= {reg1762};
                    end
                  for (forvar2021 = (1'h0); (forvar2021 < (2'h3)); forvar2021 = (forvar2021 + (1'h1)))
                    begin
                      reg2022 <= wire1813;
                      reg2023 <= (((^~(reg1794 > reg1714)) * reg1830[(4'h9):(1'h1)]) - ($signed((!reg1663)) ?
                          {reg1640} : ($signed((8'hb6)) >= (reg1700 + reg1966))));
                      reg2024 <= ($signed(forvar2008[(4'he):(4'hb)]) >> (8'hb7));
                    end
                end
            end
        end
    end
  assign wire2025 = reg1717;
  assign wire2026 = (|((-reg1711[(3'h5):(3'h5)]) ?
                        (((8'ha8) ?
                            (8'hab) : reg1563) <= {(8'hae)}) : reg1791[(1'h1):(1'h1)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3901
#(parameter param4718 = (((((8'h9f) == (8'hb2)) ? ((8'hb3) | (8'hb8)) : (|(8'hac))) == (|((8'ha4) ? (8'hb6) : (8'ha4)))) ? ((|(~&(8'h9e))) ? (((8'ha6) ? (8'had) : (8'h9f)) ? (!(8'hb9)) : ((8'ha9) + (8'ha1))) : (&((8'h9d) ? (8'ha1) : (8'hb9)))) : ({((8'hb6) >>> (8'hb7))} ? (8'hb9) : ((!(8'hab)) > (8'hb9)))))
(y, clk, wire3902, wire3903, wire3904, wire3905, wire3906);
  output wire [(32'h8dd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire3902;
  input wire [(3'h6):(1'h0)] wire3903;
  input wire [(2'h3):(1'h0)] wire3904;
  input wire [(4'hb):(1'h0)] wire3905;
  input wire [(4'h9):(1'h0)] wire3906;
  wire signed [(4'hf):(1'h0)] wire4584;
  wire [(4'h8):(1'h0)] wire4583;
  wire [(4'hd):(1'h0)] wire4545;
  wire [(4'h9):(1'h0)] wire4544;
  wire signed [(4'h8):(1'h0)] wire4543;
  wire signed [(4'ha):(1'h0)] wire4542;
  wire [(3'h5):(1'h0)] wire4541;
  wire [(3'h7):(1'h0)] wire3907;
  wire signed [(5'h10):(1'h0)] wire3908;
  wire signed [(2'h2):(1'h0)] wire3932;
  wire [(4'hb):(1'h0)] wire3933;
  wire signed [(4'hc):(1'h0)] wire3934;
  wire signed [(4'ha):(1'h0)] wire3935;
  wire signed [(4'h8):(1'h0)] wire4539;
  reg [(4'hf):(1'h0)] reg4717 = (1'h0);
  reg [(4'hf):(1'h0)] reg4715 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4714 = (1'h0);
  reg [(4'he):(1'h0)] reg4713 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4712 = (1'h0);
  reg [(3'h5):(1'h0)] reg4711 = (1'h0);
  reg [(4'hf):(1'h0)] reg4710 = (1'h0);
  reg [(4'hc):(1'h0)] reg4709 = (1'h0);
  reg [(4'ha):(1'h0)] reg4708 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4707 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4706 = (1'h0);
  reg [(3'h4):(1'h0)] reg4694 = (1'h0);
  reg [(2'h2):(1'h0)] reg4705 = (1'h0);
  reg [(3'h7):(1'h0)] reg4704 = (1'h0);
  reg [(4'ha):(1'h0)] reg4703 = (1'h0);
  reg [(4'hc):(1'h0)] reg4702 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4695 = (1'h0);
  reg [(3'h4):(1'h0)] reg4687 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4684 = (1'h0);
  reg [(4'ha):(1'h0)] reg4683 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4678 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4701 = (1'h0);
  reg [(4'hc):(1'h0)] reg4700 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4699 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4698 = (1'h0);
  reg [(3'h7):(1'h0)] reg4697 = (1'h0);
  reg [(4'hf):(1'h0)] reg4696 = (1'h0);
  reg [(3'h6):(1'h0)] reg4692 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4665 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4691 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4690 = (1'h0);
  reg [(3'h7):(1'h0)] reg4689 = (1'h0);
  reg [(4'hb):(1'h0)] reg4688 = (1'h0);
  reg [(3'h6):(1'h0)] reg4686 = (1'h0);
  reg [(4'ha):(1'h0)] reg4685 = (1'h0);
  reg [(4'hb):(1'h0)] reg4682 = (1'h0);
  reg [(3'h5):(1'h0)] reg4681 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4680 = (1'h0);
  reg [(3'h7):(1'h0)] reg4679 = (1'h0);
  reg [(3'h6):(1'h0)] reg4677 = (1'h0);
  reg [(4'hc):(1'h0)] reg4676 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4675 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4674 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4673 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4672 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4671 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4670 = (1'h0);
  reg [(2'h2):(1'h0)] reg4669 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4668 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4667 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4666 = (1'h0);
  reg [(2'h3):(1'h0)] reg4664 = (1'h0);
  reg [(4'hb):(1'h0)] reg4663 = (1'h0);
  reg [(4'he):(1'h0)] reg4662 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4661 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4660 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4659 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4658 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4651 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4649 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4657 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4656 = (1'h0);
  reg [(5'h10):(1'h0)] reg4655 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4654 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4653 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4652 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4650 = (1'h0);
  reg [(2'h2):(1'h0)] reg4648 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4646 = (1'h0);
  reg [(5'h10):(1'h0)] reg4645 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4644 = (1'h0);
  reg [(4'hd):(1'h0)] reg4643 = (1'h0);
  reg [(2'h3):(1'h0)] reg4641 = (1'h0);
  reg [(2'h3):(1'h0)] reg4640 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4639 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4638 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4637 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4636 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4635 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4634 = (1'h0);
  reg [(4'he):(1'h0)] reg4622 = (1'h0);
  reg [(2'h2):(1'h0)] reg4619 = (1'h0);
  reg [(3'h7):(1'h0)] reg4631 = (1'h0);
  reg [(4'h8):(1'h0)] reg4630 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4629 = (1'h0);
  reg [(4'ha):(1'h0)] reg4628 = (1'h0);
  reg [(4'h9):(1'h0)] reg4626 = (1'h0);
  reg [(4'hb):(1'h0)] reg4625 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4624 = (1'h0);
  reg [(5'h10):(1'h0)] reg4623 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4621 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4620 = (1'h0);
  reg [(4'hc):(1'h0)] reg4618 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4617 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4616 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4615 = (1'h0);
  reg [(4'ha):(1'h0)] reg4614 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4613 = (1'h0);
  reg [(3'h4):(1'h0)] reg4612 = (1'h0);
  reg [(5'h10):(1'h0)] reg4611 = (1'h0);
  reg [(5'h10):(1'h0)] reg4610 = (1'h0);
  reg [(4'he):(1'h0)] reg4609 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4608 = (1'h0);
  reg [(4'hf):(1'h0)] reg4607 = (1'h0);
  reg [(3'h5):(1'h0)] reg4604 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4602 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4601 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4600 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4599 = (1'h0);
  reg [(4'hb):(1'h0)] reg4598 = (1'h0);
  reg [(2'h3):(1'h0)] reg4597 = (1'h0);
  reg [(2'h2):(1'h0)] reg4596 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4594 = (1'h0);
  reg [(4'hb):(1'h0)] reg4593 = (1'h0);
  reg [(4'hd):(1'h0)] reg4592 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4591 = (1'h0);
  reg [(3'h4):(1'h0)] reg4590 = (1'h0);
  reg [(4'hf):(1'h0)] reg4585 = (1'h0);
  reg [(4'hc):(1'h0)] reg4582 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4565 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4574 = (1'h0);
  reg [(4'hc):(1'h0)] reg4571 = (1'h0);
  reg [(2'h2):(1'h0)] reg4581 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4580 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4579 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4578 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4577 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4576 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4575 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4573 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4572 = (1'h0);
  reg [(4'ha):(1'h0)] reg4570 = (1'h0);
  reg [(2'h3):(1'h0)] reg4569 = (1'h0);
  reg [(3'h7):(1'h0)] reg4568 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4567 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4566 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4564 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4563 = (1'h0);
  reg [(5'h10):(1'h0)] reg4547 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4548 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4561 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4560 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4559 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4558 = (1'h0);
  reg [(4'hf):(1'h0)] reg4556 = (1'h0);
  reg [(2'h3):(1'h0)] reg4555 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4554 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4553 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4552 = (1'h0);
  reg [(5'h10):(1'h0)] reg4551 = (1'h0);
  reg [(4'hb):(1'h0)] reg4550 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4549 = (1'h0);
  reg [(4'he):(1'h0)] reg4546 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3931 = (1'h0);
  reg [(3'h6):(1'h0)] reg3930 = (1'h0);
  reg [(4'ha):(1'h0)] reg3929 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3928 = (1'h0);
  reg [(4'h9):(1'h0)] reg3927 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3926 = (1'h0);
  reg [(2'h2):(1'h0)] reg3910 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3923 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3922 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3921 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3920 = (1'h0);
  reg [(4'hf):(1'h0)] reg3919 = (1'h0);
  reg [(4'hd):(1'h0)] reg3918 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3917 = (1'h0);
  reg [(2'h3):(1'h0)] reg3916 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3914 = (1'h0);
  reg [(3'h4):(1'h0)] reg3913 = (1'h0);
  reg [(4'ha):(1'h0)] reg3911 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4716 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4700 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4690 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4685 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4682 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4677 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4672 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4671 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4670 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4662 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4695 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4694 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4693 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4667 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4666 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4656 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4652 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4687 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4684 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4683 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4678 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4669 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4665 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4650 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4651 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4649 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4647 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4642 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4634 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4633 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4632 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4621 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4627 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4622 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4619 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4606 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4605 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4603 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4595 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4589 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4588 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4587 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4586 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4569 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4564 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4577 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4574 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4571 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4565 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4562 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4553 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4550 = (1'h0);
  reg [(4'he):(1'h0)] forvar4546 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4557 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4548 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4547 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3925 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3924 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3915 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3912 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3910 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3909 = (1'h0);
  assign y = {wire4584,
                 wire4583,
                 wire4545,
                 wire4544,
                 wire4543,
                 wire4542,
                 wire4541,
                 wire3907,
                 wire3908,
                 wire3932,
                 wire3933,
                 wire3934,
                 wire3935,
                 wire4539,
                 reg4717,
                 reg4715,
                 reg4714,
                 reg4713,
                 reg4712,
                 reg4711,
                 reg4710,
                 reg4709,
                 reg4708,
                 reg4707,
                 reg4706,
                 reg4694,
                 reg4705,
                 reg4704,
                 reg4703,
                 reg4702,
                 reg4695,
                 reg4687,
                 reg4684,
                 reg4683,
                 reg4678,
                 reg4701,
                 reg4700,
                 reg4699,
                 reg4698,
                 reg4697,
                 reg4696,
                 reg4692,
                 reg4665,
                 reg4691,
                 reg4690,
                 reg4689,
                 reg4688,
                 reg4686,
                 reg4685,
                 reg4682,
                 reg4681,
                 reg4680,
                 reg4679,
                 reg4677,
                 reg4676,
                 reg4675,
                 reg4674,
                 reg4673,
                 reg4672,
                 reg4671,
                 reg4670,
                 reg4669,
                 reg4668,
                 reg4667,
                 reg4666,
                 reg4664,
                 reg4663,
                 reg4662,
                 reg4661,
                 reg4660,
                 reg4659,
                 reg4658,
                 reg4651,
                 reg4649,
                 reg4657,
                 reg4656,
                 reg4655,
                 reg4654,
                 reg4653,
                 reg4652,
                 reg4650,
                 reg4648,
                 reg4646,
                 reg4645,
                 reg4644,
                 reg4643,
                 reg4641,
                 reg4640,
                 reg4639,
                 reg4638,
                 reg4637,
                 reg4636,
                 reg4635,
                 reg4634,
                 reg4622,
                 reg4619,
                 reg4631,
                 reg4630,
                 reg4629,
                 reg4628,
                 reg4626,
                 reg4625,
                 reg4624,
                 reg4623,
                 reg4621,
                 reg4620,
                 reg4618,
                 reg4617,
                 reg4616,
                 reg4615,
                 reg4614,
                 reg4613,
                 reg4612,
                 reg4611,
                 reg4610,
                 reg4609,
                 reg4608,
                 reg4607,
                 reg4604,
                 reg4602,
                 reg4601,
                 reg4600,
                 reg4599,
                 reg4598,
                 reg4597,
                 reg4596,
                 reg4594,
                 reg4593,
                 reg4592,
                 reg4591,
                 reg4590,
                 reg4585,
                 reg4582,
                 reg4565,
                 reg4574,
                 reg4571,
                 reg4581,
                 reg4580,
                 reg4579,
                 reg4578,
                 reg4577,
                 reg4576,
                 reg4575,
                 reg4573,
                 reg4572,
                 reg4570,
                 reg4569,
                 reg4568,
                 reg4567,
                 reg4566,
                 reg4564,
                 reg4563,
                 reg4547,
                 reg4548,
                 reg4561,
                 reg4560,
                 reg4559,
                 reg4558,
                 reg4556,
                 reg4555,
                 reg4554,
                 reg4553,
                 reg4552,
                 reg4551,
                 reg4550,
                 reg4549,
                 reg4546,
                 reg3931,
                 reg3930,
                 reg3929,
                 reg3928,
                 reg3927,
                 reg3926,
                 reg3910,
                 reg3923,
                 reg3922,
                 reg3921,
                 reg3920,
                 reg3919,
                 reg3918,
                 reg3917,
                 reg3916,
                 reg3914,
                 reg3913,
                 reg3911,
                 forvar4716,
                 forvar4700,
                 forvar4690,
                 forvar4685,
                 forvar4682,
                 forvar4677,
                 forvar4672,
                 forvar4671,
                 forvar4670,
                 forvar4662,
                 forvar4695,
                 forvar4694,
                 forvar4693,
                 forvar4667,
                 forvar4666,
                 forvar4656,
                 forvar4652,
                 forvar4687,
                 forvar4684,
                 forvar4683,
                 forvar4678,
                 forvar4669,
                 forvar4665,
                 forvar4650,
                 forvar4651,
                 forvar4649,
                 forvar4647,
                 forvar4642,
                 forvar4634,
                 forvar4633,
                 forvar4632,
                 forvar4621,
                 forvar4627,
                 forvar4622,
                 forvar4619,
                 forvar4606,
                 forvar4605,
                 forvar4603,
                 forvar4595,
                 forvar4589,
                 forvar4588,
                 forvar4587,
                 forvar4586,
                 forvar4569,
                 forvar4564,
                 forvar4577,
                 forvar4574,
                 forvar4571,
                 forvar4565,
                 forvar4562,
                 forvar4553,
                 forvar4550,
                 forvar4546,
                 forvar4557,
                 forvar4548,
                 forvar4547,
                 forvar3925,
                 forvar3924,
                 forvar3915,
                 forvar3912,
                 forvar3910,
                 forvar3909,
                 (1'h0)};
  assign wire3907 = {wire3903[(2'h3):(2'h3)]};
  assign wire3908 = $signed((wire3906 ? (&wire3904) : (|(8'haf))));
  always
    @(posedge clk) begin
      for (forvar3909 = (1'h0); (forvar3909 < (1'h1)); forvar3909 = (forvar3909 + (1'h1)))
        begin
          if (wire3905)
            begin
              for (forvar3910 = (1'h0); (forvar3910 < (1'h1)); forvar3910 = (forvar3910 + (1'h1)))
                begin
                  reg3911 <= $unsigned($signed($signed((~&wire3903))));
                  for (forvar3912 = (1'h0); (forvar3912 < (1'h1)); forvar3912 = (forvar3912 + (1'h1)))
                    begin
                      reg3913 <= $signed($unsigned($unsigned({wire3903})));
                      reg3914 <= $signed($unsigned(({wire3904} != $unsigned(wire3905))));
                    end
                end
              for (forvar3915 = (1'h0); (forvar3915 < (2'h2)); forvar3915 = (forvar3915 + (1'h1)))
                begin
                  reg3916 <= (|{reg3911});
                  if ((&($unsigned((forvar3912 * forvar3910)) ?
                      $signed($unsigned(wire3906)) : ((wire3903 ?
                          wire3908 : reg3916) + $unsigned(reg3911)))))
                    begin
                      reg3917 <= ((~|(~&$signed(wire3907))) << (($signed(wire3908) ?
                          (forvar3915 != wire3903) : $unsigned(wire3908)) ~^ (+(forvar3912 ?
                          wire3906 : wire3908))));
                      reg3918 <= wire3902[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg3917 <= reg3913;
                      reg3918 <= (((~{forvar3910}) << forvar3915) && reg3914);
                      reg3919 <= ($signed((8'hb0)) ?
                          $signed(reg3911[(1'h0):(1'h0)]) : $signed((8'hba)));
                    end
                  if ((^~(wire3906 || ({reg3919} ?
                      (&forvar3909) : $signed(wire3904)))))
                    begin
                      reg3920 <= ($signed(reg3911[(2'h2):(2'h2)]) ?
                          ((wire3908 << (reg3919 != (8'hae))) & $unsigned((reg3916 ?
                              wire3902 : wire3903))) : $unsigned((8'ha9)));
                      reg3921 <= ($signed(((reg3917 && forvar3915) ?
                              (reg3913 ?
                                  forvar3912 : reg3916) : {forvar3912})) ?
                          (reg3919 ?
                              forvar3915 : $unsigned((wire3906 ?
                                  forvar3912 : wire3907))) : ({{reg3920}} >= reg3919));
                      reg3922 <= ((($signed(forvar3912) >>> $signed(wire3906)) ^~ (~|$unsigned(wire3908))) ?
                          ((^$unsigned(reg3914)) ^ $unsigned(reg3921)) : (8'hb1));
                      reg3923 <= (-(reg3921[(3'h5):(3'h4)] != ((reg3911 ?
                          reg3917 : wire3905) >>> $unsigned(wire3906))));
                    end
                  else
                    begin
                      reg3920 <= {wire3904[(1'h0):(1'h0)]};
                    end
                end
            end
          else
            begin
              reg3910 <= ((~(~&{(8'haa)})) & $unsigned({$unsigned(wire3907)}));
            end
          for (forvar3924 = (1'h0); (forvar3924 < (2'h2)); forvar3924 = (forvar3924 + (1'h1)))
            begin
              for (forvar3925 = (1'h0); (forvar3925 < (1'h0)); forvar3925 = (forvar3925 + (1'h1)))
                begin
                  if ({$signed((~|(reg3920 ? wire3902 : (8'h9c))))})
                    begin
                      reg3926 <= $signed(({(|wire3908)} ?
                          ((~&reg3914) ?
                              $unsigned(reg3917) : (^reg3916)) : (((8'ha0) - reg3918) + wire3906[(2'h2):(1'h1)])));
                      reg3927 <= (+$signed($unsigned((reg3919 ?
                          wire3906 : wire3903))));
                    end
                  else
                    begin
                      reg3926 <= ({wire3907} >= reg3910);
                      reg3927 <= (&$unsigned((reg3918 ?
                          {wire3905} : (-reg3910))));
                      reg3928 <= $unsigned(reg3918[(4'ha):(1'h0)]);
                      reg3929 <= wire3904;
                    end
                  if ((^~forvar3912))
                    begin
                      reg3930 <= $signed(((!$signed(reg3914)) ?
                          {reg3911} : (~$signed(wire3903))));
                    end
                  else
                    begin
                      reg3930 <= (forvar3915[(2'h3):(2'h2)] ?
                          $signed(($signed(reg3911) != $signed(reg3930))) : (({forvar3912} > (reg3916 ?
                                  (8'h9f) : reg3910)) ?
                              $signed({reg3927}) : reg3917[(3'h4):(3'h4)]));
                      reg3931 <= reg3913[(1'h0):(1'h0)];
                    end
                end
            end
        end
    end
  assign wire3932 = wire3908;
  assign wire3933 = reg3911;
  assign wire3934 = (^($unsigned($signed(wire3906)) ?
                        (reg3914 ?
                            reg3922[(2'h3):(2'h2)] : (8'hb2)) : (reg3927[(3'h7):(3'h5)] ?
                            $unsigned(reg3928) : (reg3921 <<< reg3931))));
  assign wire3935 = (+(reg3914 | {((8'hb6) ? wire3904 : (8'hb1))}));
  module3936 #() modinst4540 (wire4539, clk, reg3926, reg3910, wire3902, reg3921, reg3929);
  assign wire4541 = ($signed($signed($signed(reg3914))) | (reg3929[(1'h0):(1'h0)] | $unsigned($unsigned(reg3913))));
  assign wire4542 = $signed(((|(wire4539 ?
                        wire3905 : reg3920)) ~^ $unsigned((8'ha5))));
  assign wire4543 = reg3922[(3'h5):(1'h0)];
  assign wire4544 = wire4542;
  assign wire4545 = (wire3903[(3'h5):(3'h5)] - $signed($unsigned(wire3905)));
  always
    @(posedge clk) begin
      if ((^~$signed($signed((wire3934 ? (8'had) : reg3923)))))
        begin
          reg4546 <= $unsigned((+$unsigned((~^reg3914))));
          for (forvar4547 = (1'h0); (forvar4547 < (2'h3)); forvar4547 = (forvar4547 + (1'h1)))
            begin
              if ($unsigned((reg3914 & (~|$signed(wire4541)))))
                begin
                  for (forvar4548 = (1'h0); (forvar4548 < (2'h2)); forvar4548 = (forvar4548 + (1'h1)))
                    begin
                      reg4549 <= $signed($signed(($unsigned(wire4542) ?
                          (~&wire4539) : wire4543)));
                      reg4550 <= $signed(($signed($signed(wire4545)) ?
                          ($signed(reg3916) ?
                              $unsigned(reg3926) : $unsigned(wire4543)) : reg3921[(4'hb):(3'h7)]));
                      reg4551 <= (reg3916 >= $signed(reg3914));
                    end
                  reg4552 <= (~^$unsigned((((8'hb9) == wire4544) ?
                      (wire4543 ?
                          reg3913 : wire4545) : reg3929[(3'h4):(2'h2)])));
                  if (reg3919)
                    begin
                      reg4553 <= wire3903;
                      reg4554 <= (!($signed(reg3931) >>> {reg4549}));
                    end
                  else
                    begin
                      reg4553 <= ($unsigned((8'hac)) ~^ (wire4543[(3'h6):(1'h1)] ^ $signed($unsigned(wire4543))));
                      reg4554 <= ($signed((|$signed(reg3930))) ?
                          (wire4541[(1'h1):(1'h0)] ?
                              $unsigned($unsigned((8'ha8))) : reg3910[(1'h0):(1'h0)]) : wire3908[(1'h0):(1'h0)]);
                      reg4555 <= ((~&(reg3916[(1'h0):(1'h0)] & {forvar4547})) ?
                          (wire3935[(3'h6):(3'h5)] ?
                              $signed($unsigned(reg3922)) : $signed((wire3906 * (8'hb6)))) : $unsigned(((reg3930 ?
                              reg3931 : reg3918) + {reg3921})));
                      reg4556 <= $signed((($unsigned(wire3908) ?
                          (wire4545 ?
                              reg3921 : (8'h9f)) : $signed(reg4553)) ^~ $unsigned((+reg3916))));
                    end
                  for (forvar4557 = (1'h0); (forvar4557 < (2'h3)); forvar4557 = (forvar4557 + (1'h1)))
                    begin
                      reg4558 <= reg3931[(1'h0):(1'h0)];
                      reg4559 <= ((reg3922[(1'h1):(1'h1)] <<< $unsigned($signed(wire3934))) ?
                          $signed(reg3929) : ((^reg3926) == ($signed((8'hb8)) ?
                              forvar4547[(4'h8):(3'h7)] : (8'hb4))));
                      reg4560 <= reg4549[(3'h6):(3'h5)];
                      reg4561 <= reg3914;
                    end
                end
              else
                begin
                  if ((&((wire3902[(1'h1):(1'h0)] ?
                      wire3934[(2'h3):(1'h0)] : (&(8'haa))) ~^ reg3910[(2'h2):(2'h2)])))
                    begin
                      reg4548 <= reg3911[(3'h7):(3'h6)];
                      reg4549 <= ($unsigned(reg3930[(2'h3):(1'h0)]) ?
                          ({reg4561[(3'h4):(1'h0)]} ?
                              wire3907 : $signed(reg3910[(2'h2):(2'h2)])) : reg3910);
                      reg4550 <= ($signed(($unsigned(wire3934) ?
                              $signed(reg4561) : wire3932[(1'h1):(1'h1)])) ?
                          $signed((&wire3932)) : reg3919);
                      reg4551 <= (+$unsigned($unsigned((wire4539 ?
                          reg4551 : reg4554))));
                    end
                  else
                    begin
                      reg4548 <= forvar4547[(3'h6):(2'h3)];
                      reg4549 <= ({wire3935[(1'h1):(1'h0)]} >= $unsigned($signed(reg4560)));
                    end
                  if ({reg3917[(3'h7):(3'h7)]})
                    begin
                      reg4552 <= reg4554[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg4552 <= {forvar4557[(2'h2):(1'h1)]};
                      reg4553 <= ($unsigned($unsigned({reg4548})) ?
                          ($signed($unsigned(reg3921)) * $unsigned($unsigned(reg4556))) : reg4556);
                      reg4554 <= (reg3920 | reg3917);
                    end
                end
            end
        end
      else
        begin
          if ((reg4551 ?
              (wire4544[(4'h9):(1'h0)] < $signed((reg4552 ?
                  reg3929 : reg3911))) : $unsigned(($unsigned(reg3916) && $unsigned(wire4545)))))
            begin
              for (forvar4546 = (1'h0); (forvar4546 < (2'h3)); forvar4546 = (forvar4546 + (1'h1)))
                begin
                  if ({((~(&reg3926)) ?
                          $signed((wire4545 ?
                              wire3933 : wire3906)) : (!$signed(wire3933)))})
                    begin
                      reg4547 <= {(8'h9f)};
                    end
                  else
                    begin
                      reg4547 <= (-(forvar4557[(2'h3):(2'h2)] ?
                          ((reg4555 && reg4560) ?
                              $signed((8'ha1)) : wire4541[(3'h5):(1'h1)]) : {(!reg4560)}));
                      reg4548 <= ((^~$signed(reg4548[(2'h2):(1'h1)])) <<< (forvar4547 == forvar4557));
                      reg4549 <= (~&((~&forvar4546) ?
                          {(reg4551 >>> (8'ha5))} : (reg3920[(2'h2):(2'h2)] ?
                              (&reg4560) : (wire3902 ? reg4560 : reg4550))));
                      reg4550 <= $signed($signed($unsigned((wire3906 ?
                          (8'ha0) : reg3928))));
                    end
                  if (reg3910[(1'h0):(1'h0)])
                    begin
                      reg4551 <= $signed($unsigned((~(reg3918 < reg4559))));
                      reg4552 <= $unsigned({$signed($unsigned(reg3917))});
                      reg4553 <= reg4550[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg4551 <= (!$unsigned(($signed(wire3933) >= (reg4547 ?
                          wire4543 : wire4541))));
                    end
                end
            end
          else
            begin
              for (forvar4546 = (1'h0); (forvar4546 < (1'h0)); forvar4546 = (forvar4546 + (1'h1)))
                begin
                  if ($signed(((~^wire3907[(1'h0):(1'h0)]) >>> ((reg4551 ?
                          reg3919 : (8'ha8)) ?
                      (^reg3911) : reg3929))))
                    begin
                      reg4547 <= reg4561;
                    end
                  else
                    begin
                      reg4547 <= reg4556[(3'h7):(3'h6)];
                    end
                  for (forvar4548 = (1'h0); (forvar4548 < (1'h1)); forvar4548 = (forvar4548 + (1'h1)))
                    begin
                      reg4549 <= $unsigned($signed(((wire3934 ?
                          reg3919 : (8'hb3)) > ((8'ha5) ?
                          reg4552 : wire4539))));
                    end
                  for (forvar4550 = (1'h0); (forvar4550 < (2'h2)); forvar4550 = (forvar4550 + (1'h1)))
                    begin
                      reg4551 <= reg3910;
                      reg4552 <= (~|reg4561[(2'h3):(1'h1)]);
                    end
                end
              for (forvar4553 = (1'h0); (forvar4553 < (1'h0)); forvar4553 = (forvar4553 + (1'h1)))
                begin
                  reg4554 <= $unsigned(reg4548[(3'h4):(2'h3)]);
                  if ((reg3917[(3'h5):(2'h3)] ?
                      (reg4551 ?
                          ((wire4542 <= reg4553) && $unsigned(reg3930)) : ((forvar4546 ^~ reg4555) ?
                              reg3930 : reg4561)) : $signed(((~|wire3903) - $signed(reg3927)))))
                    begin
                      reg4555 <= wire4543;
                      reg4556 <= (-forvar4557[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg4555 <= ((((reg3917 ?
                          reg3916 : reg4558) << {(8'haf)}) ^ reg4546[(4'hd):(3'h6)]) >= (forvar4550 << ((reg3911 ?
                          (8'haf) : reg4555) > (~|reg4553))));
                      reg4556 <= (^forvar4550[(2'h2):(2'h2)]);
                    end
                end
            end
        end
      for (forvar4562 = (1'h0); (forvar4562 < (2'h3)); forvar4562 = (forvar4562 + (1'h1)))
        begin
          reg4563 <= $unsigned({((wire3906 ?
                  forvar4557 : forvar4546) & forvar4546[(1'h1):(1'h0)])});
          if (reg3928)
            begin
              reg4564 <= $signed($signed(reg4550[(1'h1):(1'h1)]));
              for (forvar4565 = (1'h0); (forvar4565 < (1'h0)); forvar4565 = (forvar4565 + (1'h1)))
                begin
                  if ($signed((reg4552 ?
                      $signed($signed(wire3933)) : $unsigned((+reg4560)))))
                    begin
                      reg4566 <= reg4563;
                      reg4567 <= $signed($unsigned($unsigned({wire4544})));
                      reg4568 <= $signed($signed(((~^wire3903) ?
                          $signed(reg3926) : $unsigned(wire3902))));
                      reg4569 <= forvar4550[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg4566 <= reg4566[(2'h3):(1'h1)];
                      reg4567 <= reg4546;
                      reg4568 <= wire3932;
                    end
                end
              reg4570 <= reg4548;
              if ($unsigned($unsigned(reg3927)))
                begin
                  for (forvar4571 = (1'h0); (forvar4571 < (1'h0)); forvar4571 = (forvar4571 + (1'h1)))
                    begin
                      reg4572 <= (reg4553[(2'h2):(1'h0)] ?
                          {(-(~reg4559))} : wire3908);
                      reg4573 <= wire3935;
                    end
                  for (forvar4574 = (1'h0); (forvar4574 < (2'h3)); forvar4574 = (forvar4574 + (1'h1)))
                    begin
                      reg4575 <= (~$signed((^(reg4554 ? reg3919 : (8'hae)))));
                      reg4576 <= ((~^(forvar4546[(4'ha):(4'ha)] == $signed(reg4546))) ?
                          forvar4548[(2'h3):(2'h3)] : forvar4571);
                    end
                  reg4577 <= (+(~|($signed((8'ha6)) ?
                      (wire3902 != reg3920) : ((8'hb4) ?
                          forvar4557 : (8'ha9)))));
                  if ((wire3908 == (8'hb8)))
                    begin
                      reg4578 <= $unsigned(reg4553[(1'h0):(1'h0)]);
                      reg4579 <= (^reg4547[(3'h4):(1'h0)]);
                      reg4580 <= {reg4548};
                    end
                  else
                    begin
                      reg4578 <= $unsigned(({(forvar4548 ?
                                  reg4560 : wire4539)} ?
                          (&(~&reg4556)) : $signed((~^wire3902))));
                      reg4579 <= forvar4574;
                      reg4580 <= reg4556[(4'h9):(3'h6)];
                      reg4581 <= $unsigned(reg3931);
                    end
                end
              else
                begin
                  if ((^forvar4571))
                    begin
                      reg4571 <= $signed($unsigned($signed((reg4579 ?
                          reg4558 : (8'haa)))));
                      reg4572 <= $signed((reg4564 ?
                          (~&{wire3907}) : forvar4565[(1'h1):(1'h1)]));
                      reg4573 <= {($unsigned((reg4555 ? forvar4562 : (8'ha7))) ?
                              ({reg3920} ?
                                  (reg4546 ?
                                      wire3934 : (8'hb0)) : (reg3930 >> reg4567)) : (+reg3923))};
                    end
                  else
                    begin
                      reg4571 <= $signed($unsigned({forvar4550[(1'h0):(1'h0)]}));
                      reg4572 <= reg3916[(2'h3):(1'h0)];
                      reg4573 <= ((~^(&$unsigned((8'hb9)))) ^ $unsigned((~wire3934[(4'ha):(1'h0)])));
                    end
                  if ((~&(!(~|$signed(reg4549)))))
                    begin
                      reg4574 <= (~^reg4548[(3'h4):(3'h4)]);
                      reg4575 <= reg4570;
                      reg4576 <= (8'ha2);
                    end
                  else
                    begin
                      reg4574 <= reg3923;
                      reg4575 <= (reg4547[(3'h7):(1'h1)] > reg4578[(1'h0):(1'h0)]);
                    end
                  for (forvar4577 = (1'h0); (forvar4577 < (1'h1)); forvar4577 = (forvar4577 + (1'h1)))
                    begin
                      reg4578 <= reg4579[(3'h6):(2'h2)];
                    end
                end
            end
          else
            begin
              if ({wire4545[(4'hb):(3'h4)]})
                begin
                  for (forvar4564 = (1'h0); (forvar4564 < (1'h0)); forvar4564 = (forvar4564 + (1'h1)))
                    begin
                      reg4565 <= reg3920;
                      reg4566 <= $signed((^~$signed(reg3921)));
                      reg4567 <= $signed($unsigned((&forvar4577[(1'h1):(1'h1)])));
                    end
                  reg4568 <= $unsigned($signed((reg4546 + $unsigned(wire3908))));
                end
              else
                begin
                  for (forvar4564 = (1'h0); (forvar4564 < (1'h0)); forvar4564 = (forvar4564 + (1'h1)))
                    begin
                      reg4565 <= {(({reg4558} ?
                              (~^reg3923) : $unsigned(forvar4548)) & ((reg4566 ?
                                  reg3923 : (8'ha9)) ?
                              reg4581[(1'h1):(1'h1)] : (|wire4541)))};
                    end
                end
              for (forvar4569 = (1'h0); (forvar4569 < (2'h2)); forvar4569 = (forvar4569 + (1'h1)))
                begin
                  reg4570 <= (reg3914[(3'h6):(3'h6)] ?
                      ($unsigned((forvar4562 << reg4565)) ?
                          $unsigned((reg4556 ?
                              (8'hac) : reg3921)) : reg4564[(4'h9):(4'h9)]) : reg3914);
                end
              reg4571 <= (({(8'hba)} ? reg4568[(2'h3):(2'h2)] : wire3903) ?
                  $unsigned(((forvar4550 >> wire3933) ?
                      (forvar4547 ?
                          wire4545 : (8'hab)) : ((8'ha0) & reg4567))) : (reg4546[(4'hc):(4'ha)] ?
                      ((~&forvar4553) << (forvar4577 ^ forvar4557)) : wire4542[(4'h9):(2'h3)]));
            end
        end
      reg4582 <= $unsigned(reg4548);
    end
  assign wire4583 = $unsigned(reg3918[(4'hb):(4'h9)]);
  assign wire4584 = ((~^reg4549[(4'h9):(3'h6)]) ?
                        (reg3911[(3'h4):(1'h0)] > (!reg4556[(2'h2):(1'h1)])) : wire3903[(3'h4):(3'h4)]);
  always
    @(posedge clk) begin
      reg4585 <= (~((~&reg4546[(4'h8):(3'h7)]) ? reg4582 : reg4549));
      for (forvar4586 = (1'h0); (forvar4586 < (2'h3)); forvar4586 = (forvar4586 + (1'h1)))
        begin
          for (forvar4587 = (1'h0); (forvar4587 < (2'h2)); forvar4587 = (forvar4587 + (1'h1)))
            begin
              for (forvar4588 = (1'h0); (forvar4588 < (1'h0)); forvar4588 = (forvar4588 + (1'h1)))
                begin
                  for (forvar4589 = (1'h0); (forvar4589 < (2'h3)); forvar4589 = (forvar4589 + (1'h1)))
                    begin
                      reg4590 <= (|{(reg4559 ?
                              reg4565[(1'h0):(1'h0)] : (reg3917 * reg3927))});
                      reg4591 <= (reg4555 ?
                          {$unsigned((+reg3926))} : ($unsigned({reg4580}) & reg4578));
                    end
                  if (reg3931)
                    begin
                      reg4592 <= $signed({(~^(wire4543 ? wire3902 : (8'ha4)))});
                      reg4593 <= (&(({forvar4587} ?
                              (reg4592 ? reg3919 : reg4576) : (+reg3921)) ?
                          {(-(8'hb0))} : (~&wire4543[(2'h2):(2'h2)])));
                    end
                  else
                    begin
                      reg4592 <= (-$signed((((8'h9d) ?
                          wire4544 : reg3922) ^~ (reg4552 ?
                          reg4549 : reg4581))));
                      reg4593 <= {wire4583};
                      reg4594 <= $unsigned(reg4576);
                    end
                  for (forvar4595 = (1'h0); (forvar4595 < (1'h1)); forvar4595 = (forvar4595 + (1'h1)))
                    begin
                      reg4596 <= reg3910[(2'h2):(1'h0)];
                      reg4597 <= $unsigned({$signed((reg3921 ?
                              reg4594 : reg4579))});
                      reg4598 <= $signed(reg4593[(2'h3):(1'h0)]);
                      reg4599 <= {$unsigned(reg4551[(4'h9):(1'h0)])};
                    end
                  if (reg3923[(3'h7):(1'h1)])
                    begin
                      reg4600 <= $unsigned((^~reg4568));
                    end
                  else
                    begin
                      reg4600 <= (({$signed(forvar4588)} ?
                          {(reg4582 ?
                                  reg4548 : reg4591)} : {{reg4554}}) * wire3933);
                      reg4601 <= {$unsigned($unsigned({reg3919}))};
                      reg4602 <= reg3920;
                    end
                end
              for (forvar4603 = (1'h0); (forvar4603 < (2'h3)); forvar4603 = (forvar4603 + (1'h1)))
                begin
                  reg4604 <= reg4555;
                end
              for (forvar4605 = (1'h0); (forvar4605 < (2'h2)); forvar4605 = (forvar4605 + (1'h1)))
                begin
                  for (forvar4606 = (1'h0); (forvar4606 < (1'h0)); forvar4606 = (forvar4606 + (1'h1)))
                    begin
                      reg4607 <= (reg3918 >>> $signed($signed((reg4549 ^~ reg4594))));
                      reg4608 <= reg4598;
                      reg4609 <= (($unsigned($signed(reg4553)) ?
                              $signed((^~reg4565)) : $unsigned($signed(reg4569))) ?
                          {$signed($unsigned(reg4582))} : {($signed(reg4563) <= reg4549[(4'h9):(1'h0)])});
                      reg4610 <= (reg3919 ^ $unsigned($signed(((8'hb8) > reg4546))));
                    end
                  if (($unsigned(({wire3902} < ((8'hb2) ?
                      (8'hba) : forvar4605))) + (reg3916 >>> (&reg3926))))
                    begin
                      reg4611 <= (({wire4583} ?
                              $unsigned($unsigned((8'h9d))) : ((~forvar4588) * {wire3904})) ?
                          (($signed((8'h9c)) ?
                              (wire3934 >>> reg3911) : (wire4543 <= wire3903)) & (reg4546[(2'h2):(1'h1)] >> (reg3930 ?
                              reg4561 : reg4572))) : reg4573[(2'h3):(2'h3)]);
                      reg4612 <= (^~reg4548);
                      reg4613 <= (reg4576 ?
                          {((-reg4560) ?
                                  $unsigned(reg3910) : (~reg4556))} : $unsigned((^(^~reg4601))));
                      reg4614 <= (reg4573 ?
                          (!($unsigned(wire4539) * (~reg4582))) : {(reg3931[(3'h4):(3'h4)] >> reg4570[(4'ha):(1'h0)])});
                    end
                  else
                    begin
                      reg4611 <= (reg4556 ?
                          $unsigned($signed((reg4579 ?
                              reg3922 : reg3913))) : ({(reg3913 ~^ wire4542)} ?
                              ($unsigned((8'ha3)) | (wire3904 ?
                                  wire4539 : reg4549)) : $unsigned((|reg3927))));
                      reg4612 <= (reg4549 + $unsigned((wire3902[(3'h4):(1'h1)] ?
                          reg4555[(2'h3):(2'h3)] : reg4613)));
                    end
                  if (((~&($unsigned(reg4601) ?
                          $signed((8'ha3)) : (~reg4558))) ?
                      ((&$signed(reg4608)) != (~&(reg4612 - wire3907))) : wire4583[(2'h2):(2'h2)]))
                    begin
                      reg4615 <= (wire3908[(5'h10):(4'hb)] ?
                          reg4609[(4'hd):(4'hb)] : reg4611[(3'h6):(2'h2)]);
                      reg4616 <= ($signed((~|$unsigned(reg3928))) <<< $signed((8'h9e)));
                      reg4617 <= ({reg4570} ?
                          $signed(((~|(8'ha0)) ^~ reg3918[(2'h2):(1'h0)])) : (8'ha6));
                    end
                  else
                    begin
                      reg4615 <= $signed(reg4558);
                      reg4616 <= reg4571;
                      reg4617 <= {reg4565[(1'h1):(1'h0)]};
                      reg4618 <= $unsigned({{reg4580}});
                    end
                end
              if ($unsigned(reg4615[(2'h2):(1'h1)]))
                begin
                  for (forvar4619 = (1'h0); (forvar4619 < (2'h3)); forvar4619 = (forvar4619 + (1'h1)))
                    begin
                      reg4620 <= ($signed({{reg4599}}) ~^ {$unsigned({reg4600})});
                      reg4621 <= (($signed((8'hac)) ?
                              reg3927[(1'h0):(1'h0)] : ((wire3932 ?
                                  reg3911 : reg4592) & $unsigned((8'ha1)))) ?
                          (~$unsigned((forvar4588 ?
                              reg3910 : wire4583))) : $signed(($unsigned(reg4608) && $unsigned(reg4546))));
                    end
                  for (forvar4622 = (1'h0); (forvar4622 < (2'h2)); forvar4622 = (forvar4622 + (1'h1)))
                    begin
                      reg4623 <= (+$unsigned((reg3916[(2'h3):(1'h0)] ?
                          $unsigned(reg4607) : (8'ha0))));
                      reg4624 <= (((reg4581 ? reg4610 : {reg4615}) ?
                          reg4554[(2'h2):(2'h2)] : ($unsigned((8'ha6)) ?
                              $signed(reg4572) : reg4546)) == wire4543[(4'h8):(1'h0)]);
                      reg4625 <= ({((&wire3902) ~^ {reg3923})} <<< reg4575[(2'h3):(2'h3)]);
                      reg4626 <= (((wire3932[(1'h1):(1'h1)] ?
                                  (reg4613 ~^ forvar4606) : (+reg4555)) ?
                              $signed((reg4598 ^~ (8'hb4))) : {reg4597}) ?
                          (^~$unsigned(reg4580)) : $signed(reg3923[(1'h1):(1'h1)]));
                    end
                  for (forvar4627 = (1'h0); (forvar4627 < (1'h1)); forvar4627 = (forvar4627 + (1'h1)))
                    begin
                      reg4628 <= $signed(forvar4587);
                      reg4629 <= ({reg4565[(2'h3):(1'h1)]} ?
                          ($signed(wire3907[(1'h1):(1'h0)]) ?
                              (reg4565[(1'h0):(1'h0)] <= (reg4624 ?
                                  wire3905 : reg3926)) : $unsigned({(8'hb7)})) : reg4614);
                      reg4630 <= $unsigned($signed((~^wire3932)));
                    end
                  reg4631 <= $unsigned($unsigned(((&reg4555) ?
                      (reg3916 ? reg4594 : wire4545) : {(8'ha9)})));
                end
              else
                begin
                  reg4619 <= reg4567[(3'h7):(3'h5)];
                  if ($unsigned(forvar4595[(3'h4):(3'h4)]))
                    begin
                      reg4620 <= $unsigned($unsigned($unsigned($unsigned(reg4554))));
                    end
                  else
                    begin
                      reg4620 <= $signed(reg4559[(3'h5):(1'h1)]);
                    end
                  for (forvar4621 = (1'h0); (forvar4621 < (1'h1)); forvar4621 = (forvar4621 + (1'h1)))
                    begin
                      reg4622 <= (8'hba);
                      reg4623 <= $unsigned({reg4552[(4'hc):(1'h1)]});
                      reg4624 <= reg3918;
                      reg4625 <= (8'had);
                    end
                end
            end
        end
      for (forvar4632 = (1'h0); (forvar4632 < (2'h2)); forvar4632 = (forvar4632 + (1'h1)))
        begin
          for (forvar4633 = (1'h0); (forvar4633 < (2'h2)); forvar4633 = (forvar4633 + (1'h1)))
            begin
              if ($signed($unsigned($unsigned(reg4619[(1'h0):(1'h0)]))))
                begin
                  if ($signed(($signed((~&reg4563)) ?
                      (|(reg3917 ?
                          (8'hb5) : (8'haf))) : (^reg4554[(2'h2):(1'h1)]))))
                    begin
                      reg4634 <= {($signed($unsigned(reg3930)) ?
                              {(forvar4603 + (8'h9c))} : reg4614[(3'h7):(1'h0)])};
                    end
                  else
                    begin
                      reg4634 <= $signed((&((^~wire3934) ^~ (forvar4606 ^ reg3930))));
                    end
                  reg4635 <= {reg4611[(4'h9):(3'h5)]};
                  reg4636 <= $signed((-reg4580));
                end
              else
                begin
                  for (forvar4634 = (1'h0); (forvar4634 < (1'h1)); forvar4634 = (forvar4634 + (1'h1)))
                    begin
                      reg4635 <= (&$signed($unsigned(reg4575)));
                      reg4636 <= {(~|reg4614)};
                      reg4637 <= reg3922[(1'h1):(1'h0)];
                      reg4638 <= $signed($signed($signed($signed(reg4618))));
                    end
                  if (reg4594[(4'h8):(1'h1)])
                    begin
                      reg4639 <= (&reg3919[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg4639 <= $signed({$unsigned($unsigned(forvar4634))});
                      reg4640 <= reg4585[(2'h3):(2'h3)];
                    end
                end
              reg4641 <= reg4585;
              for (forvar4642 = (1'h0); (forvar4642 < (2'h2)); forvar4642 = (forvar4642 + (1'h1)))
                begin
                  if ($unsigned((reg4630 ?
                      ($signed(reg3923) ?
                          (reg4558 * reg4585) : $signed((8'h9c))) : ($unsigned(wire4545) ?
                          {forvar4588} : (~&reg4594)))))
                    begin
                      reg4643 <= reg4548;
                      reg4644 <= $unsigned(($signed(reg4608) ?
                          ($unsigned(reg4635) ^~ (reg4579 > (8'haf))) : ({(8'h9f)} ?
                              reg3927[(1'h0):(1'h0)] : $signed(forvar4634))));
                    end
                  else
                    begin
                      reg4643 <= (~^(8'hb0));
                    end
                  reg4645 <= wire3908[(4'h8):(1'h0)];
                end
            end
          reg4646 <= ($signed({(wire3908 ?
                  wire3904 : (8'hac))}) <<< reg4623[(4'ha):(1'h0)]);
          for (forvar4647 = (1'h0); (forvar4647 < (1'h0)); forvar4647 = (forvar4647 + (1'h1)))
            begin
              reg4648 <= ({(reg3910 ?
                          (wire3907 >> forvar4589) : (reg4625 ?
                              (8'hb4) : reg4572))} ?
                  reg4553[(1'h1):(1'h1)] : {({reg4582} >> $signed(reg3930))});
            end
        end
    end
  always
    @(posedge clk) begin
      if ((!reg3919[(4'hc):(3'h6)]))
        begin
          if ($signed(wire4541))
            begin
              if ({(($unsigned(reg4635) <= reg3928[(2'h2):(2'h2)]) ?
                      (8'hb8) : ({reg4619} ?
                          (wire3905 ?
                              wire3933 : reg4600) : $signed(wire3904)))})
                begin
                  for (forvar4649 = (1'h0); (forvar4649 < (2'h3)); forvar4649 = (forvar4649 + (1'h1)))
                    begin
                      reg4650 <= ({reg4598[(3'h5):(2'h2)]} ~^ reg4604[(3'h5):(2'h3)]);
                    end
                  for (forvar4651 = (1'h0); (forvar4651 < (2'h3)); forvar4651 = (forvar4651 + (1'h1)))
                    begin
                      reg4652 <= reg4598[(1'h0):(1'h0)];
                      reg4653 <= reg4643;
                      reg4654 <= $signed((^~$unsigned({wire3904})));
                      reg4655 <= $signed($signed((!wire3932[(1'h0):(1'h0)])));
                    end
                  reg4656 <= reg3929[(2'h2):(1'h1)];
                  reg4657 <= (reg4609 ?
                      (reg4604 ?
                          $signed((reg4630 * (8'ha5))) : $signed($signed(reg4628))) : $signed(reg4549[(3'h6):(3'h4)]));
                end
              else
                begin
                  reg4649 <= reg3916;
                  for (forvar4650 = (1'h0); (forvar4650 < (2'h3)); forvar4650 = (forvar4650 + (1'h1)))
                    begin
                      reg4651 <= reg4617[(2'h2):(2'h2)];
                      reg4652 <= $signed($unsigned(((reg3927 > reg4571) >>> $unsigned(reg4639))));
                    end
                end
              if (({(reg4612[(3'h4):(2'h3)] ?
                      reg4574[(1'h0):(1'h0)] : $signed(reg4571))} + ($signed($unsigned(wire3933)) ?
                  $signed((wire3935 ?
                      reg4635 : (8'haa))) : ($signed(reg4649) + (-(8'hab))))))
                begin
                  if (((reg3920[(1'h1):(1'h1)] ?
                      $unsigned(reg4552[(2'h2):(2'h2)]) : reg4618) == $unsigned(reg4546)))
                    begin
                      reg4658 <= $unsigned($signed((-(wire3905 & reg3929))));
                      reg4659 <= $signed($unsigned(($unsigned(reg4611) == (wire3904 >>> reg3930))));
                      reg4660 <= reg4555;
                      reg4661 <= $unsigned((~&reg4568));
                    end
                  else
                    begin
                      reg4658 <= ({reg4575[(3'h5):(1'h1)]} ^ $signed($signed($unsigned(reg4594))));
                      reg4659 <= reg4599;
                      reg4660 <= $unsigned(reg4578);
                    end
                end
              else
                begin
                  if ($signed($unsigned(($signed(reg3918) ?
                      $signed(wire3906) : reg4594))))
                    begin
                      reg4658 <= $signed($signed((8'ha5)));
                      reg4659 <= reg4625[(4'ha):(3'h4)];
                      reg4660 <= reg4558;
                      reg4661 <= $signed(((((8'h9e) >> reg4645) << (&wire3904)) ?
                          reg4554[(4'h8):(1'h0)] : $signed($unsigned((8'hba)))));
                    end
                  else
                    begin
                      reg4658 <= $signed(reg3920);
                      reg4659 <= reg4652[(1'h1):(1'h1)];
                      reg4660 <= reg4580;
                    end
                  if (reg4579)
                    begin
                      reg4662 <= {{$unsigned($unsigned(wire3902))}};
                      reg4663 <= (8'haf);
                      reg4664 <= ({(reg4612[(3'h4):(2'h2)] > reg4661[(3'h4):(3'h4)])} + (forvar4649 ?
                          $unsigned({wire3902}) : (^(reg4572 ?
                              reg3921 : reg4574))));
                    end
                  else
                    begin
                      reg4662 <= {reg3931[(3'h4):(2'h2)]};
                    end
                  for (forvar4665 = (1'h0); (forvar4665 < (2'h2)); forvar4665 = (forvar4665 + (1'h1)))
                    begin
                      reg4666 <= (8'hb7);
                      reg4667 <= {(($signed(reg4549) << {(8'had)}) ?
                              reg3913[(3'h4):(3'h4)] : $signed($signed(wire3933)))};
                      reg4668 <= (reg4558[(3'h6):(3'h5)] ?
                          $signed(reg4639[(4'ha):(3'h5)]) : reg4596);
                    end
                end
              if ((8'ha4))
                begin
                  if ($signed($signed(((~reg4548) ? (8'ha2) : (~|reg4650)))))
                    begin
                      reg4669 <= wire3932[(1'h1):(1'h0)];
                      reg4670 <= (~^reg4556[(4'h9):(2'h3)]);
                    end
                  else
                    begin
                      reg4669 <= (reg4634[(4'h9):(3'h6)] * $unsigned({reg4570[(1'h1):(1'h1)]}));
                    end
                  reg4671 <= $unsigned((((reg4560 ~^ reg4597) ?
                          $signed(reg3923) : $unsigned(reg3916)) ?
                      wire3933 : (reg4553[(2'h3):(1'h0)] >= $signed(reg4613))));
                end
              else
                begin
                  for (forvar4669 = (1'h0); (forvar4669 < (1'h0)); forvar4669 = (forvar4669 + (1'h1)))
                    begin
                      reg4670 <= wire4541[(3'h4):(2'h3)];
                    end
                  if ($signed(reg3929[(3'h4):(2'h2)]))
                    begin
                      reg4671 <= (!(8'h9c));
                    end
                  else
                    begin
                      reg4671 <= ((~^$unsigned(reg4552)) ~^ (^reg4662[(3'h6):(3'h4)]));
                      reg4672 <= (^(((reg4581 ? (8'hb4) : reg4613) ?
                          (reg4612 ? reg4669 : reg4658) : (reg3926 ?
                              reg4635 : reg4612)) > ($signed(wire4541) ?
                          (reg3923 ? reg3926 : reg4617) : (wire3907 ?
                              reg4581 : (8'ha9)))));
                      reg4673 <= {((^~reg4580[(3'h5):(3'h4)]) && $unsigned(((8'ha9) ?
                              (8'ha7) : reg4598)))};
                    end
                  if ((reg4666[(3'h7):(3'h4)] ?
                      (-($unsigned(reg4669) ^ (wire4539 != wire3906))) : $signed($signed($unsigned(reg4613)))))
                    begin
                      reg4674 <= ($unsigned(($signed((8'ha4)) ?
                          {reg4658} : $signed(reg4568))) * reg3926);
                      reg4675 <= ($unsigned((~&$unsigned(reg4653))) ^ (!reg4592[(3'h5):(3'h5)]));
                      reg4676 <= ($signed((8'h9e)) ~^ $signed({$unsigned(reg4607)}));
                    end
                  else
                    begin
                      reg4674 <= $signed(reg4611);
                      reg4675 <= ($signed((|reg4608)) & (~((reg3917 ?
                          reg4619 : reg4671) ~^ reg4666)));
                      reg4676 <= {(((reg3910 >> reg4617) ?
                              $signed(wire4543) : $signed(forvar4650)) & {(reg4660 << reg4582)})};
                      reg4677 <= reg4546[(2'h2):(1'h0)];
                    end
                  for (forvar4678 = (1'h0); (forvar4678 < (1'h0)); forvar4678 = (forvar4678 + (1'h1)))
                    begin
                      reg4679 <= ((reg4568[(3'h5):(1'h1)] ?
                          $signed(reg4623) : (^(reg4590 ?
                              reg4624 : reg4653))) << ($unsigned({reg4592}) + (+reg4671)));
                      reg4680 <= {(^reg4566)};
                      reg4681 <= $unsigned((~|{{reg3921}}));
                      reg4682 <= ({$signed((8'hb6))} ?
                          (8'hb7) : {(((8'hb5) ^~ (8'hb6)) | (reg4618 ?
                                  wire3908 : reg4662))});
                    end
                end
              for (forvar4683 = (1'h0); (forvar4683 < (1'h0)); forvar4683 = (forvar4683 + (1'h1)))
                begin
                  for (forvar4684 = (1'h0); (forvar4684 < (1'h0)); forvar4684 = (forvar4684 + (1'h1)))
                    begin
                      reg4685 <= (^(reg4579 ?
                          $unsigned($unsigned(reg3917)) : reg4548));
                      reg4686 <= forvar4683[(1'h0):(1'h0)];
                    end
                  for (forvar4687 = (1'h0); (forvar4687 < (1'h1)); forvar4687 = (forvar4687 + (1'h1)))
                    begin
                      reg4688 <= $unsigned((~reg4613[(4'he):(3'h5)]));
                      reg4689 <= (wire3905[(4'h8):(1'h0)] | (((reg4676 ^~ reg4601) ?
                              (reg4608 | reg4667) : $unsigned(reg4686)) ?
                          ((reg4662 ?
                              reg4621 : reg4639) < (~&reg4576)) : (~^(~reg4579))));
                      reg4690 <= (-(!(reg4650[(1'h1):(1'h1)] || {reg4566})));
                    end
                  reg4691 <= wire3902[(1'h0):(1'h0)];
                end
            end
          else
            begin
              if (reg4666[(3'h6):(3'h4)])
                begin
                  reg4649 <= $signed(forvar4665);
                end
              else
                begin
                  for (forvar4649 = (1'h0); (forvar4649 < (1'h0)); forvar4649 = (forvar4649 + (1'h1)))
                    begin
                      reg4650 <= (reg4569[(1'h0):(1'h0)] ?
                          (wire4542 + {(~(8'hab))}) : reg3918);
                      reg4651 <= {$signed((reg4628[(1'h1):(1'h1)] ~^ (reg4634 ?
                              reg4661 : reg4570)))};
                    end
                end
              for (forvar4652 = (1'h0); (forvar4652 < (1'h1)); forvar4652 = (forvar4652 + (1'h1)))
                begin
                  if (reg4672)
                    begin
                      reg4653 <= $signed(($unsigned($unsigned(wire4542)) ?
                          $unsigned($unsigned((8'ha9))) : $unsigned($signed(forvar4684))));
                      reg4654 <= $unsigned((8'ha3));
                      reg4655 <= (((wire3908 - reg4622[(4'h8):(2'h3)]) ?
                              $unsigned(reg4629) : ((8'hae) ^~ (reg4655 != reg4550))) ?
                          (($unsigned(reg4594) ?
                              (&reg4681) : {reg4661}) > (8'h9f)) : $signed(reg4658));
                    end
                  else
                    begin
                      reg4653 <= (^~(reg4635[(2'h3):(2'h3)] == ($unsigned(reg4577) >= (~&(8'haf)))));
                      reg4654 <= {reg4675[(1'h0):(1'h0)]};
                    end
                  for (forvar4656 = (1'h0); (forvar4656 < (1'h1)); forvar4656 = (forvar4656 + (1'h1)))
                    begin
                      reg4657 <= wire3903;
                      reg4658 <= ($signed((&{wire3932})) || reg4649[(3'h6):(2'h2)]);
                    end
                  if (reg4575)
                    begin
                      reg4659 <= ($signed((^~reg4625[(3'h5):(1'h0)])) < (&reg3918[(1'h0):(1'h0)]));
                      reg4660 <= ($unsigned((reg3919 ?
                              $unsigned(reg4548) : $unsigned(reg4622))) ?
                          {reg3921[(4'hb):(3'h4)]} : (+reg4670));
                      reg4661 <= {(8'ha9)};
                      reg4662 <= $signed($unsigned({(&reg4672)}));
                    end
                  else
                    begin
                      reg4659 <= ($unsigned((!reg4644)) ?
                          ({(^reg3910)} ?
                              (~reg4621[(3'h4):(1'h0)]) : ($signed(reg4600) << $signed(reg4646))) : $signed(reg4612[(3'h4):(1'h1)]));
                      reg4660 <= $unsigned(($unsigned(reg4614) + reg4559));
                      reg4661 <= reg4599[(2'h2):(2'h2)];
                      reg4662 <= (forvar4651 ?
                          reg4641 : (reg4674 & reg3914[(1'h1):(1'h0)]));
                    end
                  if ($signed((reg4590[(1'h1):(1'h0)] - (~^(reg4572 >> (8'hb1))))))
                    begin
                      reg4663 <= (-(!(~&{reg4636})));
                      reg4664 <= ($signed((!$unsigned(reg4664))) || (($signed(reg4680) >= (reg4573 > wire4584)) <= forvar4656[(2'h3):(2'h3)]));
                    end
                  else
                    begin
                      reg4663 <= $unsigned(reg4571[(3'h4):(2'h3)]);
                      reg4664 <= $unsigned((8'h9d));
                      reg4665 <= (&{$unsigned(reg4618[(3'h5):(2'h3)])});
                    end
                end
              for (forvar4666 = (1'h0); (forvar4666 < (2'h2)); forvar4666 = (forvar4666 + (1'h1)))
                begin
                  for (forvar4667 = (1'h0); (forvar4667 < (2'h2)); forvar4667 = (forvar4667 + (1'h1)))
                    begin
                      reg4668 <= $signed((((&reg4649) ? reg4601 : reg4577) ?
                          reg4665[(3'h5):(1'h1)] : ({wire4541} ?
                              (reg4685 ? reg4636 : reg4644) : (+reg4600))));
                    end
                  for (forvar4669 = (1'h0); (forvar4669 < (1'h1)); forvar4669 = (forvar4669 + (1'h1)))
                    begin
                      reg4670 <= (+reg4600);
                      reg4671 <= (reg4553[(1'h1):(1'h0)] * (~|(|(wire3932 ~^ reg4549))));
                      reg4672 <= $unsigned({(reg4559[(3'h6):(3'h6)] >= $unsigned(reg4596))});
                    end
                  reg4673 <= $signed((reg4660 ?
                      reg4547[(5'h10):(1'h0)] : reg4663));
                end
            end
          reg4692 <= (reg4660[(3'h7):(2'h2)] ?
              ($unsigned(reg4655[(4'ha):(3'h6)]) + ((reg4591 ?
                  (8'ha3) : reg4653) & forvar4652)) : (reg4549[(4'ha):(4'h8)] >= reg4673));
          for (forvar4693 = (1'h0); (forvar4693 < (1'h0)); forvar4693 = (forvar4693 + (1'h1)))
            begin
              for (forvar4694 = (1'h0); (forvar4694 < (2'h3)); forvar4694 = (forvar4694 + (1'h1)))
                begin
                  for (forvar4695 = (1'h0); (forvar4695 < (1'h0)); forvar4695 = (forvar4695 + (1'h1)))
                    begin
                      reg4696 <= $signed(($unsigned(forvar4649) ?
                          reg4611[(4'hc):(4'h8)] : (reg3922[(4'h9):(3'h6)] + (-reg4578))));
                      reg4697 <= forvar4656[(4'h9):(3'h7)];
                      reg4698 <= (forvar4652[(2'h3):(2'h3)] ?
                          ($signed($unsigned(reg4679)) ?
                              reg4610 : reg4672[(3'h7):(3'h7)]) : {((reg4666 ?
                                  reg3918 : reg4676) <= {(8'hb1)})});
                      reg4699 <= $unsigned($signed({(reg3926 ?
                              reg4622 : reg3914)}));
                    end
                  if (reg4639)
                    begin
                      reg4700 <= $signed($unsigned((forvar4666 ?
                          (~^reg4566) : (^~reg4567))));
                    end
                  else
                    begin
                      reg4700 <= reg4699;
                    end
                end
            end
          reg4701 <= $unsigned({reg4670[(1'h1):(1'h0)]});
        end
      else
        begin
          for (forvar4649 = (1'h0); (forvar4649 < (1'h0)); forvar4649 = (forvar4649 + (1'h1)))
            begin
              reg4650 <= (^wire4542);
              if (reg4697[(3'h4):(2'h3)])
                begin
                  for (forvar4651 = (1'h0); (forvar4651 < (2'h2)); forvar4651 = (forvar4651 + (1'h1)))
                    begin
                      reg4652 <= (!reg3913);
                      reg4653 <= $signed(reg4692);
                      reg4654 <= ($signed($unsigned({reg4582})) ?
                          reg4613 : reg4658[(1'h1):(1'h1)]);
                      reg4655 <= ($unsigned((!(!reg4566))) ?
                          (~^{forvar4669}) : reg4631[(2'h2):(1'h0)]);
                    end
                end
              else
                begin
                  if ($signed(reg4581[(2'h2):(2'h2)]))
                    begin
                      reg4651 <= (forvar4665[(1'h0):(1'h0)] ?
                          reg4655[(4'hb):(4'ha)] : ($unsigned(reg4582) ?
                              $signed(reg4682) : (reg4671[(2'h3):(1'h1)] <= reg4673)));
                      reg4652 <= $unsigned({$signed($unsigned(reg4575))});
                    end
                  else
                    begin
                      reg4651 <= {$signed(forvar4695[(4'h8):(1'h1)])};
                    end
                  reg4653 <= reg4688[(3'h6):(3'h6)];
                end
              for (forvar4656 = (1'h0); (forvar4656 < (1'h0)); forvar4656 = (forvar4656 + (1'h1)))
                begin
                  if ($signed({$signed((wire3932 + reg4690))}))
                    begin
                      reg4657 <= (~|$signed(((reg3928 ? reg4685 : reg4624) ?
                          (^~reg4547) : {reg4636})));
                    end
                  else
                    begin
                      reg4657 <= (($signed($unsigned((8'h9d))) & ({(8'ha0)} ?
                              (~|forvar4666) : reg3911)) ?
                          ($signed((|reg4629)) != (|(!(8'hba)))) : ((forvar4669[(2'h2):(1'h0)] ^ reg4629) ?
                              $signed($unsigned((8'h9d))) : reg3930[(1'h0):(1'h0)]));
                      reg4658 <= $unsigned(($signed(reg4651) ?
                          (wire3933 ?
                              (-reg4648) : (reg4607 >> reg4624)) : (^~$unsigned(reg3923))));
                      reg4659 <= $signed((($unsigned(reg4591) && (forvar4652 ?
                              reg4649 : reg4641)) ?
                          $signed($signed((8'ha2))) : ((reg4552 ?
                                  reg4690 : reg4608) ?
                              wire4541[(2'h3):(1'h0)] : reg4585)));
                    end
                  reg4660 <= ($unsigned({reg4551[(2'h2):(1'h0)]}) | (8'ha2));
                  reg4661 <= $unsigned({reg4692[(1'h0):(1'h0)]});
                end
              for (forvar4662 = (1'h0); (forvar4662 < (2'h3)); forvar4662 = (forvar4662 + (1'h1)))
                begin
                  if ($signed($unsigned(reg4674)))
                    begin
                      reg4663 <= $signed($signed($unsigned($signed(reg4641))));
                      reg4664 <= reg3930;
                      reg4665 <= reg4669;
                    end
                  else
                    begin
                      reg4663 <= reg4689[(3'h6):(3'h5)];
                      reg4664 <= $signed($signed((|{wire4584})));
                      reg4665 <= (reg4613 ? reg4560 : reg3923);
                    end
                  if (($unsigned((((8'hac) ? reg4677 : reg4576) ?
                      (reg4656 & forvar4665) : $signed((8'haa)))) >> {{reg4548[(3'h6):(2'h3)]}}))
                    begin
                      reg4666 <= $signed($unsigned({(reg4574 ?
                              wire4583 : reg4558)}));
                      reg4667 <= $unsigned(reg4622[(1'h1):(1'h0)]);
                      reg4668 <= reg4561;
                    end
                  else
                    begin
                      reg4666 <= reg4690[(1'h1):(1'h1)];
                      reg4667 <= (~|$signed(wire3907));
                      reg4668 <= (wire4583 < $unsigned($signed((^(8'hb4)))));
                    end
                  reg4669 <= ($signed($signed((~^reg4564))) ?
                      ((~&(~^reg3930)) != ({reg4680} ?
                          reg4573 : reg3928[(1'h1):(1'h0)])) : reg4624[(2'h2):(2'h2)]);
                end
            end
          for (forvar4670 = (1'h0); (forvar4670 < (1'h1)); forvar4670 = (forvar4670 + (1'h1)))
            begin
              for (forvar4671 = (1'h0); (forvar4671 < (1'h1)); forvar4671 = (forvar4671 + (1'h1)))
                begin
                  for (forvar4672 = (1'h0); (forvar4672 < (2'h3)); forvar4672 = (forvar4672 + (1'h1)))
                    begin
                      reg4673 <= $signed((~&reg4567[(3'h7):(1'h1)]));
                      reg4674 <= wire4542[(1'h1):(1'h0)];
                      reg4675 <= $signed($unsigned({$signed(reg3920)}));
                    end
                  reg4676 <= (reg4688 ?
                      (-$unsigned($unsigned(reg4578))) : $unsigned((-(!reg4560))));
                  for (forvar4677 = (1'h0); (forvar4677 < (2'h3)); forvar4677 = (forvar4677 + (1'h1)))
                    begin
                      reg4678 <= (-reg4608);
                      reg4679 <= (8'hb1);
                    end
                  reg4680 <= reg3927[(2'h2):(2'h2)];
                end
              reg4681 <= (reg4568[(3'h4):(3'h4)] ?
                  ((~|$unsigned(reg4640)) ?
                      wire4539 : $signed((reg4690 ?
                          reg4644 : reg4645))) : ((^~$signed(reg4679)) ?
                      reg4621[(1'h1):(1'h0)] : $unsigned(reg4602)));
              if (reg4688)
                begin
                  reg4682 <= $unsigned(forvar4651[(2'h3):(2'h2)]);
                end
              else
                begin
                  for (forvar4682 = (1'h0); (forvar4682 < (1'h1)); forvar4682 = (forvar4682 + (1'h1)))
                    begin
                      reg4683 <= reg4622[(4'hb):(3'h5)];
                      reg4684 <= (~(~&{$unsigned(reg4553)}));
                    end
                  for (forvar4685 = (1'h0); (forvar4685 < (2'h3)); forvar4685 = (forvar4685 + (1'h1)))
                    begin
                      reg4686 <= (({reg4546} < reg4625) > $signed(reg4552));
                      reg4687 <= $unsigned($unsigned((~{reg4688})));
                      reg4688 <= reg4646;
                      reg4689 <= $unsigned(reg4601[(2'h3):(2'h3)]);
                    end
                  for (forvar4690 = (1'h0); (forvar4690 < (1'h0)); forvar4690 = (forvar4690 + (1'h1)))
                    begin
                      reg4691 <= $unsigned(($unsigned($unsigned((8'ha3))) ?
                          $unsigned($signed(reg4665)) : reg4645[(4'ha):(2'h3)]));
                      reg4692 <= reg4564[(1'h1):(1'h1)];
                    end
                end
            end
          for (forvar4693 = (1'h0); (forvar4693 < (1'h1)); forvar4693 = (forvar4693 + (1'h1)))
            begin
              if ($signed(((^~(reg4575 >>> reg4554)) == ($unsigned(reg4698) ?
                  (wire3905 == (8'hae)) : (^~(8'h9c))))))
                begin
                  for (forvar4694 = (1'h0); (forvar4694 < (1'h1)); forvar4694 = (forvar4694 + (1'h1)))
                    begin
                      reg4695 <= (~&$signed($unsigned((~&reg3920))));
                      reg4696 <= $signed($unsigned((8'ha5)));
                      reg4697 <= ((-wire3904[(2'h2):(2'h2)]) ?
                          ($signed(reg4622[(4'he):(4'hc)]) ?
                              reg4582 : (reg4654[(4'hd):(3'h4)] ?
                                  $unsigned(reg3923) : (reg3919 ?
                                      reg4611 : reg4619))) : $unsigned((~&$signed(reg4697))));
                      reg4698 <= (~^((8'hac) ?
                          {$unsigned(reg4691)} : (forvar4670[(4'h8):(2'h2)] >= $unsigned(reg4682))));
                    end
                  reg4699 <= (|reg4617[(1'h1):(1'h1)]);
                  for (forvar4700 = (1'h0); (forvar4700 < (1'h0)); forvar4700 = (forvar4700 + (1'h1)))
                    begin
                      reg4701 <= reg4565[(1'h0):(1'h0)];
                      reg4702 <= reg4658;
                    end
                  if (($signed($signed(reg3919[(3'h4):(3'h4)])) ?
                      ({$unsigned(reg4553)} & {wire4542}) : $signed(wire3935[(3'h4):(1'h0)])))
                    begin
                      reg4703 <= $signed(reg4698);
                      reg4704 <= ((reg4676 ?
                              (~^reg4638[(1'h1):(1'h0)]) : $unsigned($unsigned(reg4619))) ?
                          (~|$signed((reg4660 || reg4697))) : (~|((reg4570 ?
                                  reg4592 : (8'hba)) ?
                              $signed(reg4698) : reg3926[(4'hb):(3'h7)])));
                      reg4705 <= $signed({(wire4583 ?
                              (reg4673 ? (8'hb6) : (8'h9d)) : (reg4687 ?
                                  reg3919 : reg4704))});
                    end
                  else
                    begin
                      reg4703 <= $signed((~^reg3928[(1'h1):(1'h1)]));
                    end
                end
              else
                begin
                  reg4694 <= reg4601;
                  reg4695 <= $signed((8'ha2));
                  if ({$unsigned((reg4594 ?
                          (reg3918 ? reg4682 : forvar4662) : (reg4672 ?
                              reg4654 : wire3903)))})
                    begin
                      reg4696 <= (^(~$signed(wire3904[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg4696 <= reg4567;
                      reg4697 <= (^$unsigned({reg4622[(1'h1):(1'h0)]}));
                    end
                  reg4698 <= reg4592[(3'h5):(2'h3)];
                end
              reg4706 <= forvar4652[(1'h1):(1'h0)];
              if ($signed(($signed((|reg4681)) ?
                  ($unsigned(forvar4687) >> reg4660) : ($signed(forvar4672) ?
                      $unsigned(forvar4649) : (reg4704 ? reg4690 : reg4701)))))
                begin
                  reg4707 <= reg4613[(2'h3):(1'h1)];
                  reg4708 <= reg4700[(4'h8):(2'h3)];
                  if ($unsigned((~^(reg4634[(1'h0):(1'h0)] ?
                      (reg3929 - reg3931) : reg4665[(1'h1):(1'h0)]))))
                    begin
                      reg4709 <= (reg4656 ^ {$unsigned($unsigned(reg3923))});
                      reg4710 <= ($unsigned((reg4697[(3'h5):(2'h2)] ?
                          reg4695 : ((8'ha7) && reg4556))) == reg4561[(3'h6):(3'h5)]);
                    end
                  else
                    begin
                      reg4709 <= ($signed({$unsigned((8'hb6))}) < (reg4575[(1'h0):(1'h0)] & reg3922[(1'h1):(1'h0)]));
                      reg4710 <= (~^$signed($unsigned({(8'hb7)})));
                      reg4711 <= ((!(-reg4610)) ?
                          $signed((((8'hae) ? forvar4670 : reg4704) ?
                              (reg4634 ^~ (8'hb6)) : {reg4654})) : wire4544[(1'h1):(1'h0)]);
                    end
                  if ({(-$signed(reg4656[(3'h6):(2'h3)]))})
                    begin
                      reg4712 <= reg4658;
                      reg4713 <= (($unsigned($signed(forvar4672)) != forvar4669[(1'h0):(1'h0)]) * (($signed((8'hb6)) << reg4621[(2'h3):(1'h1)]) == (^$signed(reg4670))));
                      reg4714 <= reg4607[(4'h9):(3'h5)];
                      reg4715 <= forvar4665[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg4712 <= reg4552;
                      reg4713 <= reg4684;
                    end
                end
              else
                begin
                  if ($signed($unsigned((reg4571 ?
                      (forvar4700 ? reg4599 : reg4685) : $signed((8'hac))))))
                    begin
                      reg4707 <= (^(~^$unsigned((^reg4599))));
                    end
                  else
                    begin
                      reg4707 <= $unsigned($unsigned(($signed(reg4563) ^ (wire4544 ?
                          reg4575 : reg4578))));
                      reg4708 <= (~$unsigned(forvar4687[(4'hb):(3'h6)]));
                      reg4709 <= $signed((8'hb4));
                      reg4710 <= {$unsigned({(reg4675 - reg3910)})};
                    end
                  reg4711 <= reg4681[(3'h5):(1'h1)];
                end
            end
          for (forvar4716 = (1'h0); (forvar4716 < (1'h0)); forvar4716 = (forvar4716 + (1'h1)))
            begin
              reg4717 <= wire4539;
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3414  (y, clk, wire3415, wire3416, wire3417, wire3418, wire3419);
  output wire [(32'h7e6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire3415;
  input wire [(5'h10):(1'h0)] wire3416;
  input wire signed [(4'hc):(1'h0)] wire3417;
  input wire [(5'h10):(1'h0)] wire3418;
  input wire signed [(4'hd):(1'h0)] wire3419;
  wire [(4'hf):(1'h0)] wire3897;
  wire [(3'h6):(1'h0)] wire3896;
  wire signed [(4'ha):(1'h0)] wire3895;
  wire signed [(3'h5):(1'h0)] wire3894;
  wire [(4'ha):(1'h0)] wire3829;
  wire signed [(2'h3):(1'h0)] wire3828;
  wire signed [(4'hf):(1'h0)] wire3420;
  wire [(4'he):(1'h0)] wire3714;
  reg [(2'h3):(1'h0)] reg3893 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3892 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3891 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3890 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3889 = (1'h0);
  reg [(2'h3):(1'h0)] reg3887 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3885 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3884 = (1'h0);
  reg [(2'h2):(1'h0)] reg3883 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3881 = (1'h0);
  reg [(4'h8):(1'h0)] reg3880 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3879 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3878 = (1'h0);
  reg [(4'h9):(1'h0)] reg3872 = (1'h0);
  reg [(4'hf):(1'h0)] reg3877 = (1'h0);
  reg [(4'h8):(1'h0)] reg3875 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3874 = (1'h0);
  reg [(4'hc):(1'h0)] reg3873 = (1'h0);
  reg [(3'h5):(1'h0)] reg3867 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3863 = (1'h0);
  reg [(4'h8):(1'h0)] reg3856 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3845 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3832 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3871 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3870 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3869 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3868 = (1'h0);
  reg [(2'h2):(1'h0)] reg3866 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3865 = (1'h0);
  reg [(4'h8):(1'h0)] reg3864 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3862 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3861 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3860 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3859 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3857 = (1'h0);
  reg [(2'h2):(1'h0)] reg3841 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3836 = (1'h0);
  reg [(4'ha):(1'h0)] reg3830 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3853 = (1'h0);
  reg [(3'h5):(1'h0)] reg3851 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3855 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3854 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3852 = (1'h0);
  reg [(3'h7):(1'h0)] reg3850 = (1'h0);
  reg [(3'h6):(1'h0)] reg3849 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3848 = (1'h0);
  reg [(4'hd):(1'h0)] reg3847 = (1'h0);
  reg [(4'hb):(1'h0)] reg3846 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3844 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3843 = (1'h0);
  reg [(3'h5):(1'h0)] reg3842 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3840 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3839 = (1'h0);
  reg [(4'hb):(1'h0)] reg3838 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3837 = (1'h0);
  reg [(2'h2):(1'h0)] reg3835 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3834 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3833 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3831 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3827 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3826 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3824 = (1'h0);
  reg [(4'hb):(1'h0)] reg3823 = (1'h0);
  reg [(4'ha):(1'h0)] reg3822 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3821 = (1'h0);
  reg [(3'h7):(1'h0)] reg3820 = (1'h0);
  reg [(4'hc):(1'h0)] reg3818 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3817 = (1'h0);
  reg [(4'h9):(1'h0)] reg3816 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3815 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3814 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3813 = (1'h0);
  reg [(2'h2):(1'h0)] reg3812 = (1'h0);
  reg [(4'he):(1'h0)] reg3811 = (1'h0);
  reg [(3'h7):(1'h0)] reg3781 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3809 = (1'h0);
  reg [(4'hf):(1'h0)] reg3808 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3807 = (1'h0);
  reg [(4'hd):(1'h0)] reg3806 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3804 = (1'h0);
  reg [(4'hf):(1'h0)] reg3803 = (1'h0);
  reg [(4'hc):(1'h0)] reg3802 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3801 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3800 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3799 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3798 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3789 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3796 = (1'h0);
  reg [(3'h6):(1'h0)] reg3795 = (1'h0);
  reg [(4'h8):(1'h0)] reg3794 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3793 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3792 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3791 = (1'h0);
  reg [(2'h3):(1'h0)] reg3790 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3788 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3787 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3785 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3784 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3783 = (1'h0);
  reg [(4'hf):(1'h0)] reg3780 = (1'h0);
  reg [(4'hb):(1'h0)] reg3778 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3777 = (1'h0);
  reg [(5'h10):(1'h0)] reg3775 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3774 = (1'h0);
  reg [(3'h4):(1'h0)] reg3773 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3772 = (1'h0);
  reg [(2'h3):(1'h0)] reg3771 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3769 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3766 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3764 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3762 = (1'h0);
  reg [(3'h6):(1'h0)] reg3761 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3760 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3759 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3758 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3757 = (1'h0);
  reg [(3'h5):(1'h0)] reg3756 = (1'h0);
  reg [(3'h6):(1'h0)] reg3755 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3754 = (1'h0);
  reg [(4'hf):(1'h0)] reg3752 = (1'h0);
  reg [(4'ha):(1'h0)] reg3751 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3749 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3748 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3747 = (1'h0);
  reg [(5'h10):(1'h0)] reg3745 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3742 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3741 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3740 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3739 = (1'h0);
  reg [(4'he):(1'h0)] reg3738 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3737 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3736 = (1'h0);
  reg [(4'hb):(1'h0)] reg3735 = (1'h0);
  reg [(4'hf):(1'h0)] reg3734 = (1'h0);
  reg [(5'h10):(1'h0)] reg3733 = (1'h0);
  reg [(3'h7):(1'h0)] reg3731 = (1'h0);
  reg [(3'h4):(1'h0)] reg3729 = (1'h0);
  reg [(4'hd):(1'h0)] reg3727 = (1'h0);
  reg [(4'h8):(1'h0)] reg3723 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3721 = (1'h0);
  reg [(4'hf):(1'h0)] reg3728 = (1'h0);
  reg [(4'ha):(1'h0)] reg3726 = (1'h0);
  reg [(4'ha):(1'h0)] reg3725 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3724 = (1'h0);
  reg [(4'hf):(1'h0)] reg3722 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3720 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3719 = (1'h0);
  reg [(3'h5):(1'h0)] reg3718 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3717 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3716 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3888 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3886 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3882 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3875 = (1'h0);
  reg [(4'he):(1'h0)] forvar3871 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3870 = (1'h0);
  reg [(4'he):(1'h0)] forvar3865 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3876 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3872 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3869 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3866 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3848 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3834 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3849 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3846 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3831 = (1'h0);
  reg [(4'he):(1'h0)] forvar3867 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3863 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3858 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3856 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3837 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3850 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3853 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3851 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3845 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3841 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3836 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3832 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3830 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3825 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3819 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3812 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3810 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3805 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3797 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3792 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3789 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3786 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3782 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3781 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3779 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3776 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3770 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3768 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3767 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3765 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3763 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3755 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3753 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3750 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3746 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3744 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3743 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3732 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3730 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3725 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3719 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3717 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3727 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3723 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3721 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3716 = (1'h0);
  assign y = {wire3897,
                 wire3896,
                 wire3895,
                 wire3894,
                 wire3829,
                 wire3828,
                 wire3420,
                 wire3714,
                 reg3893,
                 reg3892,
                 reg3891,
                 reg3890,
                 reg3889,
                 reg3887,
                 reg3885,
                 reg3884,
                 reg3883,
                 reg3881,
                 reg3880,
                 reg3879,
                 reg3878,
                 reg3872,
                 reg3877,
                 reg3875,
                 reg3874,
                 reg3873,
                 reg3867,
                 reg3863,
                 reg3856,
                 reg3845,
                 reg3832,
                 reg3871,
                 reg3870,
                 reg3869,
                 reg3868,
                 reg3866,
                 reg3865,
                 reg3864,
                 reg3862,
                 reg3861,
                 reg3860,
                 reg3859,
                 reg3857,
                 reg3841,
                 reg3836,
                 reg3830,
                 reg3853,
                 reg3851,
                 reg3855,
                 reg3854,
                 reg3852,
                 reg3850,
                 reg3849,
                 reg3848,
                 reg3847,
                 reg3846,
                 reg3844,
                 reg3843,
                 reg3842,
                 reg3840,
                 reg3839,
                 reg3838,
                 reg3837,
                 reg3835,
                 reg3834,
                 reg3833,
                 reg3831,
                 reg3827,
                 reg3826,
                 reg3824,
                 reg3823,
                 reg3822,
                 reg3821,
                 reg3820,
                 reg3818,
                 reg3817,
                 reg3816,
                 reg3815,
                 reg3814,
                 reg3813,
                 reg3812,
                 reg3811,
                 reg3781,
                 reg3809,
                 reg3808,
                 reg3807,
                 reg3806,
                 reg3804,
                 reg3803,
                 reg3802,
                 reg3801,
                 reg3800,
                 reg3799,
                 reg3798,
                 reg3789,
                 reg3796,
                 reg3795,
                 reg3794,
                 reg3793,
                 reg3792,
                 reg3791,
                 reg3790,
                 reg3788,
                 reg3787,
                 reg3785,
                 reg3784,
                 reg3783,
                 reg3780,
                 reg3778,
                 reg3777,
                 reg3775,
                 reg3774,
                 reg3773,
                 reg3772,
                 reg3771,
                 reg3769,
                 reg3766,
                 reg3764,
                 reg3762,
                 reg3761,
                 reg3760,
                 reg3759,
                 reg3758,
                 reg3757,
                 reg3756,
                 reg3755,
                 reg3754,
                 reg3752,
                 reg3751,
                 reg3749,
                 reg3748,
                 reg3747,
                 reg3745,
                 reg3742,
                 reg3741,
                 reg3740,
                 reg3739,
                 reg3738,
                 reg3737,
                 reg3736,
                 reg3735,
                 reg3734,
                 reg3733,
                 reg3731,
                 reg3729,
                 reg3727,
                 reg3723,
                 reg3721,
                 reg3728,
                 reg3726,
                 reg3725,
                 reg3724,
                 reg3722,
                 reg3720,
                 reg3719,
                 reg3718,
                 reg3717,
                 reg3716,
                 forvar3888,
                 forvar3886,
                 forvar3882,
                 forvar3875,
                 forvar3871,
                 forvar3870,
                 forvar3865,
                 forvar3876,
                 forvar3872,
                 forvar3869,
                 forvar3866,
                 forvar3848,
                 forvar3834,
                 forvar3849,
                 forvar3846,
                 forvar3831,
                 forvar3867,
                 forvar3863,
                 forvar3858,
                 forvar3856,
                 forvar3837,
                 forvar3850,
                 forvar3853,
                 forvar3851,
                 forvar3845,
                 forvar3841,
                 forvar3836,
                 forvar3832,
                 forvar3830,
                 forvar3825,
                 forvar3819,
                 forvar3812,
                 forvar3810,
                 forvar3805,
                 forvar3797,
                 forvar3792,
                 forvar3789,
                 forvar3786,
                 forvar3782,
                 forvar3781,
                 forvar3779,
                 forvar3776,
                 forvar3770,
                 forvar3768,
                 forvar3767,
                 forvar3765,
                 forvar3763,
                 forvar3755,
                 forvar3753,
                 forvar3750,
                 forvar3746,
                 forvar3744,
                 forvar3743,
                 forvar3732,
                 forvar3730,
                 forvar3725,
                 forvar3719,
                 forvar3717,
                 forvar3727,
                 forvar3723,
                 forvar3721,
                 forvar3716,
                 (1'h0)};
  assign wire3420 = ($signed(((|wire3418) - (wire3419 < (8'had)))) ?
                        {$unsigned(wire3415[(3'h5):(3'h5)])} : wire3415[(3'h5):(1'h1)]);
  module3421 #() modinst3715 (.clk(clk), .wire3425(wire3417), .wire3423(wire3420), .wire3424(wire3419), .wire3426(wire3415), .y(wire3714), .wire3422(wire3418));
  always
    @(posedge clk) begin
      if (wire3419[(3'h6):(3'h5)])
        begin
          reg3716 <= (~($signed((wire3416 ^~ wire3416)) == wire3420[(1'h1):(1'h1)]));
        end
      else
        begin
          for (forvar3716 = (1'h0); (forvar3716 < (2'h2)); forvar3716 = (forvar3716 + (1'h1)))
            begin
              if ((wire3418 < (forvar3716[(2'h2):(2'h2)] ?
                  wire3714 : {(wire3420 ? wire3416 : wire3419)})))
                begin
                  if (($unsigned((wire3419[(2'h3):(2'h3)] + wire3415[(3'h5):(3'h4)])) ?
                      reg3716[(2'h2):(1'h0)] : wire3418))
                    begin
                      reg3717 <= ($signed(((forvar3716 ? wire3415 : wire3416) ?
                              wire3415 : wire3418[(4'hc):(2'h3)])) ?
                          wire3417 : (|(^~wire3417[(2'h2):(2'h2)])));
                      reg3718 <= forvar3716[(1'h1):(1'h0)];
                      reg3719 <= wire3714[(4'hb):(3'h4)];
                    end
                  else
                    begin
                      reg3717 <= ((|($signed(reg3719) ?
                          (wire3418 >> (8'hb5)) : forvar3716[(1'h1):(1'h0)])) != ((8'h9e) << ((wire3417 | reg3716) ?
                          (&forvar3716) : wire3714[(1'h0):(1'h0)])));
                      reg3718 <= reg3717[(3'h7):(2'h3)];
                      reg3719 <= reg3717[(3'h5):(1'h1)];
                      reg3720 <= reg3718;
                    end
                  for (forvar3721 = (1'h0); (forvar3721 < (1'h0)); forvar3721 = (forvar3721 + (1'h1)))
                    begin
                      reg3722 <= (~|(|{(reg3719 ? forvar3716 : wire3714)}));
                    end
                  for (forvar3723 = (1'h0); (forvar3723 < (2'h2)); forvar3723 = (forvar3723 + (1'h1)))
                    begin
                      reg3724 <= $unsigned((^~($signed(wire3417) <= {wire3417})));
                      reg3725 <= ($unsigned(reg3716[(3'h7):(3'h5)]) ?
                          (8'haf) : (~^wire3415[(4'h8):(2'h3)]));
                      reg3726 <= (reg3718 ?
                          (!($signed(reg3724) ?
                              wire3418 : forvar3721[(4'he):(2'h3)])) : ((forvar3716 <<< (!wire3415)) ?
                              $signed(wire3417[(4'hb):(4'h8)]) : reg3716[(3'h5):(2'h3)]));
                    end
                  for (forvar3727 = (1'h0); (forvar3727 < (2'h3)); forvar3727 = (forvar3727 + (1'h1)))
                    begin
                      reg3728 <= $signed($unsigned(((wire3417 >>> wire3415) >= wire3415[(2'h3):(1'h1)])));
                    end
                end
              else
                begin
                  for (forvar3717 = (1'h0); (forvar3717 < (1'h0)); forvar3717 = (forvar3717 + (1'h1)))
                    begin
                      reg3718 <= {$unsigned((~^(~^reg3718)))};
                    end
                  for (forvar3719 = (1'h0); (forvar3719 < (1'h1)); forvar3719 = (forvar3719 + (1'h1)))
                    begin
                      reg3720 <= forvar3721;
                      reg3721 <= {$unsigned($signed((!wire3416)))};
                      reg3722 <= {(forvar3721 ?
                              (reg3722 ?
                                  ((8'hb2) ?
                                      wire3415 : reg3726) : $signed(reg3718)) : wire3417)};
                      reg3723 <= $unsigned(($unsigned(forvar3721) | ((8'hb8) ?
                          reg3719[(4'ha):(2'h3)] : (wire3415 ^~ reg3725))));
                    end
                  reg3724 <= $unsigned((((!reg3723) ?
                          reg3722 : wire3419[(3'h6):(1'h0)]) ?
                      reg3720 : (wire3714 ?
                          (reg3718 - wire3417) : (|(8'ha6)))));
                  for (forvar3725 = (1'h0); (forvar3725 < (2'h2)); forvar3725 = (forvar3725 + (1'h1)))
                    begin
                      reg3726 <= forvar3727[(4'h8):(4'h8)];
                      reg3727 <= (^(+{reg3719[(1'h0):(1'h0)]}));
                    end
                end
              if ($unsigned((($signed(forvar3716) || {forvar3719}) ?
                  {reg3716} : $unsigned((wire3416 ? (8'haf) : reg3722)))))
                begin
                  reg3729 <= {forvar3717};
                end
              else
                begin
                  reg3729 <= $signed((((forvar3716 != (8'ha0)) > $unsigned(wire3714)) <= reg3723));
                end
              for (forvar3730 = (1'h0); (forvar3730 < (1'h0)); forvar3730 = (forvar3730 + (1'h1)))
                begin
                  reg3731 <= {(8'ha6)};
                  for (forvar3732 = (1'h0); (forvar3732 < (2'h2)); forvar3732 = (forvar3732 + (1'h1)))
                    begin
                      reg3733 <= ((~{reg3726}) >> reg3728[(3'h6):(1'h1)]);
                      reg3734 <= (8'ha4);
                      reg3735 <= $unsigned({$unsigned((+forvar3732))});
                      reg3736 <= reg3718[(2'h3):(2'h3)];
                    end
                  if ((^((|(wire3416 >= reg3726)) ~^ $signed(reg3735[(3'h7):(1'h1)]))))
                    begin
                      reg3737 <= reg3720[(4'hb):(1'h0)];
                      reg3738 <= reg3735[(3'h7):(2'h3)];
                      reg3739 <= reg3724;
                      reg3740 <= $signed($signed({(wire3420 == (8'h9c))}));
                    end
                  else
                    begin
                      reg3737 <= (!$unsigned($signed(forvar3716[(1'h0):(1'h0)])));
                      reg3738 <= forvar3723[(2'h2):(1'h1)];
                      reg3739 <= (8'ha8);
                      reg3740 <= $signed(reg3723[(2'h3):(2'h2)]);
                    end
                  reg3741 <= reg3729[(3'h4):(1'h0)];
                end
            end
          reg3742 <= (reg3724[(4'h8):(4'h8)] ?
              (((8'h9e) ?
                  (reg3733 ?
                      wire3714 : reg3727) : $unsigned(forvar3732)) != (8'hae)) : $signed($signed($signed(forvar3721))));
          for (forvar3743 = (1'h0); (forvar3743 < (2'h2)); forvar3743 = (forvar3743 + (1'h1)))
            begin
              for (forvar3744 = (1'h0); (forvar3744 < (1'h1)); forvar3744 = (forvar3744 + (1'h1)))
                begin
                  reg3745 <= wire3420;
                  for (forvar3746 = (1'h0); (forvar3746 < (2'h3)); forvar3746 = (forvar3746 + (1'h1)))
                    begin
                      reg3747 <= ((8'ha8) == {{$signed(wire3415)}});
                      reg3748 <= $signed({$unsigned(forvar3725[(1'h1):(1'h1)])});
                      reg3749 <= forvar3730[(3'h5):(2'h2)];
                    end
                  for (forvar3750 = (1'h0); (forvar3750 < (1'h0)); forvar3750 = (forvar3750 + (1'h1)))
                    begin
                      reg3751 <= forvar3743[(4'ha):(1'h1)];
                      reg3752 <= reg3751[(4'h8):(3'h6)];
                    end
                end
              for (forvar3753 = (1'h0); (forvar3753 < (2'h2)); forvar3753 = (forvar3753 + (1'h1)))
                begin
                  reg3754 <= ((^((forvar3730 << reg3717) ?
                      reg3748[(1'h1):(1'h1)] : reg3741)) ~^ reg3727[(3'h6):(3'h6)]);
                end
              if (($signed(reg3724) ? (&forvar3723[(2'h2):(1'h0)]) : reg3722))
                begin
                  if ((reg3734[(1'h0):(1'h0)] ?
                      reg3742[(1'h0):(1'h0)] : $unsigned({(reg3754 << wire3420)})))
                    begin
                      reg3755 <= (reg3741[(4'h9):(4'h8)] <= $signed(($unsigned(reg3717) ?
                          reg3749[(2'h2):(1'h1)] : $signed(wire3418))));
                      reg3756 <= ((~|(~&(^~reg3755))) || $unsigned(reg3735[(3'h5):(3'h4)]));
                      reg3757 <= $unsigned((($unsigned(wire3714) != $unsigned((8'haf))) <<< (|$signed(reg3721))));
                    end
                  else
                    begin
                      reg3755 <= (&$signed((~(reg3716 ? reg3723 : wire3714))));
                    end
                  if (({((forvar3732 & reg3742) ? reg3728 : {wire3416})} ?
                      reg3751[(4'h8):(4'h8)] : (forvar3732[(2'h3):(1'h1)] | (^$signed(reg3734)))))
                    begin
                      reg3758 <= (($unsigned((8'hb2)) - $signed((reg3723 ?
                              (8'ha2) : wire3714))) ?
                          (^~(wire3419 - reg3741[(4'hc):(3'h7)])) : (!reg3723[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg3758 <= (|reg3726);
                    end
                  if ($signed($unsigned((reg3741 ?
                      reg3758[(2'h3):(1'h1)] : $signed(wire3418)))))
                    begin
                      reg3759 <= {(!(!(forvar3727 ? forvar3753 : reg3748)))};
                      reg3760 <= $signed($signed(($unsigned(forvar3721) ?
                          (!reg3756) : $signed(reg3738))));
                    end
                  else
                    begin
                      reg3759 <= $unsigned((({reg3745} ?
                          {(8'ha2)} : ((8'hac) ?
                              forvar3750 : forvar3743)) * $signed((reg3741 ?
                          reg3759 : (8'hb6)))));
                    end
                  reg3761 <= $unsigned(((reg3720[(4'he):(1'h0)] && reg3740) ?
                      {$signed(reg3723)} : (wire3415 ^ (reg3741 <<< reg3752))));
                end
              else
                begin
                  for (forvar3755 = (1'h0); (forvar3755 < (2'h3)); forvar3755 = (forvar3755 + (1'h1)))
                    begin
                      reg3756 <= forvar3723;
                    end
                  if (reg3729)
                    begin
                      reg3757 <= ({(^~{reg3727})} + (^~$unsigned((reg3754 ?
                          forvar3727 : wire3419))));
                      reg3758 <= (reg3759[(3'h5):(2'h2)] ?
                          {$unsigned(reg3758)} : $unsigned((~reg3740[(1'h0):(1'h0)])));
                      reg3759 <= ((~|reg3737) || $signed(reg3727));
                      reg3760 <= $unsigned(($unsigned((reg3738 ?
                              reg3719 : forvar3727)) ?
                          $unsigned(reg3719) : $unsigned($unsigned(reg3725))));
                    end
                  else
                    begin
                      reg3757 <= reg3728;
                    end
                  if (({((^forvar3723) + $unsigned(reg3759))} >> reg3756[(1'h1):(1'h0)]))
                    begin
                      reg3761 <= $unsigned(wire3418);
                      reg3762 <= $unsigned((~reg3733[(4'h8):(2'h3)]));
                    end
                  else
                    begin
                      reg3761 <= $signed(($unsigned((forvar3730 <= forvar3721)) << reg3755));
                    end
                  for (forvar3763 = (1'h0); (forvar3763 < (1'h0)); forvar3763 = (forvar3763 + (1'h1)))
                    begin
                      reg3764 <= (8'hb8);
                    end
                end
            end
        end
      for (forvar3765 = (1'h0); (forvar3765 < (2'h2)); forvar3765 = (forvar3765 + (1'h1)))
        begin
          reg3766 <= $unsigned($unsigned((forvar3723[(1'h0):(1'h0)] * {(8'ha5)})));
          for (forvar3767 = (1'h0); (forvar3767 < (2'h2)); forvar3767 = (forvar3767 + (1'h1)))
            begin
              for (forvar3768 = (1'h0); (forvar3768 < (1'h0)); forvar3768 = (forvar3768 + (1'h1)))
                begin
                  reg3769 <= (|($unsigned((forvar3723 & reg3759)) >> reg3726));
                end
              for (forvar3770 = (1'h0); (forvar3770 < (1'h0)); forvar3770 = (forvar3770 + (1'h1)))
                begin
                  if (({((wire3418 >>> (8'haa)) ? {(8'hb9)} : (~&forvar3743))} ?
                      (wire3419 ?
                          $signed((forvar3765 ?
                              forvar3717 : (8'hb3))) : $unsigned($unsigned((8'hb3)))) : forvar3770))
                    begin
                      reg3771 <= $signed($unsigned({{reg3755}}));
                      reg3772 <= ($signed(reg3731[(1'h1):(1'h0)]) < $unsigned(reg3760));
                    end
                  else
                    begin
                      reg3771 <= $signed($unsigned((~(|reg3764))));
                      reg3772 <= $unsigned(((reg3739 ?
                          (reg3738 ?
                              (8'hb2) : (8'hb7)) : (forvar3765 < reg3737)) ^ $unsigned(reg3726[(1'h0):(1'h0)])));
                    end
                  if ((~&(reg3737 >> $signed((forvar3763 && forvar3765)))))
                    begin
                      reg3773 <= (8'ha6);
                      reg3774 <= (($unsigned((forvar3753 == reg3721)) ?
                              reg3722 : $unsigned((|reg3734))) ?
                          (~^((!forvar3727) >= reg3734)) : ((~reg3725[(2'h2):(1'h0)]) ^~ $signed((reg3724 ^ wire3415))));
                      reg3775 <= reg3757;
                    end
                  else
                    begin
                      reg3773 <= reg3733[(2'h3):(2'h2)];
                      reg3774 <= (($signed((~&(8'ha3))) >= ((reg3775 == reg3736) < (reg3769 ?
                              (8'ha3) : (8'ha5)))) ?
                          reg3749[(1'h0):(1'h0)] : {(reg3747[(3'h7):(2'h3)] && $unsigned(forvar3746))});
                    end
                end
              for (forvar3776 = (1'h0); (forvar3776 < (2'h3)); forvar3776 = (forvar3776 + (1'h1)))
                begin
                  if ((^reg3771))
                    begin
                      reg3777 <= $signed(($signed((reg3760 ?
                          forvar3719 : reg3725)) >> ($signed(reg3761) ?
                          (!forvar3763) : (reg3772 ? (8'haa) : reg3725))));
                    end
                  else
                    begin
                      reg3777 <= (reg3733[(5'h10):(4'he)] ?
                          $signed(reg3737[(1'h0):(1'h0)]) : reg3721);
                    end
                end
            end
        end
      reg3778 <= reg3749[(2'h3):(1'h0)];
      for (forvar3779 = (1'h0); (forvar3779 < (2'h2)); forvar3779 = (forvar3779 + (1'h1)))
        begin
          reg3780 <= $unsigned({(&reg3766[(3'h5):(1'h1)])});
          if ((forvar3716 ? forvar3779[(3'h6):(1'h1)] : $signed(reg3773)))
            begin
              for (forvar3781 = (1'h0); (forvar3781 < (2'h3)); forvar3781 = (forvar3781 + (1'h1)))
                begin
                  for (forvar3782 = (1'h0); (forvar3782 < (2'h3)); forvar3782 = (forvar3782 + (1'h1)))
                    begin
                      reg3783 <= (~^$unsigned((~&$signed((8'hba)))));
                      reg3784 <= reg3722[(4'he):(4'he)];
                    end
                  reg3785 <= (forvar3782 ?
                      (!((reg3720 * forvar3730) - $signed(reg3734))) : reg3752);
                  for (forvar3786 = (1'h0); (forvar3786 < (1'h1)); forvar3786 = (forvar3786 + (1'h1)))
                    begin
                      reg3787 <= $unsigned($unsigned((&(~forvar3730))));
                      reg3788 <= ({({forvar3767} ?
                              (reg3772 <<< forvar3776) : $signed(reg3773))} > (-((8'ha9) ?
                          reg3761 : reg3734[(1'h0):(1'h0)])));
                    end
                end
              if (reg3721[(1'h0):(1'h0)])
                begin
                  for (forvar3789 = (1'h0); (forvar3789 < (2'h2)); forvar3789 = (forvar3789 + (1'h1)))
                    begin
                      reg3790 <= ({$signed(((8'hb0) * reg3780))} > ($unsigned({reg3740}) == wire3418));
                      reg3791 <= $signed(reg3726);
                      reg3792 <= (reg3760[(2'h2):(1'h0)] != reg3791);
                    end
                  if ($unsigned(forvar3717[(3'h4):(2'h2)]))
                    begin
                      reg3793 <= $signed(forvar3755[(1'h1):(1'h0)]);
                      reg3794 <= reg3769[(4'h9):(1'h1)];
                      reg3795 <= $unsigned(forvar3781[(1'h0):(1'h0)]);
                      reg3796 <= (|forvar3732[(3'h6):(1'h1)]);
                    end
                  else
                    begin
                      reg3793 <= reg3745;
                      reg3794 <= $signed(reg3755[(3'h6):(2'h2)]);
                      reg3795 <= {$unsigned(($signed(wire3418) ?
                              (reg3737 & forvar3753) : reg3747))};
                      reg3796 <= ((($signed(forvar3779) ~^ reg3795[(1'h1):(1'h0)]) >>> (^{reg3721})) >>> ((reg3780 ?
                          (reg3793 ?
                              forvar3786 : reg3762) : (forvar3743 && forvar3721)) * reg3785[(2'h2):(2'h2)]));
                    end
                end
              else
                begin
                  if (((({reg3791} ?
                      (reg3716 * reg3721) : $signed(reg3760)) == reg3757) >> (($signed(reg3723) ?
                      $unsigned(reg3736) : $unsigned(reg3719)) >= reg3757[(4'he):(1'h0)])))
                    begin
                      reg3789 <= {forvar3781};
                      reg3790 <= {(~$signed(reg3791))};
                      reg3791 <= $signed(((&(+forvar3746)) < (&(8'hb6))));
                    end
                  else
                    begin
                      reg3789 <= {forvar3779};
                    end
                  for (forvar3792 = (1'h0); (forvar3792 < (1'h0)); forvar3792 = (forvar3792 + (1'h1)))
                    begin
                      reg3793 <= reg3738[(4'hb):(3'h6)];
                      reg3794 <= (-{reg3735[(2'h2):(2'h2)]});
                      reg3795 <= $signed(($unsigned({reg3719}) ?
                          (~^((8'haa) == (8'h9f))) : reg3747[(2'h3):(1'h1)]));
                      reg3796 <= $unsigned({(~|$unsigned(reg3754))});
                    end
                end
              for (forvar3797 = (1'h0); (forvar3797 < (1'h0)); forvar3797 = (forvar3797 + (1'h1)))
                begin
                  if ($unsigned(reg3783[(2'h2):(1'h0)]))
                    begin
                      reg3798 <= reg3736[(4'hb):(1'h0)];
                    end
                  else
                    begin
                      reg3798 <= $signed(reg3717);
                      reg3799 <= {forvar3716[(2'h2):(1'h1)]};
                      reg3800 <= reg3774[(1'h1):(1'h0)];
                    end
                  if (($signed(((reg3778 ^ reg3728) << forvar3725)) ?
                      reg3798 : (~(^(forvar3744 | reg3764)))))
                    begin
                      reg3801 <= (+(wire3416 ? {reg3723} : $unsigned((8'ha5))));
                      reg3802 <= (-($signed($signed(wire3420)) * $signed({reg3784})));
                      reg3803 <= {$signed(reg3752)};
                      reg3804 <= (($unsigned(reg3745) >> reg3761) ?
                          reg3739[(4'ha):(1'h0)] : ({(reg3733 >= reg3778)} <<< $signed(forvar3717)));
                    end
                  else
                    begin
                      reg3801 <= $signed(forvar3725[(1'h0):(1'h0)]);
                    end
                  for (forvar3805 = (1'h0); (forvar3805 < (1'h1)); forvar3805 = (forvar3805 + (1'h1)))
                    begin
                      reg3806 <= $unsigned((~|reg3742[(2'h2):(1'h0)]));
                      reg3807 <= (($unsigned(wire3420) + (8'hba)) ?
                          $unsigned((forvar3763[(3'h6):(3'h6)] ?
                              (!reg3726) : (wire3416 != reg3792))) : (reg3720 >= forvar3782[(3'h5):(1'h1)]));
                    end
                  if ({($signed((reg3734 ?
                          reg3784 : reg3759)) <<< ((+(8'hb3)) > (^~wire3417)))})
                    begin
                      reg3808 <= reg3755;
                    end
                  else
                    begin
                      reg3808 <= ((8'hb1) + (forvar3723[(1'h1):(1'h0)] == reg3726));
                      reg3809 <= ((-(~reg3727[(1'h0):(1'h0)])) ?
                          reg3749 : $unsigned(((forvar3727 << (8'had)) < forvar3725)));
                    end
                end
            end
          else
            begin
              reg3781 <= reg3717[(3'h6):(3'h5)];
            end
          for (forvar3810 = (1'h0); (forvar3810 < (1'h1)); forvar3810 = (forvar3810 + (1'h1)))
            begin
              reg3811 <= $signed(wire3420[(3'h5):(3'h5)]);
              if ($signed(((~|$signed(reg3771)) ?
                  $unsigned($unsigned((8'hab))) : {(reg3796 | (8'hba))})))
                begin
                  reg3812 <= reg3789[(2'h3):(2'h3)];
                end
              else
                begin
                  for (forvar3812 = (1'h0); (forvar3812 < (1'h1)); forvar3812 = (forvar3812 + (1'h1)))
                    begin
                      reg3813 <= $unsigned($signed((~^(reg3716 && reg3761))));
                      reg3814 <= (((reg3724[(2'h2):(2'h2)] ?
                              $unsigned((8'hb3)) : $signed(forvar3755)) ?
                          ((!forvar3789) ?
                              (~^reg3778) : ((8'hb3) ?
                                  reg3777 : reg3751)) : (~|reg3795[(3'h5):(1'h0)])) <<< (^reg3739));
                    end
                  if ((($unsigned(reg3802) ^~ ((-forvar3776) && (forvar3768 | reg3813))) ?
                      $unsigned($unsigned($unsigned((8'ha4)))) : ($unsigned(reg3735[(4'ha):(3'h7)]) << ($signed(reg3726) - $signed(reg3788)))))
                    begin
                      reg3815 <= {((~^(forvar3792 * reg3809)) ?
                              reg3733[(1'h0):(1'h0)] : (forvar3753[(4'hd):(1'h0)] & $unsigned(reg3780)))};
                      reg3816 <= $unsigned($signed($unsigned((8'haa))));
                      reg3817 <= $signed(($unsigned(reg3727[(3'h4):(2'h3)]) ?
                          reg3798[(1'h1):(1'h1)] : reg3725[(4'h8):(3'h5)]));
                    end
                  else
                    begin
                      reg3815 <= {$signed($unsigned((reg3745 ?
                              forvar3716 : wire3415)))};
                      reg3816 <= $unsigned($unsigned($unsigned((+(8'ha1)))));
                    end
                end
              reg3818 <= {((((8'haf) == (8'hba)) == (reg3717 + wire3416)) ~^ $unsigned(forvar3812[(4'h9):(3'h7)]))};
              for (forvar3819 = (1'h0); (forvar3819 < (2'h3)); forvar3819 = (forvar3819 + (1'h1)))
                begin
                  reg3820 <= ((($unsigned(forvar3789) ?
                          ((8'ha4) ~^ (8'haa)) : (reg3751 ?
                              reg3802 : forvar3781)) ?
                      (reg3741[(3'h5):(3'h4)] ?
                          reg3720 : {(8'ha4)}) : (+(wire3419 ?
                          reg3725 : (8'ha3)))) && ((^(forvar3727 ?
                          reg3752 : reg3764)) ?
                      (+(reg3760 ? reg3729 : forvar3725)) : reg3740));
                  if (({$unsigned(forvar3819[(2'h3):(2'h3)])} ?
                      (8'hb4) : $signed(reg3816)))
                    begin
                      reg3821 <= reg3748[(2'h2):(1'h1)];
                      reg3822 <= (~|reg3727[(2'h3):(2'h3)]);
                      reg3823 <= reg3716[(3'h6):(1'h1)];
                      reg3824 <= ({$unsigned((!reg3718))} ?
                          reg3804[(4'h9):(3'h7)] : $signed($signed(((8'ha0) ?
                              forvar3744 : reg3735))));
                    end
                  else
                    begin
                      reg3821 <= forvar3763;
                      reg3822 <= (!forvar3819);
                      reg3823 <= reg3747;
                      reg3824 <= forvar3810[(3'h4):(1'h0)];
                    end
                end
            end
          for (forvar3825 = (1'h0); (forvar3825 < (1'h0)); forvar3825 = (forvar3825 + (1'h1)))
            begin
              reg3826 <= (8'ha9);
              reg3827 <= reg3731[(1'h0):(1'h0)];
            end
        end
    end
  assign wire3828 = reg3764;
  assign wire3829 = $unsigned((|(~^(reg3808 && (8'ha3)))));
  always
    @(posedge clk) begin
      if (($unsigned(((reg3722 | reg3735) ? (~|reg3751) : (&reg3804))) ?
          ((~$signed((8'ha0))) != $signed(reg3723)) : (reg3752 <= reg3725)))
        begin
          if ($signed({((reg3824 ? reg3724 : reg3775) ?
                  {(8'ha2)} : {reg3769})}))
            begin
              for (forvar3830 = (1'h0); (forvar3830 < (2'h2)); forvar3830 = (forvar3830 + (1'h1)))
                begin
                  reg3831 <= ((($signed(reg3747) ?
                              (!reg3800) : (wire3420 ? reg3781 : reg3793)) ?
                          {(~^reg3821)} : {reg3754[(1'h0):(1'h0)]}) ?
                      (((reg3798 ? reg3756 : reg3788) ?
                          (^reg3772) : reg3827) <= $unsigned($unsigned(reg3809))) : $unsigned(reg3822));
                end
              for (forvar3832 = (1'h0); (forvar3832 < (2'h3)); forvar3832 = (forvar3832 + (1'h1)))
                begin
                  if ({(~|($unsigned(reg3739) ? (~^reg3781) : (~reg3749)))})
                    begin
                      reg3833 <= $signed($signed(reg3814));
                      reg3834 <= ($signed($signed((&reg3831))) ?
                          ((!{reg3760}) << $signed($unsigned((8'hb8)))) : $signed({(reg3749 ?
                                  reg3820 : reg3794)}));
                      reg3835 <= (!reg3822);
                    end
                  else
                    begin
                      reg3833 <= (~^reg3811[(4'hc):(3'h4)]);
                      reg3834 <= (reg3745[(2'h3):(1'h1)] ?
                          ((((8'ha3) >> (8'haa)) < reg3724) >= reg3741) : $unsigned(reg3790[(2'h3):(1'h1)]));
                      reg3835 <= reg3739[(4'h8):(3'h7)];
                    end
                end
              for (forvar3836 = (1'h0); (forvar3836 < (2'h2)); forvar3836 = (forvar3836 + (1'h1)))
                begin
                  if ({$unsigned(({wire3419} >> {(8'h9c)}))})
                    begin
                      reg3837 <= $unsigned(($unsigned((!forvar3832)) <= $unsigned((reg3739 & reg3823))));
                      reg3838 <= (($unsigned({reg3823}) && $unsigned(((8'h9c) + (8'hac)))) ?
                          reg3742 : ({(wire3714 * (8'h9e))} ?
                              $unsigned(reg3814[(3'h5):(2'h3)]) : $unsigned(reg3727[(3'h6):(3'h6)])));
                      reg3839 <= reg3784[(3'h4):(2'h2)];
                      reg3840 <= {reg3766[(4'hd):(4'h9)]};
                    end
                  else
                    begin
                      reg3837 <= reg3833;
                    end
                  for (forvar3841 = (1'h0); (forvar3841 < (1'h1)); forvar3841 = (forvar3841 + (1'h1)))
                    begin
                      reg3842 <= (~reg3794);
                      reg3843 <= ($unsigned($unsigned({reg3751})) ?
                          (|((^reg3755) ?
                              (reg3826 ?
                                  reg3754 : reg3824) : reg3833)) : (~((reg3785 >> reg3774) + (^~reg3760))));
                      reg3844 <= (8'hb3);
                    end
                  for (forvar3845 = (1'h0); (forvar3845 < (1'h1)); forvar3845 = (forvar3845 + (1'h1)))
                    begin
                      reg3846 <= $signed(reg3795);
                      reg3847 <= reg3724[(3'h4):(2'h2)];
                      reg3848 <= (&$signed(wire3418[(3'h4):(1'h1)]));
                      reg3849 <= ($unsigned((((8'ha4) ^ reg3806) ?
                              reg3727[(3'h7):(1'h1)] : reg3839)) ?
                          ($signed((+reg3838)) ?
                              {reg3718[(1'h0):(1'h0)]} : {(reg3801 ?
                                      reg3812 : reg3754)}) : (reg3843 ?
                              ((~&reg3760) == (+reg3772)) : ((reg3728 <<< reg3725) ?
                                  (reg3817 | reg3788) : {reg3727})));
                    end
                end
              if ((reg3798 < ($signed(reg3754) == $signed((reg3725 ?
                  reg3784 : reg3716)))))
                begin
                  reg3850 <= ($unsigned($signed(reg3722[(1'h1):(1'h1)])) ?
                      $signed((^(reg3760 ?
                          reg3778 : (8'ha8)))) : (~&(+reg3807[(1'h0):(1'h0)])));
                  for (forvar3851 = (1'h0); (forvar3851 < (2'h3)); forvar3851 = (forvar3851 + (1'h1)))
                    begin
                      reg3852 <= ($unsigned({(~^reg3816)}) ^ reg3774);
                    end
                  for (forvar3853 = (1'h0); (forvar3853 < (2'h3)); forvar3853 = (forvar3853 + (1'h1)))
                    begin
                      reg3854 <= $signed(reg3741[(2'h3):(2'h3)]);
                      reg3855 <= (reg3814 > {forvar3830});
                    end
                end
              else
                begin
                  for (forvar3850 = (1'h0); (forvar3850 < (2'h3)); forvar3850 = (forvar3850 + (1'h1)))
                    begin
                      reg3851 <= (($signed(((8'hb1) == reg3760)) | reg3727[(4'hb):(3'h7)]) != $unsigned($unsigned((reg3761 ?
                          reg3790 : reg3725))));
                      reg3852 <= (^~$signed((~(wire3420 ? reg3820 : reg3783))));
                    end
                  if ((~&(^~reg3737[(1'h1):(1'h1)])))
                    begin
                      reg3853 <= $unsigned({(~^(reg3759 | reg3793))});
                    end
                  else
                    begin
                      reg3853 <= $signed(reg3848);
                      reg3854 <= ((~|$signed($unsigned(reg3783))) ?
                          ((wire3420[(1'h0):(1'h0)] ?
                              reg3747 : $signed((8'ha0))) * ((reg3784 << wire3828) ?
                              reg3762 : (reg3824 + reg3834))) : (reg3818 || ((reg3814 ?
                              reg3756 : reg3843) << (~|reg3754))));
                    end
                end
            end
          else
            begin
              reg3830 <= $unsigned(reg3814);
              reg3831 <= ($unsigned(($signed(reg3772) ?
                  (-reg3799) : (-(8'hb0)))) >>> {(reg3752[(2'h3):(1'h0)] ?
                      {reg3777} : reg3814)});
              for (forvar3832 = (1'h0); (forvar3832 < (1'h1)); forvar3832 = (forvar3832 + (1'h1)))
                begin
                  if (reg3757)
                    begin
                      reg3833 <= reg3849[(1'h1):(1'h0)];
                      reg3834 <= reg3830;
                      reg3835 <= reg3851;
                      reg3836 <= $unsigned(reg3853);
                    end
                  else
                    begin
                      reg3833 <= reg3741[(3'h4):(3'h4)];
                      reg3834 <= ((($unsigned(reg3831) ?
                                  {reg3756} : $signed(reg3760)) ?
                              $signed((~&reg3801)) : $unsigned($unsigned((8'hab)))) ?
                          (&$signed(reg3764)) : $signed((~|{reg3842})));
                    end
                  for (forvar3837 = (1'h0); (forvar3837 < (2'h2)); forvar3837 = (forvar3837 + (1'h1)))
                    begin
                      reg3838 <= (~$signed((reg3725 ? (|reg3793) : {(8'ha7)})));
                      reg3839 <= forvar3853[(4'hc):(4'h8)];
                      reg3840 <= (reg3762 | {(+(reg3739 > (8'hba)))});
                      reg3841 <= (~|reg3785);
                    end
                  reg3842 <= reg3799;
                end
            end
          for (forvar3856 = (1'h0); (forvar3856 < (1'h0)); forvar3856 = (forvar3856 + (1'h1)))
            begin
              reg3857 <= (8'h9d);
              for (forvar3858 = (1'h0); (forvar3858 < (1'h1)); forvar3858 = (forvar3858 + (1'h1)))
                begin
                  if (($unsigned($signed({reg3762})) ?
                      $signed(((reg3842 | (8'ha8)) - (reg3747 ?
                          reg3792 : reg3837))) : $unsigned(reg3775)))
                    begin
                      reg3859 <= $unsigned($unsigned(({(8'h9f)} == $unsigned(reg3771))));
                    end
                  else
                    begin
                      reg3859 <= reg3771[(2'h2):(1'h1)];
                      reg3860 <= (reg3775[(4'ha):(1'h0)] ?
                          (((reg3761 ? reg3726 : reg3798) ?
                                  (reg3754 ?
                                      reg3780 : reg3716) : $unsigned((8'hb9))) ?
                              (reg3847 > (~&reg3834)) : (+(reg3854 ?
                                  (8'ha4) : reg3759))) : $signed($unsigned(reg3759[(3'h5):(2'h3)])));
                      reg3861 <= reg3719;
                      reg3862 <= reg3846[(1'h1):(1'h1)];
                    end
                  for (forvar3863 = (1'h0); (forvar3863 < (1'h0)); forvar3863 = (forvar3863 + (1'h1)))
                    begin
                      reg3864 <= $signed(reg3740[(3'h5):(2'h2)]);
                      reg3865 <= ($signed($unsigned((^~reg3837))) ?
                          (|($unsigned(reg3842) + (^reg3739))) : $signed(reg3864[(4'h8):(4'h8)]));
                      reg3866 <= $unsigned(forvar3830[(1'h0):(1'h0)]);
                    end
                end
              for (forvar3867 = (1'h0); (forvar3867 < (2'h2)); forvar3867 = (forvar3867 + (1'h1)))
                begin
                  if (((reg3808[(1'h0):(1'h0)] ?
                          ((forvar3830 != reg3848) & reg3839) : (~|reg3865[(1'h1):(1'h1)])) ?
                      $unsigned((^~reg3778[(4'h9):(3'h7)])) : $unsigned($signed(forvar3836[(2'h2):(1'h1)]))))
                    begin
                      reg3868 <= reg3804;
                      reg3869 <= $signed(reg3726[(3'h5):(2'h3)]);
                      reg3870 <= $unsigned(reg3766);
                    end
                  else
                    begin
                      reg3868 <= {$unsigned(reg3784[(4'hd):(4'ha)])};
                      reg3869 <= $unsigned(forvar3858[(4'h9):(1'h0)]);
                    end
                end
            end
          reg3871 <= (!reg3738[(4'hc):(4'h8)]);
        end
      else
        begin
          if (reg3716)
            begin
              for (forvar3830 = (1'h0); (forvar3830 < (1'h0)); forvar3830 = (forvar3830 + (1'h1)))
                begin
                  for (forvar3831 = (1'h0); (forvar3831 < (2'h2)); forvar3831 = (forvar3831 + (1'h1)))
                    begin
                      reg3832 <= reg3812;
                      reg3833 <= $unsigned((8'h9e));
                      reg3834 <= forvar3856[(4'ha):(1'h1)];
                      reg3835 <= reg3838;
                    end
                  if (reg3751)
                    begin
                      reg3836 <= ((forvar3837[(2'h2):(1'h0)] - $unsigned($signed(reg3855))) + (~&({(8'hb2)} - $signed(reg3756))));
                      reg3837 <= $unsigned((!$unsigned(forvar3836[(2'h3):(2'h3)])));
                      reg3838 <= (|(reg3759 != reg3785));
                      reg3839 <= reg3848;
                    end
                  else
                    begin
                      reg3836 <= ($signed((reg3788 ^ (!reg3794))) | reg3788);
                      reg3837 <= (^reg3731);
                    end
                  reg3840 <= reg3784[(4'hc):(3'h4)];
                  for (forvar3841 = (1'h0); (forvar3841 < (1'h0)); forvar3841 = (forvar3841 + (1'h1)))
                    begin
                      reg3842 <= $unsigned($signed((reg3781 | {wire3828})));
                      reg3843 <= ($unsigned($signed(((8'hb6) >>> reg3866))) ?
                          (!forvar3845) : reg3736);
                    end
                end
              if (reg3837)
                begin
                  if (forvar3831[(3'h7):(3'h7)])
                    begin
                      reg3844 <= $unsigned({(~$unsigned(reg3734))});
                    end
                  else
                    begin
                      reg3844 <= {$signed((((8'ha8) ^ reg3853) ?
                              {wire3417} : $unsigned((8'ha0))))};
                    end
                  reg3845 <= ((~&$unsigned((reg3722 | reg3725))) - reg3777[(4'ha):(3'h5)]);
                  for (forvar3846 = (1'h0); (forvar3846 < (2'h3)); forvar3846 = (forvar3846 + (1'h1)))
                    begin
                      reg3847 <= ($signed(reg3755) != reg3820[(2'h2):(2'h2)]);
                      reg3848 <= reg3724[(4'h8):(3'h6)];
                      reg3849 <= reg3762;
                      reg3850 <= $unsigned(forvar3851);
                    end
                end
              else
                begin
                  reg3844 <= reg3807[(5'h10):(2'h2)];
                  reg3845 <= {$signed((8'hab))};
                  if ((reg3737 ?
                      ($unsigned($signed(reg3817)) - $signed((^reg3848))) : (~&{(reg3826 ?
                              reg3745 : reg3784)})))
                    begin
                      reg3846 <= reg3793[(1'h1):(1'h0)];
                      reg3847 <= $signed($signed(reg3835));
                      reg3848 <= (~&(8'hb2));
                    end
                  else
                    begin
                      reg3846 <= $signed(wire3418);
                      reg3847 <= $unsigned(({{reg3868}} * reg3740));
                    end
                  for (forvar3849 = (1'h0); (forvar3849 < (1'h1)); forvar3849 = (forvar3849 + (1'h1)))
                    begin
                      reg3850 <= reg3716[(1'h1):(1'h0)];
                      reg3851 <= (((forvar3863[(1'h0):(1'h0)] ~^ (reg3800 ?
                              reg3847 : (8'hba))) <= forvar3849[(2'h2):(2'h2)]) ?
                          {reg3836} : (($unsigned((8'h9e)) && reg3731[(1'h1):(1'h0)]) <<< $signed(((8'hae) - reg3751))));
                      reg3852 <= $signed((forvar3849[(2'h3):(1'h0)] ?
                          $unsigned((reg3784 ?
                              reg3818 : reg3800)) : $unsigned({reg3729})));
                    end
                end
            end
          else
            begin
              if ((reg3804 ^~ (8'h9d)))
                begin
                  for (forvar3830 = (1'h0); (forvar3830 < (2'h2)); forvar3830 = (forvar3830 + (1'h1)))
                    begin
                      reg3831 <= (~(((reg3811 >>> (8'hb5)) ?
                              reg3795 : (reg3734 * reg3737)) ?
                          ((reg3833 <<< reg3787) ?
                              $unsigned((8'hb3)) : {forvar3831}) : reg3784));
                      reg3832 <= (~&reg3859[(3'h4):(1'h1)]);
                      reg3833 <= (+reg3827[(2'h3):(1'h1)]);
                    end
                  for (forvar3834 = (1'h0); (forvar3834 < (2'h3)); forvar3834 = (forvar3834 + (1'h1)))
                    begin
                      reg3835 <= reg3731;
                      reg3836 <= (8'hb8);
                      reg3837 <= ({({reg3723} >= reg3824[(3'h7):(1'h0)])} < (reg3839[(2'h3):(2'h3)] ?
                          (reg3837 ? (-reg3731) : reg3738) : {(reg3815 ?
                                  reg3741 : reg3771)}));
                      reg3838 <= (8'h9f);
                    end
                  if (reg3773[(1'h0):(1'h0)])
                    begin
                      reg3839 <= {((((8'hb7) ~^ (8'had)) ?
                                  wire3420[(4'hd):(3'h5)] : reg3728[(4'hc):(4'hb)]) ?
                              forvar3831[(4'h9):(4'h9)] : ($unsigned(reg3846) ^~ (reg3791 != reg3847)))};
                    end
                  else
                    begin
                      reg3839 <= (!($unsigned($unsigned(reg3718)) ?
                          ($signed(reg3756) ?
                              $signed((8'ha3)) : (reg3781 ?
                                  forvar3841 : reg3756)) : reg3736));
                      reg3840 <= reg3803[(3'h4):(2'h3)];
                    end
                  if ((&reg3736))
                    begin
                      reg3841 <= (reg3745 + reg3844);
                      reg3842 <= (reg3844[(4'hd):(2'h3)] ?
                          (|$unsigned(reg3812)) : reg3836[(2'h2):(1'h0)]);
                      reg3843 <= $unsigned((+$unsigned((forvar3851 ?
                          (8'hb3) : reg3841))));
                    end
                  else
                    begin
                      reg3841 <= (($unsigned((reg3847 | reg3764)) ?
                          reg3861 : reg3740) - reg3742[(3'h4):(2'h2)]);
                      reg3842 <= (reg3850 - (reg3803[(4'h8):(1'h1)] ?
                          $unsigned(reg3831) : ($signed((8'ha5)) ?
                              (^(8'ha1)) : $unsigned(reg3862))));
                      reg3843 <= reg3840;
                    end
                end
              else
                begin
                  if ($signed(((~|(reg3843 != reg3812)) ?
                      reg3868 : (~^reg3860[(2'h3):(2'h2)]))))
                    begin
                      reg3830 <= $unsigned((~|(((8'ha8) ?
                          reg3781 : forvar3836) && $signed((8'hba)))));
                      reg3831 <= (~&reg3771);
                      reg3832 <= (&$unsigned(reg3836));
                    end
                  else
                    begin
                      reg3830 <= (reg3742[(2'h3):(1'h1)] ?
                          reg3814 : forvar3851[(4'h8):(3'h7)]);
                      reg3831 <= reg3761[(3'h5):(2'h2)];
                    end
                  if ($unsigned(reg3806))
                    begin
                      reg3833 <= (|$signed($unsigned((8'ha2))));
                      reg3834 <= (+(~&(+(reg3784 << reg3722))));
                      reg3835 <= reg3781;
                    end
                  else
                    begin
                      reg3833 <= (~reg3865[(2'h3):(1'h0)]);
                      reg3834 <= {{(reg3775[(4'he):(2'h3)] & $unsigned(forvar3832))}};
                    end
                  for (forvar3836 = (1'h0); (forvar3836 < (1'h1)); forvar3836 = (forvar3836 + (1'h1)))
                    begin
                      reg3837 <= reg3812[(1'h0):(1'h0)];
                      reg3838 <= ((reg3809 ~^ ($signed(reg3853) == (reg3869 | reg3795))) * (($unsigned(reg3838) < (reg3775 ?
                              reg3727 : reg3733)) ?
                          forvar3867 : $unsigned($signed(reg3727))));
                      reg3839 <= reg3758[(3'h4):(2'h3)];
                    end
                  if ($signed((~reg3820)))
                    begin
                      reg3840 <= {($signed(((8'h9c) <<< reg3783)) || forvar3858)};
                      reg3841 <= $signed(((reg3745[(2'h3):(2'h2)] ?
                          $unsigned(reg3758) : reg3826[(1'h0):(1'h0)]) >> (~|(reg3821 ?
                          (8'hba) : reg3733))));
                      reg3842 <= ($unsigned($unsigned({wire3418})) ?
                          (-(8'h9c)) : ((!{reg3834}) ?
                              {forvar3849} : (&reg3838[(3'h5):(1'h0)])));
                    end
                  else
                    begin
                      reg3840 <= wire3419[(4'ha):(4'ha)];
                      reg3841 <= reg3759;
                      reg3842 <= $unsigned((&reg3846[(2'h2):(1'h1)]));
                    end
                end
              reg3844 <= ({$unsigned(reg3755)} <<< $signed(((-reg3766) << reg3738[(3'h4):(2'h3)])));
              if (reg3742[(1'h1):(1'h0)])
                begin
                  if (($signed(reg3757) ?
                      {(|((8'ha8) << reg3804))} : $unsigned({reg3717[(4'h8):(3'h4)]})))
                    begin
                      reg3845 <= ((|reg3798) * ($unsigned(reg3795[(1'h0):(1'h0)]) ?
                          $unsigned((|reg3781)) : $signed(reg3739)));
                    end
                  else
                    begin
                      reg3845 <= (reg3716 ?
                          $unsigned(({reg3852} == (reg3745 <= forvar3856))) : reg3741[(4'ha):(3'h7)]);
                      reg3846 <= (reg3741[(3'h6):(1'h1)] & (-$unsigned((8'hb8))));
                      reg3847 <= $unsigned(reg3857[(3'h4):(3'h4)]);
                    end
                end
              else
                begin
                  for (forvar3845 = (1'h0); (forvar3845 < (1'h0)); forvar3845 = (forvar3845 + (1'h1)))
                    begin
                      reg3846 <= reg3848;
                      reg3847 <= (reg3789 > reg3802[(3'h4):(1'h0)]);
                    end
                  for (forvar3848 = (1'h0); (forvar3848 < (1'h0)); forvar3848 = (forvar3848 + (1'h1)))
                    begin
                      reg3849 <= (($unsigned((reg3803 > reg3777)) << (!(reg3794 ?
                              reg3822 : reg3729))) ?
                          (-(~|wire3420[(4'h9):(1'h1)])) : $unsigned(({reg3762} <<< (^reg3719))));
                      reg3850 <= ($unsigned(((reg3822 + reg3848) ?
                          $unsigned(reg3800) : (~|(8'hb7)))) == {((|forvar3845) ?
                              (reg3724 ~^ (8'ha6)) : reg3812)});
                    end
                end
              for (forvar3851 = (1'h0); (forvar3851 < (2'h2)); forvar3851 = (forvar3851 + (1'h1)))
                begin
                  reg3852 <= $unsigned($signed(reg3728[(4'hc):(2'h3)]));
                  for (forvar3853 = (1'h0); (forvar3853 < (2'h2)); forvar3853 = (forvar3853 + (1'h1)))
                    begin
                      reg3854 <= reg3728;
                      reg3855 <= reg3811;
                      reg3856 <= {(reg3717[(3'h7):(3'h7)] + reg3864[(2'h3):(2'h3)])};
                      reg3857 <= (~($unsigned((forvar3832 ?
                          (8'hb7) : forvar3841)) * ((8'hb9) == (reg3785 ?
                          reg3859 : reg3843))));
                    end
                  for (forvar3858 = (1'h0); (forvar3858 < (2'h3)); forvar3858 = (forvar3858 + (1'h1)))
                    begin
                      reg3859 <= (&reg3736[(3'h5):(2'h3)]);
                      reg3860 <= forvar3837;
                      reg3861 <= reg3739;
                      reg3862 <= {(($unsigned(reg3723) <= $unsigned(wire3828)) <= ((reg3817 ?
                              (8'hb5) : reg3780) <<< $unsigned(reg3719)))};
                    end
                end
            end
          if ((~&$signed(((reg3795 << forvar3863) ?
              $unsigned(reg3761) : (|reg3723)))))
            begin
              if (reg3719)
                begin
                  if ($signed($signed($unsigned($unsigned(reg3794)))))
                    begin
                      reg3863 <= reg3827;
                      reg3864 <= reg3856[(1'h1):(1'h0)];
                      reg3865 <= ((-$signed((!reg3740))) ?
                          wire3829[(2'h3):(2'h3)] : (^reg3802[(4'hc):(4'h9)]));
                    end
                  else
                    begin
                      reg3863 <= {reg3834[(4'h8):(3'h6)]};
                      reg3864 <= (wire3714 ? (+wire3714) : reg3844);
                      reg3865 <= {wire3828};
                    end
                end
              else
                begin
                  for (forvar3863 = (1'h0); (forvar3863 < (1'h1)); forvar3863 = (forvar3863 + (1'h1)))
                    begin
                      reg3864 <= $signed(reg3833[(3'h5):(2'h3)]);
                      reg3865 <= $signed(((~&(8'hb5)) < ($unsigned(reg3806) ^~ {(8'hb6)})));
                    end
                  for (forvar3866 = (1'h0); (forvar3866 < (1'h0)); forvar3866 = (forvar3866 + (1'h1)))
                    begin
                      reg3867 <= forvar3832;
                      reg3868 <= (reg3818 >> (((reg3831 <<< reg3794) ?
                              (&reg3799) : (reg3728 > reg3852)) ?
                          ($signed(reg3814) ~^ {reg3727}) : {(~|reg3868)}));
                    end
                  for (forvar3869 = (1'h0); (forvar3869 < (2'h2)); forvar3869 = (forvar3869 + (1'h1)))
                    begin
                      reg3870 <= $signed($signed(((+reg3807) ?
                          reg3800 : $unsigned((8'ha2)))));
                      reg3871 <= (reg3836 ~^ reg3824[(1'h0):(1'h0)]);
                    end
                end
              for (forvar3872 = (1'h0); (forvar3872 < (1'h1)); forvar3872 = (forvar3872 + (1'h1)))
                begin
                  if ({forvar3863})
                    begin
                      reg3873 <= (reg3773[(1'h1):(1'h1)] <<< forvar3849);
                      reg3874 <= reg3852;
                    end
                  else
                    begin
                      reg3873 <= (((~^(!reg3735)) ?
                          $unsigned((reg3865 ?
                              reg3836 : reg3822)) : (~reg3866)) | $unsigned(reg3764));
                      reg3874 <= $signed($signed((~^forvar3858)));
                      reg3875 <= $unsigned((^~{reg3752[(4'he):(3'h4)]}));
                    end
                  for (forvar3876 = (1'h0); (forvar3876 < (1'h1)); forvar3876 = (forvar3876 + (1'h1)))
                    begin
                      reg3877 <= (~&reg3787[(3'h4):(3'h4)]);
                    end
                end
            end
          else
            begin
              if ($unsigned(({reg3859} ~^ (~(~^reg3780)))))
                begin
                  for (forvar3863 = (1'h0); (forvar3863 < (1'h0)); forvar3863 = (forvar3863 + (1'h1)))
                    begin
                      reg3864 <= reg3844[(5'h10):(4'hd)];
                    end
                  for (forvar3865 = (1'h0); (forvar3865 < (2'h3)); forvar3865 = (forvar3865 + (1'h1)))
                    begin
                      reg3866 <= $signed((^~$unsigned((^~reg3842))));
                      reg3867 <= $signed(reg3857);
                      reg3868 <= forvar3830[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar3863 = (1'h0); (forvar3863 < (1'h0)); forvar3863 = (forvar3863 + (1'h1)))
                    begin
                      reg3864 <= $unsigned(reg3803);
                      reg3865 <= $unsigned((((reg3848 ?
                              reg3877 : forvar3869) <<< (!reg3834)) ?
                          (&(forvar3865 ? reg3777 : reg3748)) : {(~&reg3762)}));
                    end
                  for (forvar3866 = (1'h0); (forvar3866 < (1'h1)); forvar3866 = (forvar3866 + (1'h1)))
                    begin
                      reg3867 <= {(^~$unsigned($signed(reg3757)))};
                    end
                  if ((reg3853 ?
                      $unsigned(reg3817[(2'h2):(2'h2)]) : ($unsigned($signed((8'hb8))) ?
                          reg3749[(2'h3):(1'h1)] : $signed((^~reg3851)))))
                    begin
                      reg3868 <= $unsigned($signed(reg3774[(3'h4):(3'h4)]));
                    end
                  else
                    begin
                      reg3868 <= forvar3845;
                      reg3869 <= {(forvar3867[(4'he):(4'hc)] ?
                              {forvar3865[(1'h1):(1'h0)]} : reg3792[(3'h6):(2'h3)])};
                    end
                end
              for (forvar3870 = (1'h0); (forvar3870 < (1'h1)); forvar3870 = (forvar3870 + (1'h1)))
                begin
                  for (forvar3871 = (1'h0); (forvar3871 < (1'h1)); forvar3871 = (forvar3871 + (1'h1)))
                    begin
                      reg3872 <= reg3771;
                      reg3873 <= reg3832[(3'h4):(2'h2)];
                      reg3874 <= (8'hb1);
                    end
                end
              for (forvar3875 = (1'h0); (forvar3875 < (1'h0)); forvar3875 = (forvar3875 + (1'h1)))
                begin
                  for (forvar3876 = (1'h0); (forvar3876 < (2'h2)); forvar3876 = (forvar3876 + (1'h1)))
                    begin
                      reg3877 <= forvar3850[(4'h8):(3'h4)];
                      reg3878 <= {$unsigned(((~reg3735) ?
                              $unsigned(reg3823) : $signed(reg3824)))};
                    end
                  if ($signed(reg3849))
                    begin
                      reg3879 <= $unsigned($unsigned(forvar3867[(2'h2):(1'h1)]));
                      reg3880 <= $unsigned((+($unsigned(reg3771) ?
                          $unsigned(reg3859) : $signed(reg3830))));
                    end
                  else
                    begin
                      reg3879 <= ((((8'hb8) ^ (reg3771 <= reg3815)) ~^ {$unsigned((8'haa))}) ?
                          ($signed((&(8'hb3))) ?
                              forvar3832 : ((~reg3799) ?
                                  forvar3865[(1'h1):(1'h0)] : reg3841)) : $unsigned($unsigned($signed(reg3757))));
                      reg3880 <= wire3415[(2'h2):(2'h2)];
                      reg3881 <= reg3817;
                    end
                  for (forvar3882 = (1'h0); (forvar3882 < (2'h2)); forvar3882 = (forvar3882 + (1'h1)))
                    begin
                      reg3883 <= $signed(forvar3876[(1'h1):(1'h0)]);
                      reg3884 <= $unsigned($unsigned($signed({reg3806})));
                      reg3885 <= reg3788[(2'h2):(2'h2)];
                    end
                end
              for (forvar3886 = (1'h0); (forvar3886 < (2'h3)); forvar3886 = (forvar3886 + (1'h1)))
                begin
                  reg3887 <= ((|$signed($signed((8'h9d)))) ?
                      (&$signed($unsigned(reg3777))) : forvar3865);
                  for (forvar3888 = (1'h0); (forvar3888 < (2'h2)); forvar3888 = (forvar3888 + (1'h1)))
                    begin
                      reg3889 <= (forvar3850 ?
                          ((~^(^reg3769)) ?
                              reg3811[(4'ha):(4'ha)] : (reg3803[(2'h2):(2'h2)] ?
                                  $signed(forvar3832) : $unsigned(reg3840))) : (~&forvar3869[(2'h2):(1'h0)]));
                      reg3890 <= ((forvar3851 == $signed(reg3769)) < (reg3836 * ((~|reg3733) ?
                          (!(8'hb8)) : forvar3886[(5'h10):(2'h2)])));
                    end
                  reg3891 <= $unsigned(reg3723);
                  reg3892 <= reg3769;
                end
            end
          reg3893 <= {(|(^~$signed((8'ha8))))};
        end
    end
  assign wire3894 = reg3754[(3'h4):(1'h1)];
  assign wire3895 = $unsigned(((~|reg3815) ?
                        reg3787 : ($signed(reg3729) > reg3871[(4'ha):(4'ha)])));
  assign wire3896 = (~reg3742[(1'h0):(1'h0)]);
  assign wire3897 = (~^{$signed((&reg3861))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3421  (y, clk, wire3426, wire3425, wire3424, wire3423, wire3422);
  output wire [(32'hc65):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire3426;
  input wire signed [(4'hc):(1'h0)] wire3425;
  input wire signed [(4'hc):(1'h0)] wire3424;
  input wire signed [(4'h8):(1'h0)] wire3423;
  input wire signed [(2'h3):(1'h0)] wire3422;
  wire [(3'h4):(1'h0)] wire3713;
  wire signed [(3'h6):(1'h0)] wire3526;
  wire [(4'hc):(1'h0)] wire3525;
  wire signed [(4'he):(1'h0)] wire3524;
  wire signed [(3'h5):(1'h0)] wire3523;
  wire signed [(4'hd):(1'h0)] wire3522;
  reg signed [(2'h2):(1'h0)] reg3635 = (1'h0);
  reg [(2'h2):(1'h0)] reg3712 = (1'h0);
  reg [(3'h4):(1'h0)] reg3708 = (1'h0);
  reg [(3'h5):(1'h0)] reg3704 = (1'h0);
  reg [(4'hc):(1'h0)] reg3711 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3710 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3709 = (1'h0);
  reg [(4'hb):(1'h0)] reg3707 = (1'h0);
  reg [(4'hb):(1'h0)] reg3706 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3705 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3703 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3702 = (1'h0);
  reg [(4'hd):(1'h0)] reg3701 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3700 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3699 = (1'h0);
  reg [(3'h6):(1'h0)] reg3698 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3697 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3693 = (1'h0);
  reg [(4'ha):(1'h0)] reg3692 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3691 = (1'h0);
  reg [(5'h10):(1'h0)] reg3690 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3689 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3688 = (1'h0);
  reg [(4'hc):(1'h0)] reg3684 = (1'h0);
  reg [(4'hf):(1'h0)] reg3681 = (1'h0);
  reg [(4'hb):(1'h0)] reg3687 = (1'h0);
  reg [(4'hc):(1'h0)] reg3686 = (1'h0);
  reg [(4'h9):(1'h0)] reg3685 = (1'h0);
  reg [(4'hc):(1'h0)] reg3683 = (1'h0);
  reg [(4'hf):(1'h0)] reg3682 = (1'h0);
  reg [(5'h10):(1'h0)] reg3680 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3679 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3678 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3676 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3674 = (1'h0);
  reg [(4'hd):(1'h0)] reg3670 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3660 = (1'h0);
  reg [(4'ha):(1'h0)] reg3666 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3663 = (1'h0);
  reg [(3'h4):(1'h0)] reg3662 = (1'h0);
  reg [(3'h7):(1'h0)] reg3675 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3673 = (1'h0);
  reg [(2'h3):(1'h0)] reg3672 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3671 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3669 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3668 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3667 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3665 = (1'h0);
  reg [(4'hd):(1'h0)] reg3664 = (1'h0);
  reg [(5'h10):(1'h0)] reg3661 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3659 = (1'h0);
  reg [(2'h2):(1'h0)] reg3657 = (1'h0);
  reg [(4'h8):(1'h0)] reg3656 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3655 = (1'h0);
  reg [(4'hd):(1'h0)] reg3654 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3653 = (1'h0);
  reg [(2'h3):(1'h0)] reg3652 = (1'h0);
  reg [(4'hb):(1'h0)] reg3651 = (1'h0);
  reg [(4'h9):(1'h0)] reg3649 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3636 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3641 = (1'h0);
  reg [(3'h4):(1'h0)] reg3650 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3648 = (1'h0);
  reg [(2'h2):(1'h0)] reg3647 = (1'h0);
  reg [(5'h10):(1'h0)] reg3646 = (1'h0);
  reg [(4'hc):(1'h0)] reg3645 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3644 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3643 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3642 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3640 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3639 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3638 = (1'h0);
  reg [(5'h10):(1'h0)] reg3637 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3634 = (1'h0);
  reg [(3'h6):(1'h0)] reg3633 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3632 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3631 = (1'h0);
  reg [(4'h9):(1'h0)] reg3630 = (1'h0);
  reg [(4'hf):(1'h0)] reg3624 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3628 = (1'h0);
  reg [(4'hb):(1'h0)] reg3627 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3626 = (1'h0);
  reg [(4'he):(1'h0)] reg3625 = (1'h0);
  reg [(3'h6):(1'h0)] reg3623 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3619 = (1'h0);
  reg [(4'he):(1'h0)] reg3611 = (1'h0);
  reg [(4'h8):(1'h0)] reg3618 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3617 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3616 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3615 = (1'h0);
  reg [(4'hf):(1'h0)] reg3614 = (1'h0);
  reg [(5'h10):(1'h0)] reg3613 = (1'h0);
  reg [(4'he):(1'h0)] reg3612 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3610 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3609 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3608 = (1'h0);
  reg [(3'h7):(1'h0)] reg3605 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3604 = (1'h0);
  reg [(4'h9):(1'h0)] reg3583 = (1'h0);
  reg [(4'ha):(1'h0)] reg3574 = (1'h0);
  reg [(3'h5):(1'h0)] reg3571 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3553 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3529 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3528 = (1'h0);
  reg [(4'h9):(1'h0)] reg3599 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3603 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3602 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3601 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3600 = (1'h0);
  reg [(4'hb):(1'h0)] reg3598 = (1'h0);
  reg [(2'h2):(1'h0)] reg3597 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3595 = (1'h0);
  reg [(2'h3):(1'h0)] reg3594 = (1'h0);
  reg [(3'h5):(1'h0)] reg3592 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3591 = (1'h0);
  reg [(4'he):(1'h0)] reg3590 = (1'h0);
  reg [(4'he):(1'h0)] reg3589 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3587 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3586 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3585 = (1'h0);
  reg [(4'he):(1'h0)] reg3584 = (1'h0);
  reg [(3'h6):(1'h0)] reg3578 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3582 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3581 = (1'h0);
  reg [(5'h10):(1'h0)] reg3580 = (1'h0);
  reg [(4'hd):(1'h0)] reg3579 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3576 = (1'h0);
  reg [(4'h8):(1'h0)] reg3575 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3573 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3572 = (1'h0);
  reg [(4'hb):(1'h0)] reg3570 = (1'h0);
  reg [(4'he):(1'h0)] reg3569 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3566 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3561 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3568 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3567 = (1'h0);
  reg [(2'h2):(1'h0)] reg3565 = (1'h0);
  reg [(3'h7):(1'h0)] reg3564 = (1'h0);
  reg [(3'h7):(1'h0)] reg3563 = (1'h0);
  reg [(3'h4):(1'h0)] reg3562 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3559 = (1'h0);
  reg [(4'he):(1'h0)] reg3558 = (1'h0);
  reg [(3'h6):(1'h0)] reg3557 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3556 = (1'h0);
  reg [(4'ha):(1'h0)] reg3555 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3554 = (1'h0);
  reg [(2'h2):(1'h0)] reg3552 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3551 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3550 = (1'h0);
  reg [(3'h6):(1'h0)] reg3548 = (1'h0);
  reg [(2'h2):(1'h0)] reg3537 = (1'h0);
  reg [(3'h6):(1'h0)] reg3549 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3547 = (1'h0);
  reg [(2'h2):(1'h0)] reg3546 = (1'h0);
  reg [(3'h5):(1'h0)] reg3545 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3544 = (1'h0);
  reg [(3'h4):(1'h0)] reg3543 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3542 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3541 = (1'h0);
  reg [(2'h3):(1'h0)] reg3540 = (1'h0);
  reg [(3'h5):(1'h0)] reg3539 = (1'h0);
  reg [(2'h3):(1'h0)] reg3538 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3536 = (1'h0);
  reg [(2'h3):(1'h0)] reg3535 = (1'h0);
  reg [(4'hf):(1'h0)] reg3534 = (1'h0);
  reg [(4'hc):(1'h0)] reg3533 = (1'h0);
  reg [(3'h5):(1'h0)] reg3532 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3531 = (1'h0);
  reg [(4'hd):(1'h0)] reg3530 = (1'h0);
  reg [(4'hd):(1'h0)] reg3497 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3521 = (1'h0);
  reg [(4'he):(1'h0)] reg3520 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3519 = (1'h0);
  reg [(3'h7):(1'h0)] reg3518 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3517 = (1'h0);
  reg [(4'he):(1'h0)] reg3516 = (1'h0);
  reg [(3'h4):(1'h0)] reg3514 = (1'h0);
  reg [(4'he):(1'h0)] reg3513 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3512 = (1'h0);
  reg [(2'h3):(1'h0)] reg3511 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3510 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3509 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3508 = (1'h0);
  reg [(5'h10):(1'h0)] reg3507 = (1'h0);
  reg [(5'h10):(1'h0)] reg3506 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3504 = (1'h0);
  reg [(2'h2):(1'h0)] reg3503 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3501 = (1'h0);
  reg [(4'h9):(1'h0)] reg3500 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3499 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3498 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3427 = (1'h0);
  reg [(4'he):(1'h0)] reg3468 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3466 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3457 = (1'h0);
  reg [(4'hd):(1'h0)] reg3456 = (1'h0);
  reg [(3'h4):(1'h0)] reg3494 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3493 = (1'h0);
  reg [(3'h6):(1'h0)] reg3492 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3491 = (1'h0);
  reg [(3'h6):(1'h0)] reg3490 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3489 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3488 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3487 = (1'h0);
  reg [(3'h5):(1'h0)] reg3486 = (1'h0);
  reg [(3'h4):(1'h0)] reg3484 = (1'h0);
  reg [(4'hc):(1'h0)] reg3483 = (1'h0);
  reg [(3'h6):(1'h0)] reg3482 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3481 = (1'h0);
  reg [(3'h4):(1'h0)] reg3478 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3477 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3476 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3475 = (1'h0);
  reg [(5'h10):(1'h0)] reg3474 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3472 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3471 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3470 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3469 = (1'h0);
  reg [(4'hb):(1'h0)] reg3467 = (1'h0);
  reg [(2'h3):(1'h0)] reg3465 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3464 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3463 = (1'h0);
  reg [(4'he):(1'h0)] reg3462 = (1'h0);
  reg [(4'hd):(1'h0)] reg3461 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3460 = (1'h0);
  reg [(5'h10):(1'h0)] reg3459 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3458 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3455 = (1'h0);
  reg [(4'hb):(1'h0)] reg3445 = (1'h0);
  reg [(4'hd):(1'h0)] reg3454 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3453 = (1'h0);
  reg [(2'h2):(1'h0)] reg3452 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3451 = (1'h0);
  reg [(3'h7):(1'h0)] reg3450 = (1'h0);
  reg [(5'h10):(1'h0)] reg3449 = (1'h0);
  reg [(2'h2):(1'h0)] reg3448 = (1'h0);
  reg [(3'h6):(1'h0)] reg3447 = (1'h0);
  reg [(4'ha):(1'h0)] reg3446 = (1'h0);
  reg [(4'ha):(1'h0)] reg3436 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3434 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3444 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3443 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3442 = (1'h0);
  reg [(3'h4):(1'h0)] reg3441 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3440 = (1'h0);
  reg [(3'h6):(1'h0)] reg3439 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3438 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3437 = (1'h0);
  reg [(4'hf):(1'h0)] reg3435 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3433 = (1'h0);
  reg [(4'hb):(1'h0)] reg3432 = (1'h0);
  reg [(4'hc):(1'h0)] reg3431 = (1'h0);
  reg [(3'h4):(1'h0)] reg3430 = (1'h0);
  reg [(4'h9):(1'h0)] reg3429 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3428 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3708 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3704 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3696 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3695 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3694 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3685 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3684 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3681 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3677 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3672 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3671 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3668 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3665 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3674 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3670 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3666 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3663 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3662 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3660 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3658 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3650 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3642 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3638 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3645 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3649 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3641 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3636 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3635 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3629 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3624 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3622 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3621 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3620 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3611 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3607 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3606 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3604 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3585 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3581 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3568 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3544 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3555 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3545 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3540 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3536 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3599 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3596 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3593 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3588 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3583 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3578 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3577 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3574 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3571 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3567 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3566 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3561 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3560 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3553 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3551 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3549 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3541 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3548 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3537 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3529 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3528 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3527 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3515 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3505 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3502 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3497 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3496 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3495 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3460 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3459 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3455 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3448 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3447 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3444 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3441 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3433 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3465 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3462 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3485 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3480 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3479 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3473 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3468 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3466 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3457 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3456 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3442 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3445 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3437 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3436 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3434 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3427 = (1'h0);
  assign y = {wire3713,
                 wire3526,
                 wire3525,
                 wire3524,
                 wire3523,
                 wire3522,
                 reg3635,
                 reg3712,
                 reg3708,
                 reg3704,
                 reg3711,
                 reg3710,
                 reg3709,
                 reg3707,
                 reg3706,
                 reg3705,
                 reg3703,
                 reg3702,
                 reg3701,
                 reg3700,
                 reg3699,
                 reg3698,
                 reg3697,
                 reg3693,
                 reg3692,
                 reg3691,
                 reg3690,
                 reg3689,
                 reg3688,
                 reg3684,
                 reg3681,
                 reg3687,
                 reg3686,
                 reg3685,
                 reg3683,
                 reg3682,
                 reg3680,
                 reg3679,
                 reg3678,
                 reg3676,
                 reg3674,
                 reg3670,
                 reg3660,
                 reg3666,
                 reg3663,
                 reg3662,
                 reg3675,
                 reg3673,
                 reg3672,
                 reg3671,
                 reg3669,
                 reg3668,
                 reg3667,
                 reg3665,
                 reg3664,
                 reg3661,
                 reg3659,
                 reg3657,
                 reg3656,
                 reg3655,
                 reg3654,
                 reg3653,
                 reg3652,
                 reg3651,
                 reg3649,
                 reg3636,
                 reg3641,
                 reg3650,
                 reg3648,
                 reg3647,
                 reg3646,
                 reg3645,
                 reg3644,
                 reg3643,
                 reg3642,
                 reg3640,
                 reg3639,
                 reg3638,
                 reg3637,
                 reg3634,
                 reg3633,
                 reg3632,
                 reg3631,
                 reg3630,
                 reg3624,
                 reg3628,
                 reg3627,
                 reg3626,
                 reg3625,
                 reg3623,
                 reg3619,
                 reg3611,
                 reg3618,
                 reg3617,
                 reg3616,
                 reg3615,
                 reg3614,
                 reg3613,
                 reg3612,
                 reg3610,
                 reg3609,
                 reg3608,
                 reg3605,
                 reg3604,
                 reg3583,
                 reg3574,
                 reg3571,
                 reg3553,
                 reg3529,
                 reg3528,
                 reg3599,
                 reg3603,
                 reg3602,
                 reg3601,
                 reg3600,
                 reg3598,
                 reg3597,
                 reg3595,
                 reg3594,
                 reg3592,
                 reg3591,
                 reg3590,
                 reg3589,
                 reg3587,
                 reg3586,
                 reg3585,
                 reg3584,
                 reg3578,
                 reg3582,
                 reg3581,
                 reg3580,
                 reg3579,
                 reg3576,
                 reg3575,
                 reg3573,
                 reg3572,
                 reg3570,
                 reg3569,
                 reg3566,
                 reg3561,
                 reg3568,
                 reg3567,
                 reg3565,
                 reg3564,
                 reg3563,
                 reg3562,
                 reg3559,
                 reg3558,
                 reg3557,
                 reg3556,
                 reg3555,
                 reg3554,
                 reg3552,
                 reg3551,
                 reg3550,
                 reg3548,
                 reg3537,
                 reg3549,
                 reg3547,
                 reg3546,
                 reg3545,
                 reg3544,
                 reg3543,
                 reg3542,
                 reg3541,
                 reg3540,
                 reg3539,
                 reg3538,
                 reg3536,
                 reg3535,
                 reg3534,
                 reg3533,
                 reg3532,
                 reg3531,
                 reg3530,
                 reg3497,
                 reg3521,
                 reg3520,
                 reg3519,
                 reg3518,
                 reg3517,
                 reg3516,
                 reg3514,
                 reg3513,
                 reg3512,
                 reg3511,
                 reg3510,
                 reg3509,
                 reg3508,
                 reg3507,
                 reg3506,
                 reg3504,
                 reg3503,
                 reg3501,
                 reg3500,
                 reg3499,
                 reg3498,
                 reg3427,
                 reg3468,
                 reg3466,
                 reg3457,
                 reg3456,
                 reg3494,
                 reg3493,
                 reg3492,
                 reg3491,
                 reg3490,
                 reg3489,
                 reg3488,
                 reg3487,
                 reg3486,
                 reg3484,
                 reg3483,
                 reg3482,
                 reg3481,
                 reg3478,
                 reg3477,
                 reg3476,
                 reg3475,
                 reg3474,
                 reg3472,
                 reg3471,
                 reg3470,
                 reg3469,
                 reg3467,
                 reg3465,
                 reg3464,
                 reg3463,
                 reg3462,
                 reg3461,
                 reg3460,
                 reg3459,
                 reg3458,
                 reg3455,
                 reg3445,
                 reg3454,
                 reg3453,
                 reg3452,
                 reg3451,
                 reg3450,
                 reg3449,
                 reg3448,
                 reg3447,
                 reg3446,
                 reg3436,
                 reg3434,
                 reg3444,
                 reg3443,
                 reg3442,
                 reg3441,
                 reg3440,
                 reg3439,
                 reg3438,
                 reg3437,
                 reg3435,
                 reg3433,
                 reg3432,
                 reg3431,
                 reg3430,
                 reg3429,
                 reg3428,
                 forvar3708,
                 forvar3704,
                 forvar3696,
                 forvar3695,
                 forvar3694,
                 forvar3685,
                 forvar3684,
                 forvar3681,
                 forvar3677,
                 forvar3672,
                 forvar3671,
                 forvar3668,
                 forvar3665,
                 forvar3674,
                 forvar3670,
                 forvar3666,
                 forvar3663,
                 forvar3662,
                 forvar3660,
                 forvar3658,
                 forvar3650,
                 forvar3642,
                 forvar3638,
                 forvar3645,
                 forvar3649,
                 forvar3641,
                 forvar3636,
                 forvar3635,
                 forvar3629,
                 forvar3624,
                 forvar3622,
                 forvar3621,
                 forvar3620,
                 forvar3611,
                 forvar3607,
                 forvar3606,
                 forvar3604,
                 forvar3585,
                 forvar3581,
                 forvar3568,
                 forvar3544,
                 forvar3555,
                 forvar3545,
                 forvar3540,
                 forvar3536,
                 forvar3599,
                 forvar3596,
                 forvar3593,
                 forvar3588,
                 forvar3583,
                 forvar3578,
                 forvar3577,
                 forvar3574,
                 forvar3571,
                 forvar3567,
                 forvar3566,
                 forvar3561,
                 forvar3560,
                 forvar3553,
                 forvar3551,
                 forvar3549,
                 forvar3541,
                 forvar3548,
                 forvar3537,
                 forvar3529,
                 forvar3528,
                 forvar3527,
                 forvar3515,
                 forvar3505,
                 forvar3502,
                 forvar3497,
                 forvar3496,
                 forvar3495,
                 forvar3460,
                 forvar3459,
                 forvar3455,
                 forvar3448,
                 forvar3447,
                 forvar3444,
                 forvar3441,
                 forvar3433,
                 forvar3465,
                 forvar3462,
                 forvar3485,
                 forvar3480,
                 forvar3479,
                 forvar3473,
                 forvar3468,
                 forvar3466,
                 forvar3457,
                 forvar3456,
                 forvar3442,
                 forvar3445,
                 forvar3437,
                 forvar3436,
                 forvar3434,
                 forvar3427,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($signed({wire3424[(4'h8):(3'h5)]}))
        begin
          if ((((8'ha5) ?
              wire3426[(3'h7):(1'h0)] : {(wire3424 ?
                      (8'hab) : wire3423)}) + wire3423[(3'h4):(1'h0)]))
            begin
              for (forvar3427 = (1'h0); (forvar3427 < (1'h0)); forvar3427 = (forvar3427 + (1'h1)))
                begin
                  reg3428 <= $signed(wire3425[(2'h2):(1'h1)]);
                  reg3429 <= ((((wire3423 ?
                          (8'hb6) : wire3425) >= {forvar3427}) - ({wire3426} < (wire3425 ?
                          wire3423 : wire3424))) ?
                      (^~$unsigned((wire3424 > wire3426))) : (wire3422[(2'h3):(2'h3)] >= (wire3426 ?
                          $unsigned(wire3425) : (wire3426 ^ reg3428))));
                  if ((reg3428[(3'h5):(3'h5)] ? $unsigned(wire3426) : reg3429))
                    begin
                      reg3430 <= ((~^$unsigned($unsigned(wire3423))) ?
                          (((|forvar3427) >> $signed(wire3425)) ?
                              (wire3425[(4'hb):(4'h8)] + (8'ha6)) : $signed($unsigned(wire3426))) : (^wire3425[(3'h7):(1'h1)]));
                      reg3431 <= $unsigned(($unsigned($unsigned(wire3422)) ?
                          $signed({reg3429}) : (~$unsigned(reg3430))));
                      reg3432 <= (-$signed(({(8'hb3)} ?
                          $signed((8'haf)) : wire3424)));
                      reg3433 <= (-(!((wire3423 <= wire3422) ?
                          $unsigned(wire3424) : (reg3430 - wire3424))));
                    end
                  else
                    begin
                      reg3430 <= $unsigned($signed(($signed(wire3425) << wire3426)));
                      reg3431 <= (wire3426 ?
                          (({wire3423} & (&wire3425)) * ((wire3422 & wire3422) ?
                              $unsigned(wire3423) : (8'ha8))) : {wire3423[(3'h5):(3'h4)]});
                    end
                end
              for (forvar3434 = (1'h0); (forvar3434 < (1'h0)); forvar3434 = (forvar3434 + (1'h1)))
                begin
                  reg3435 <= ((-(&(wire3425 < forvar3427))) ?
                      (+wire3422) : ((reg3431 <= wire3424[(4'h9):(3'h7)]) ?
                          ((forvar3434 - (8'ha9)) ?
                              wire3423[(3'h4):(1'h0)] : $signed(reg3431)) : $unsigned((reg3431 ?
                              wire3425 : reg3429))));
                  for (forvar3436 = (1'h0); (forvar3436 < (1'h1)); forvar3436 = (forvar3436 + (1'h1)))
                    begin
                      reg3437 <= (+(-$unsigned((reg3435 ?
                          reg3433 : wire3426))));
                      reg3438 <= (&forvar3427[(1'h1):(1'h0)]);
                      reg3439 <= reg3430[(1'h0):(1'h0)];
                      reg3440 <= (forvar3427[(1'h0):(1'h0)] ?
                          $signed(reg3438[(1'h1):(1'h0)]) : (~|reg3438[(1'h1):(1'h1)]));
                    end
                  if (reg3428[(3'h5):(3'h4)])
                    begin
                      reg3441 <= $unsigned($unsigned(({(8'hb4)} ?
                          $unsigned((8'hb2)) : $unsigned(reg3440))));
                      reg3442 <= $unsigned($unsigned($signed(reg3433)));
                      reg3443 <= {forvar3436};
                    end
                  else
                    begin
                      reg3441 <= reg3433[(3'h6):(2'h3)];
                      reg3442 <= reg3433[(4'h8):(2'h3)];
                      reg3443 <= forvar3427[(1'h0):(1'h0)];
                    end
                  if ((~^((reg3438 ?
                      (8'hb4) : (reg3441 < reg3443)) ^~ wire3422)))
                    begin
                      reg3444 <= $unsigned(wire3422[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg3444 <= (reg3442[(4'hc):(1'h0)] ^~ ((reg3441 >> $unsigned(reg3439)) ^~ reg3444));
                    end
                end
            end
          else
            begin
              for (forvar3427 = (1'h0); (forvar3427 < (1'h0)); forvar3427 = (forvar3427 + (1'h1)))
                begin
                  if (wire3424[(1'h1):(1'h0)])
                    begin
                      reg3428 <= wire3423[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg3428 <= ((reg3439 ?
                          (((8'ha8) > reg3435) || $signed(reg3430)) : reg3429) + $signed($unsigned($signed(reg3437))));
                      reg3429 <= (8'hb2);
                      reg3430 <= reg3443[(3'h7):(2'h3)];
                      reg3431 <= {$unsigned((forvar3434 >>> $unsigned(reg3428)))};
                    end
                  reg3432 <= forvar3436[(1'h0):(1'h0)];
                end
              if ($signed($signed($signed((reg3444 ? wire3424 : wire3425)))))
                begin
                  if ({(reg3428[(1'h0):(1'h0)] < ($unsigned(reg3439) ?
                          (8'h9f) : (wire3423 ? (8'h9d) : wire3426)))})
                    begin
                      reg3433 <= $signed(reg3431);
                      reg3434 <= $signed(reg3437);
                    end
                  else
                    begin
                      reg3433 <= ({reg3438[(1'h0):(1'h0)]} ?
                          reg3440[(4'hc):(2'h3)] : ((^~(~^reg3443)) ?
                              ((~&(8'hb8)) ?
                                  forvar3427[(1'h0):(1'h0)] : (forvar3434 ?
                                      forvar3434 : reg3443)) : forvar3436[(3'h7):(1'h0)]));
                      reg3434 <= $unsigned((~$signed($signed(reg3432))));
                      reg3435 <= $unsigned(($signed({reg3441}) ?
                          (forvar3427 ?
                              (reg3442 ?
                                  reg3434 : reg3444) : (wire3422 << reg3439)) : (reg3435[(4'he):(1'h0)] ?
                              $signed(forvar3427) : $unsigned(reg3433))));
                      reg3436 <= {$unsigned({(wire3423 ? wire3426 : reg3432)})};
                    end
                  for (forvar3437 = (1'h0); (forvar3437 < (2'h3)); forvar3437 = (forvar3437 + (1'h1)))
                    begin
                      reg3438 <= (!wire3426);
                      reg3439 <= wire3423[(2'h2):(2'h2)];
                    end
                end
              else
                begin
                  if ({$signed(((wire3422 >= (8'h9e)) && (reg3440 < forvar3436)))})
                    begin
                      reg3433 <= (|$unsigned($unsigned({reg3441})));
                      reg3434 <= {(-wire3424)};
                    end
                  else
                    begin
                      reg3433 <= (wire3424[(3'h7):(2'h3)] ?
                          forvar3427[(2'h2):(2'h2)] : forvar3427);
                      reg3434 <= (($signed((reg3443 ?
                              (8'ha6) : reg3437)) != (|reg3441[(1'h1):(1'h1)])) ?
                          (~^((forvar3427 * reg3433) ?
                              {forvar3427} : (wire3425 & wire3423))) : (8'ha8));
                      reg3435 <= reg3429[(3'h6):(1'h0)];
                    end
                  for (forvar3436 = (1'h0); (forvar3436 < (2'h2)); forvar3436 = (forvar3436 + (1'h1)))
                    begin
                      reg3437 <= $unsigned(($unsigned((~&wire3422)) ^ reg3440[(3'h5):(3'h4)]));
                      reg3438 <= $signed(reg3433);
                      reg3439 <= ($unsigned((|$signed((8'hb3)))) > (~&(^reg3431)));
                      reg3440 <= reg3438;
                    end
                  reg3441 <= $unsigned($signed((forvar3434 ?
                      $signed(reg3429) : (8'haa))));
                end
              if ({$unsigned($unsigned((+reg3430)))})
                begin
                  if ((wire3426[(3'h4):(3'h4)] > reg3429))
                    begin
                      reg3442 <= ((reg3441 < $signed((&reg3433))) * ($unsigned(reg3431) <<< reg3439[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg3442 <= ((|(reg3437[(2'h2):(1'h1)] != (~^wire3425))) ?
                          $signed(((8'hb0) - (forvar3436 < (8'hb4)))) : (reg3433 >>> reg3430));
                      reg3443 <= (^(((reg3432 ?
                              reg3433 : wire3425) >= ((8'haf) > reg3441)) ?
                          (&reg3443[(1'h1):(1'h1)]) : (~&(reg3444 < reg3439))));
                      reg3444 <= (~reg3444);
                    end
                  for (forvar3445 = (1'h0); (forvar3445 < (2'h3)); forvar3445 = (forvar3445 + (1'h1)))
                    begin
                      reg3446 <= {$unsigned(((reg3428 ? reg3441 : forvar3434) ?
                              reg3435 : reg3437[(2'h3):(1'h1)]))};
                      reg3447 <= $signed(reg3439);
                      reg3448 <= wire3426[(2'h3):(2'h3)];
                    end
                  if (reg3433)
                    begin
                      reg3449 <= ($unsigned($unsigned((8'hb0))) ?
                          (|$signed($signed(forvar3445))) : forvar3436[(3'h4):(2'h2)]);
                      reg3450 <= ($signed(reg3447) ?
                          forvar3445 : $signed((~$signed(wire3423))));
                    end
                  else
                    begin
                      reg3449 <= $unsigned(($signed((~&wire3422)) & reg3428));
                      reg3450 <= reg3438[(1'h1):(1'h1)];
                    end
                  if ($signed($unsigned(((reg3448 - wire3425) ?
                      forvar3436[(3'h6):(2'h3)] : ((8'ha0) ~^ reg3444)))))
                    begin
                      reg3451 <= ($unsigned({(reg3435 ?
                              reg3439 : reg3449)}) * $unsigned(((~(8'hb5)) ?
                          (reg3441 < reg3448) : wire3422[(1'h0):(1'h0)])));
                      reg3452 <= (^$signed(wire3426[(3'h4):(3'h4)]));
                      reg3453 <= {reg3438[(1'h1):(1'h1)]};
                      reg3454 <= reg3447[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3451 <= (8'hac);
                      reg3452 <= wire3426;
                      reg3453 <= reg3440[(4'hb):(3'h4)];
                    end
                end
              else
                begin
                  for (forvar3442 = (1'h0); (forvar3442 < (2'h3)); forvar3442 = (forvar3442 + (1'h1)))
                    begin
                      reg3443 <= reg3454;
                    end
                  if ((^~forvar3436))
                    begin
                      reg3444 <= (~(((reg3435 * reg3449) << $unsigned(wire3422)) ?
                          reg3441 : (-$signed(forvar3445))));
                      reg3445 <= (^(((wire3424 & reg3444) <<< wire3423[(2'h3):(2'h3)]) & reg3442[(3'h6):(3'h6)]));
                    end
                  else
                    begin
                      reg3444 <= (reg3449 ~^ (reg3432 ?
                          ($signed(reg3445) > {reg3440}) : reg3437));
                      reg3445 <= $signed((((reg3436 ?
                          (8'hb0) : reg3446) <<< forvar3442[(2'h2):(2'h2)]) || ((~&reg3444) ?
                          (reg3442 ? reg3454 : forvar3445) : (-reg3443))));
                    end
                  reg3446 <= $unsigned((({reg3445} >> $signed(forvar3434)) ^ $unsigned($unsigned(reg3439))));
                  reg3447 <= ($signed(((reg3430 ? reg3444 : reg3451) ?
                          (-wire3422) : (wire3425 && (8'hae)))) ?
                      reg3430 : reg3430);
                end
              reg3455 <= forvar3445;
            end
          if (reg3440[(4'h8):(2'h2)])
            begin
              for (forvar3456 = (1'h0); (forvar3456 < (2'h2)); forvar3456 = (forvar3456 + (1'h1)))
                begin
                  for (forvar3457 = (1'h0); (forvar3457 < (1'h0)); forvar3457 = (forvar3457 + (1'h1)))
                    begin
                      reg3458 <= forvar3427;
                      reg3459 <= reg3454[(3'h6):(3'h6)];
                      reg3460 <= $unsigned(reg3443);
                      reg3461 <= $unsigned((8'haa));
                    end
                  if ((~&(!(8'h9e))))
                    begin
                      reg3462 <= ({reg3431[(4'ha):(3'h5)]} ?
                          (8'h9c) : ($unsigned((~|reg3435)) | ((reg3442 <= forvar3442) ?
                              (reg3455 && forvar3445) : (8'ha9))));
                      reg3463 <= reg3448[(2'h2):(1'h0)];
                      reg3464 <= ($unsigned((~|$signed(reg3436))) == $signed((forvar3434 ?
                          $signed(reg3460) : $unsigned(reg3434))));
                      reg3465 <= (^~($unsigned((reg3429 * (8'ha0))) << reg3449[(4'hc):(4'hc)]));
                    end
                  else
                    begin
                      reg3462 <= ($signed(($unsigned(reg3446) < (wire3426 ^~ forvar3456))) != (((forvar3457 ?
                                  reg3436 : reg3436) ?
                              $unsigned(forvar3427) : $unsigned(forvar3437)) ?
                          reg3442 : ({reg3439} ?
                              (^~forvar3457) : reg3455[(1'h1):(1'h0)])));
                      reg3463 <= reg3439[(3'h5):(3'h4)];
                      reg3464 <= ({wire3425[(3'h7):(1'h1)]} - $unsigned({$signed(reg3444)}));
                    end
                end
              for (forvar3466 = (1'h0); (forvar3466 < (2'h3)); forvar3466 = (forvar3466 + (1'h1)))
                begin
                  reg3467 <= reg3463;
                  for (forvar3468 = (1'h0); (forvar3468 < (2'h2)); forvar3468 = (forvar3468 + (1'h1)))
                    begin
                      reg3469 <= (+$unsigned($signed(reg3462[(4'h8):(1'h1)])));
                      reg3470 <= $signed($signed(reg3465[(2'h3):(1'h0)]));
                      reg3471 <= (({(wire3425 * (8'ha9))} >= ($unsigned(reg3443) != (forvar3434 ?
                              wire3422 : reg3455))) ?
                          $signed(reg3463[(2'h2):(1'h0)]) : $unsigned($signed($unsigned(reg3461))));
                      reg3472 <= forvar3468[(1'h1):(1'h0)];
                    end
                  for (forvar3473 = (1'h0); (forvar3473 < (2'h2)); forvar3473 = (forvar3473 + (1'h1)))
                    begin
                      reg3474 <= reg3462[(4'ha):(3'h6)];
                      reg3475 <= $signed($unsigned(wire3424[(3'h5):(1'h1)]));
                      reg3476 <= (^~((8'ha8) ? reg3438 : {(^~reg3469)}));
                      reg3477 <= $unsigned($unsigned(reg3450[(3'h7):(2'h2)]));
                    end
                end
              reg3478 <= ($signed($unsigned((!forvar3457))) ?
                  (($signed(reg3436) ?
                      (forvar3457 ? reg3474 : (8'h9e)) : (reg3455 ?
                          reg3446 : reg3435)) ^ (~^((8'ha5) ~^ reg3443))) : reg3459);
              for (forvar3479 = (1'h0); (forvar3479 < (1'h1)); forvar3479 = (forvar3479 + (1'h1)))
                begin
                  for (forvar3480 = (1'h0); (forvar3480 < (2'h2)); forvar3480 = (forvar3480 + (1'h1)))
                    begin
                      reg3481 <= (~(reg3463 <= forvar3437));
                      reg3482 <= reg3465[(2'h3):(1'h1)];
                      reg3483 <= (({reg3450[(2'h3):(1'h1)]} ?
                          ((~forvar3456) || $unsigned(reg3459)) : (~|wire3425)) ^~ $signed(reg3432[(3'h7):(3'h4)]));
                      reg3484 <= $signed(reg3469[(4'ha):(3'h5)]);
                    end
                  for (forvar3485 = (1'h0); (forvar3485 < (1'h1)); forvar3485 = (forvar3485 + (1'h1)))
                    begin
                      reg3486 <= reg3431;
                    end
                  if ($unsigned((!reg3474[(4'ha):(3'h4)])))
                    begin
                      reg3487 <= $signed($unsigned(({reg3448} | (forvar3468 ?
                          (8'hb9) : forvar3473))));
                      reg3488 <= (reg3464 ?
                          {(~(reg3487 ~^ reg3471))} : $unsigned(reg3459));
                    end
                  else
                    begin
                      reg3487 <= $unsigned(({$signed(reg3438)} <= $unsigned($signed(forvar3437))));
                      reg3488 <= $signed((+((!wire3424) ?
                          $unsigned((8'ha6)) : reg3477)));
                      reg3489 <= $signed(($unsigned(reg3483[(3'h6):(2'h2)]) & (8'ha4)));
                      reg3490 <= reg3447;
                    end
                  if ({$unsigned(((forvar3445 ?
                          forvar3434 : reg3431) << {reg3444}))})
                    begin
                      reg3491 <= ((&$unsigned($unsigned(reg3477))) ?
                          $signed((reg3437 ?
                              reg3437 : $signed((8'had)))) : reg3450);
                      reg3492 <= $signed($unsigned(({reg3488} ~^ $signed(reg3460))));
                      reg3493 <= $signed(($unsigned($signed(reg3481)) >> (8'h9e)));
                    end
                  else
                    begin
                      reg3491 <= ($signed($signed((&reg3428))) ?
                          (((~&reg3490) ^~ (|reg3438)) + (!reg3445)) : $unsigned(((reg3447 ?
                                  reg3474 : reg3459) ?
                              (reg3477 <<< reg3438) : {reg3451})));
                      reg3492 <= (forvar3442[(1'h1):(1'h0)] ?
                          reg3487[(4'hc):(2'h2)] : $unsigned((((8'h9f) ?
                                  forvar3427 : forvar3434) ?
                              $signed(reg3442) : (reg3440 ?
                                  forvar3442 : reg3439))));
                      reg3493 <= $unsigned(({(!reg3475)} ?
                          (8'had) : {reg3478[(1'h1):(1'h0)]}));
                      reg3494 <= {$unsigned(({reg3448} ^ (8'had)))};
                    end
                end
            end
          else
            begin
              if (((((8'ha3) ?
                      $signed(reg3494) : (forvar3468 ? reg3449 : reg3447)) ?
                  (~$unsigned(forvar3434)) : (-(reg3465 > (8'ha5)))) < reg3488))
                begin
                  if (wire3422)
                    begin
                      reg3456 <= $unsigned((&forvar3437[(1'h0):(1'h0)]));
                      reg3457 <= reg3433;
                    end
                  else
                    begin
                      reg3456 <= $unsigned(reg3438);
                      reg3457 <= reg3484;
                    end
                  if ((forvar3442 == wire3424))
                    begin
                      reg3458 <= (^~{(reg3469 ?
                              reg3450[(1'h0):(1'h0)] : $unsigned(reg3444))});
                      reg3459 <= reg3428[(3'h4):(2'h3)];
                      reg3460 <= reg3489;
                      reg3461 <= $signed(($unsigned({reg3475}) > ((forvar3442 << reg3431) ?
                          (reg3436 ? forvar3436 : reg3432) : (reg3437 ?
                              reg3447 : forvar3434))));
                    end
                  else
                    begin
                      reg3458 <= $unsigned($signed(($unsigned(reg3432) ^~ wire3425)));
                    end
                  for (forvar3462 = (1'h0); (forvar3462 < (2'h3)); forvar3462 = (forvar3462 + (1'h1)))
                    begin
                      reg3463 <= (^{reg3454[(3'h7):(3'h4)]});
                      reg3464 <= $signed((-forvar3462));
                    end
                  for (forvar3465 = (1'h0); (forvar3465 < (2'h3)); forvar3465 = (forvar3465 + (1'h1)))
                    begin
                      reg3466 <= ($unsigned((reg3477[(2'h2):(2'h2)] ?
                          {reg3489} : {reg3447})) << ((!((8'hb8) * reg3451)) ^ forvar3479));
                      reg3467 <= reg3446[(1'h0):(1'h0)];
                      reg3468 <= $signed($signed($unsigned(reg3440[(3'h4):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar3456 = (1'h0); (forvar3456 < (1'h0)); forvar3456 = (forvar3456 + (1'h1)))
                    begin
                      reg3457 <= (^~(~&reg3465));
                      reg3458 <= ({(~(reg3494 ?
                              forvar3457 : reg3494))} * reg3457[(2'h2):(1'h0)]);
                    end
                end
            end
        end
      else
        begin
          if ((!$signed(reg3455)))
            begin
              for (forvar3427 = (1'h0); (forvar3427 < (2'h2)); forvar3427 = (forvar3427 + (1'h1)))
                begin
                  reg3428 <= (!(8'hba));
                  if ((|$signed(reg3474[(4'h9):(1'h1)])))
                    begin
                      reg3429 <= reg3445;
                    end
                  else
                    begin
                      reg3429 <= reg3478[(2'h3):(1'h0)];
                      reg3430 <= $signed(reg3458);
                      reg3431 <= reg3462[(3'h7):(3'h6)];
                      reg3432 <= ($unsigned(((8'h9d) ?
                          (&forvar3466) : (^(8'ha3)))) | (8'hb6));
                    end
                  for (forvar3433 = (1'h0); (forvar3433 < (1'h0)); forvar3433 = (forvar3433 + (1'h1)))
                    begin
                      reg3434 <= ((($unsigned(reg3475) ?
                          wire3423 : (~(8'hb6))) ^~ {reg3481}) <<< $unsigned($unsigned(forvar3456[(3'h6):(2'h3)])));
                      reg3435 <= $signed((~^reg3493[(4'h9):(1'h0)]));
                      reg3436 <= reg3441;
                    end
                  if (forvar3437[(1'h0):(1'h0)])
                    begin
                      reg3437 <= (~^$unsigned((8'ha3)));
                      reg3438 <= $unsigned($signed((forvar3457 & (8'hb1))));
                      reg3439 <= $signed((^~$unsigned(reg3447[(2'h3):(1'h0)])));
                      reg3440 <= {(8'ha4)};
                    end
                  else
                    begin
                      reg3437 <= reg3483[(2'h3):(2'h2)];
                      reg3438 <= forvar3427;
                      reg3439 <= (^(|forvar3473[(1'h1):(1'h0)]));
                    end
                end
              if (reg3461)
                begin
                  for (forvar3441 = (1'h0); (forvar3441 < (1'h1)); forvar3441 = (forvar3441 + (1'h1)))
                    begin
                      reg3442 <= (!($unsigned(reg3464[(3'h4):(3'h4)]) ?
                          ((|(8'hb3)) <= (forvar3445 ?
                              reg3470 : reg3456)) : $signed(reg3455)));
                    end
                  reg3443 <= (+$unsigned(($unsigned((8'ha7)) <= ((8'ha0) > (8'ha4)))));
                  for (forvar3444 = (1'h0); (forvar3444 < (1'h1)); forvar3444 = (forvar3444 + (1'h1)))
                    begin
                      reg3445 <= {forvar3465[(3'h4):(2'h2)]};
                    end
                end
              else
                begin
                  if ((8'hae))
                    begin
                      reg3441 <= reg3466;
                      reg3442 <= $unsigned((reg3449 ?
                          ((+reg3452) ?
                              reg3484[(2'h3):(1'h0)] : $unsigned(forvar3427)) : (~|(forvar3465 < forvar3462))));
                    end
                  else
                    begin
                      reg3441 <= (forvar3445[(3'h6):(2'h3)] < forvar3433);
                      reg3442 <= $unsigned((reg3455 ?
                          reg3463[(1'h0):(1'h0)] : ((reg3477 ?
                                  reg3451 : (8'haa)) ?
                              (reg3475 ? (8'h9d) : reg3470) : reg3447)));
                      reg3443 <= {reg3442};
                      reg3444 <= (^~($signed((~^reg3478)) >> reg3445));
                    end
                end
            end
          else
            begin
              if ((|reg3432))
                begin
                  for (forvar3427 = (1'h0); (forvar3427 < (2'h2)); forvar3427 = (forvar3427 + (1'h1)))
                    begin
                      reg3428 <= forvar3457[(4'h8):(2'h3)];
                      reg3429 <= reg3460;
                      reg3430 <= reg3493[(3'h5):(1'h0)];
                    end
                  if ($unsigned($unsigned($unsigned($signed(forvar3437)))))
                    begin
                      reg3431 <= forvar3442[(1'h0):(1'h0)];
                      reg3432 <= (+($signed(forvar3457) ?
                          reg3445 : (!{reg3490})));
                      reg3433 <= {(+(reg3433[(3'h4):(2'h2)] ?
                              reg3446[(4'h9):(3'h6)] : $signed(forvar3433)))};
                      reg3434 <= wire3426;
                    end
                  else
                    begin
                      reg3431 <= reg3442;
                    end
                  if ((reg3477 > ({((8'ha7) >= (8'haf))} * $unsigned(reg3438))))
                    begin
                      reg3435 <= (!(((reg3449 < reg3468) ?
                              wire3425[(4'h8):(2'h2)] : (forvar3479 & forvar3485)) ?
                          (forvar3457[(3'h5):(2'h3)] == (reg3481 ?
                              reg3433 : forvar3462)) : $unsigned($signed(reg3462))));
                      reg3436 <= (^$unsigned(forvar3434));
                    end
                  else
                    begin
                      reg3435 <= (~&(($unsigned(reg3482) ?
                              (reg3437 != (8'ha3)) : (reg3494 ?
                                  reg3459 : forvar3466)) ?
                          (wire3422[(2'h3):(2'h2)] ?
                              $unsigned((8'ha4)) : $signed(wire3424)) : $unsigned((~forvar3434))));
                    end
                  for (forvar3437 = (1'h0); (forvar3437 < (2'h3)); forvar3437 = (forvar3437 + (1'h1)))
                    begin
                      reg3438 <= $unsigned($signed({$signed(reg3453)}));
                      reg3439 <= reg3435;
                      reg3440 <= {forvar3437[(3'h4):(2'h2)]};
                      reg3441 <= ((((~^wire3425) ?
                              $unsigned(wire3426) : $signed(reg3435)) || {(-(8'h9e))}) ?
                          $signed(reg3444) : reg3468);
                    end
                end
              else
                begin
                  if ($signed((reg3467[(2'h2):(1'h1)] * (~(forvar3457 ?
                      reg3487 : reg3491)))))
                    begin
                      reg3427 <= $unsigned($signed({forvar3444[(1'h0):(1'h0)]}));
                      reg3428 <= (!($signed((+reg3484)) >> (reg3438 ?
                          (~reg3489) : (|(8'ha1)))));
                      reg3429 <= $unsigned((~^(((8'hab) | reg3457) << ((8'ha1) && reg3456))));
                    end
                  else
                    begin
                      reg3427 <= $signed({(~|(reg3467 ? reg3472 : reg3467))});
                    end
                  if ((~&$unsigned((^(reg3427 <<< reg3491)))))
                    begin
                      reg3430 <= (reg3461 <<< (^$unsigned((&forvar3456))));
                      reg3431 <= reg3452;
                      reg3432 <= ($unsigned((reg3481 < $unsigned(reg3429))) ?
                          {((reg3478 ? reg3464 : reg3444) ?
                                  $signed(reg3464) : reg3494)} : $signed($unsigned((reg3466 != reg3466))));
                      reg3433 <= $signed((&$signed(forvar3457)));
                    end
                  else
                    begin
                      reg3430 <= $unsigned($signed(((8'h9e) ?
                          (8'hb8) : $unsigned(reg3478))));
                      reg3431 <= {reg3455[(3'h5):(2'h3)]};
                    end
                  for (forvar3434 = (1'h0); (forvar3434 < (1'h0)); forvar3434 = (forvar3434 + (1'h1)))
                    begin
                      reg3435 <= $unsigned($unsigned(reg3448));
                      reg3436 <= $signed($unsigned($signed(reg3455[(2'h2):(1'h1)])));
                    end
                  for (forvar3437 = (1'h0); (forvar3437 < (1'h0)); forvar3437 = (forvar3437 + (1'h1)))
                    begin
                      reg3438 <= $unsigned(($unsigned($signed(reg3484)) ?
                          $signed((-wire3426)) : ((forvar3466 <<< forvar3436) ~^ reg3466)));
                      reg3439 <= (~|forvar3436);
                      reg3440 <= reg3481;
                      reg3441 <= (((~$unsigned(reg3492)) ?
                              forvar3427 : (~|$unsigned(forvar3441))) ?
                          $signed(reg3452) : wire3426[(3'h6):(2'h3)]);
                    end
                end
            end
          reg3446 <= {($signed(reg3469[(4'ha):(1'h0)]) & reg3458[(3'h5):(1'h1)])};
          if ({(~|({forvar3434} << {forvar3456}))})
            begin
              if (reg3475)
                begin
                  reg3447 <= $signed(({(-forvar3462)} | forvar3433[(4'h8):(3'h6)]));
                end
              else
                begin
                  for (forvar3447 = (1'h0); (forvar3447 < (1'h0)); forvar3447 = (forvar3447 + (1'h1)))
                    begin
                      reg3448 <= ($signed($unsigned({forvar3444})) ?
                          forvar3445 : (~$unsigned((reg3446 ?
                              forvar3462 : reg3489))));
                      reg3449 <= $signed($signed($unsigned((reg3444 ?
                          wire3423 : reg3489))));
                      reg3450 <= reg3465;
                      reg3451 <= (~&reg3447[(2'h2):(1'h1)]);
                    end
                end
            end
          else
            begin
              for (forvar3447 = (1'h0); (forvar3447 < (2'h3)); forvar3447 = (forvar3447 + (1'h1)))
                begin
                  for (forvar3448 = (1'h0); (forvar3448 < (2'h2)); forvar3448 = (forvar3448 + (1'h1)))
                    begin
                      reg3449 <= $signed((($signed(forvar3444) ?
                          forvar3479 : reg3439) * $unsigned($signed(wire3423))));
                    end
                  if ((|($signed((forvar3444 ? reg3467 : reg3455)) ?
                      reg3447[(3'h4):(3'h4)] : $unsigned((reg3477 + reg3450)))))
                    begin
                      reg3450 <= forvar3468;
                      reg3451 <= reg3427[(3'h4):(1'h0)];
                      reg3452 <= reg3457[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg3450 <= (~^reg3470);
                      reg3451 <= forvar3447[(4'h8):(3'h4)];
                      reg3452 <= (~^(~|$signed((~reg3443))));
                      reg3453 <= reg3462;
                    end
                  reg3454 <= ({$unsigned(reg3477)} >> $unsigned(($signed(reg3456) ?
                      $signed(wire3425) : wire3426)));
                  for (forvar3455 = (1'h0); (forvar3455 < (2'h3)); forvar3455 = (forvar3455 + (1'h1)))
                    begin
                      reg3456 <= (((!(reg3493 ?
                          reg3460 : forvar3465)) || (reg3463 < forvar3480[(1'h0):(1'h0)])) | (8'hb9));
                      reg3457 <= ($signed(reg3431[(2'h2):(1'h0)]) ?
                          ($signed({reg3430}) ?
                              $unsigned(forvar3445[(3'h5):(2'h2)]) : (reg3448[(2'h2):(1'h1)] ^~ ((8'h9c) - (8'h9e)))) : (!reg3446[(1'h1):(1'h1)]));
                    end
                end
              reg3458 <= $unsigned((-{(reg3442 ? reg3430 : (8'hb0))}));
              for (forvar3459 = (1'h0); (forvar3459 < (1'h1)); forvar3459 = (forvar3459 + (1'h1)))
                begin
                  for (forvar3460 = (1'h0); (forvar3460 < (2'h2)); forvar3460 = (forvar3460 + (1'h1)))
                    begin
                      reg3461 <= forvar3437;
                      reg3462 <= $unsigned((~|(((8'had) + forvar3485) ?
                          $unsigned((8'ha7)) : $signed(reg3436))));
                      reg3463 <= {{$unsigned($signed(reg3457))}};
                      reg3464 <= ($unsigned($unsigned((reg3442 < (8'ha7)))) > {{{reg3470}}});
                    end
                end
              reg3465 <= reg3483;
            end
        end
      if ((($unsigned((reg3448 ? reg3482 : reg3488)) - $signed(reg3471)) ?
          reg3461[(4'ha):(2'h2)] : $signed(($signed(forvar3436) > $signed(forvar3448)))))
        begin
          for (forvar3495 = (1'h0); (forvar3495 < (1'h0)); forvar3495 = (forvar3495 + (1'h1)))
            begin
              for (forvar3496 = (1'h0); (forvar3496 < (2'h3)); forvar3496 = (forvar3496 + (1'h1)))
                begin
                  for (forvar3497 = (1'h0); (forvar3497 < (2'h3)); forvar3497 = (forvar3497 + (1'h1)))
                    begin
                      reg3498 <= $unsigned({{(8'hb9)}});
                    end
                  if ($signed((forvar3436 ^ ($unsigned(reg3442) << reg3476))))
                    begin
                      reg3499 <= ((~|({forvar3442} < (reg3433 != forvar3445))) ?
                          (reg3460[(1'h1):(1'h1)] << ((reg3451 > reg3448) << (~&reg3494))) : $signed($unsigned((reg3454 ?
                              reg3490 : reg3453))));
                      reg3500 <= forvar3455;
                      reg3501 <= reg3443[(4'ha):(4'ha)];
                    end
                  else
                    begin
                      reg3499 <= $unsigned(($signed($unsigned(reg3481)) ?
                          reg3482 : forvar3445));
                      reg3500 <= reg3443[(1'h0):(1'h0)];
                      reg3501 <= (^(((forvar3456 || reg3467) >= $signed(reg3462)) ?
                          $signed(reg3448) : (~^$signed(forvar3462))));
                    end
                  for (forvar3502 = (1'h0); (forvar3502 < (2'h3)); forvar3502 = (forvar3502 + (1'h1)))
                    begin
                      reg3503 <= ((-($signed((8'h9d)) ?
                          $signed(reg3468) : reg3491[(2'h2):(2'h2)])) - (~^{(|reg3487)}));
                      reg3504 <= wire3423;
                    end
                  for (forvar3505 = (1'h0); (forvar3505 < (2'h2)); forvar3505 = (forvar3505 + (1'h1)))
                    begin
                      reg3506 <= $signed({$unsigned($unsigned(reg3471))});
                      reg3507 <= (({forvar3505[(2'h3):(1'h1)]} ?
                          ($unsigned(forvar3456) == $signed(reg3460)) : reg3490[(2'h3):(2'h2)]) != (reg3451[(1'h1):(1'h0)] + $unsigned(reg3477[(1'h0):(1'h0)])));
                      reg3508 <= (($unsigned(reg3484) ?
                          {reg3459[(1'h0):(1'h0)]} : $unsigned(reg3476[(2'h2):(1'h0)])) << ($signed((reg3437 | reg3466)) ?
                          reg3467 : (8'hb4)));
                      reg3509 <= $unsigned(reg3489[(2'h3):(1'h0)]);
                    end
                end
              reg3510 <= $signed(((&(reg3446 & forvar3465)) - $signed($signed(wire3424))));
              if (reg3449)
                begin
                  if ((~(^reg3437)))
                    begin
                      reg3511 <= reg3442[(4'hc):(3'h5)];
                    end
                  else
                    begin
                      reg3511 <= (~&$unsigned($signed({reg3475})));
                      reg3512 <= (+($unsigned((reg3478 ?
                          wire3426 : reg3474)) | $signed(reg3468)));
                      reg3513 <= {({(&reg3452)} ?
                              $unsigned(reg3449[(3'h7):(3'h7)]) : forvar3456)};
                    end
                end
              else
                begin
                  if (wire3423)
                    begin
                      reg3511 <= {$signed((~^$signed(reg3471)))};
                      reg3512 <= $unsigned({({(8'hab)} ?
                              (reg3452 ?
                                  reg3498 : reg3469) : $signed((8'hb1)))});
                      reg3513 <= $unsigned(reg3486[(3'h5):(3'h4)]);
                      reg3514 <= reg3490[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg3511 <= forvar3465[(4'h9):(3'h4)];
                      reg3512 <= ({(reg3433[(1'h0):(1'h0)] ?
                              (reg3500 ?
                                  forvar3457 : reg3452) : (^reg3454))} < ((+(forvar3447 ?
                              reg3432 : forvar3434)) ?
                          reg3449 : (reg3449[(4'hb):(3'h5)] ?
                              $signed((8'hb6)) : ((8'hb2) ?
                                  reg3490 : reg3432))));
                      reg3513 <= {(~&($signed(reg3461) >>> $signed(reg3444)))};
                      reg3514 <= $unsigned((-$unsigned((^~(8'ha3)))));
                    end
                end
              for (forvar3515 = (1'h0); (forvar3515 < (1'h1)); forvar3515 = (forvar3515 + (1'h1)))
                begin
                  reg3516 <= $signed($unsigned($unsigned((-forvar3437))));
                  if (reg3472[(3'h4):(1'h0)])
                    begin
                      reg3517 <= ($signed($unsigned(reg3457[(4'hb):(3'h4)])) >= (&reg3441[(1'h1):(1'h1)]));
                      reg3518 <= {reg3472[(1'h1):(1'h1)]};
                      reg3519 <= forvar3460;
                    end
                  else
                    begin
                      reg3517 <= (forvar3465[(2'h2):(1'h0)] ?
                          reg3467[(2'h2):(1'h1)] : (|(~|(~&forvar3448))));
                      reg3518 <= {$unsigned(reg3430[(2'h2):(2'h2)])};
                    end
                  reg3520 <= wire3426[(3'h5):(2'h3)];
                  reg3521 <= $signed((reg3499 == reg3481[(2'h2):(1'h1)]));
                end
            end
        end
      else
        begin
          for (forvar3495 = (1'h0); (forvar3495 < (2'h3)); forvar3495 = (forvar3495 + (1'h1)))
            begin
              for (forvar3496 = (1'h0); (forvar3496 < (1'h1)); forvar3496 = (forvar3496 + (1'h1)))
                begin
                  if ($unsigned({reg3519[(1'h1):(1'h0)]}))
                    begin
                      reg3497 <= reg3492[(2'h2):(2'h2)];
                      reg3498 <= (reg3508 >= (~|reg3483[(2'h3):(2'h2)]));
                      reg3499 <= (forvar3427 ?
                          $unsigned(reg3441[(2'h3):(2'h2)]) : reg3440);
                    end
                  else
                    begin
                      reg3497 <= $unsigned(reg3429);
                      reg3498 <= reg3468[(4'he):(4'hd)];
                      reg3499 <= (~&forvar3502);
                    end
                end
            end
        end
    end
  assign wire3522 = (8'ha6);
  assign wire3523 = reg3450[(3'h7):(2'h2)];
  assign wire3524 = ($signed((reg3428 ? (~|reg3464) : (^reg3451))) ?
                        reg3440 : {((^~reg3478) ~^ (~wire3422))});
  assign wire3525 = reg3477[(2'h2):(1'h0)];
  assign wire3526 = (^$signed(reg3521));
  always
    @(posedge clk) begin
      if (((((reg3478 ? (8'hb4) : reg3492) ?
                  (reg3469 ? reg3478 : reg3484) : (reg3516 ?
                      reg3474 : reg3433)) ?
              ($signed(reg3456) ?
                  reg3449 : $signed(wire3526)) : {$unsigned(reg3442)}) ?
          $signed(((reg3451 ? reg3471 : wire3525) ?
              $signed((8'hb9)) : (|reg3445))) : (-reg3428[(2'h3):(2'h3)])))
        begin
          for (forvar3527 = (1'h0); (forvar3527 < (1'h0)); forvar3527 = (forvar3527 + (1'h1)))
            begin
              for (forvar3528 = (1'h0); (forvar3528 < (2'h2)); forvar3528 = (forvar3528 + (1'h1)))
                begin
                  for (forvar3529 = (1'h0); (forvar3529 < (2'h2)); forvar3529 = (forvar3529 + (1'h1)))
                    begin
                      reg3530 <= ($unsigned((reg3454[(2'h2):(1'h1)] ?
                          $unsigned(wire3523) : {reg3481})) >> (8'hba));
                      reg3531 <= $unsigned((~&({reg3509} * reg3461[(3'h5):(2'h2)])));
                      reg3532 <= ({($unsigned(reg3450) ?
                              (8'hb7) : (reg3491 == reg3465))} | reg3467);
                      reg3533 <= reg3448;
                    end
                  reg3534 <= (({((8'ha0) ? reg3518 : reg3471)} ?
                      ((~^reg3448) ?
                          (wire3525 ~^ wire3526) : reg3508[(3'h5):(2'h3)]) : $unsigned(reg3481)) == $unsigned(($signed(reg3451) ?
                      reg3475 : reg3483)));
                  reg3535 <= reg3499[(1'h0):(1'h0)];
                  reg3536 <= reg3475;
                end
            end
          if ($signed((&{(|reg3472)})))
            begin
              if ((reg3489[(2'h2):(2'h2)] ?
                  $unsigned((reg3509[(1'h0):(1'h0)] ?
                      (~&reg3429) : reg3429[(4'h9):(2'h2)])) : reg3463))
                begin
                  for (forvar3537 = (1'h0); (forvar3537 < (2'h3)); forvar3537 = (forvar3537 + (1'h1)))
                    begin
                      reg3538 <= reg3486[(1'h1):(1'h1)];
                      reg3539 <= (-$unsigned((^(-(8'hb8)))));
                      reg3540 <= reg3501;
                      reg3541 <= $signed((~|((reg3509 >> reg3513) != (-reg3430))));
                    end
                end
              else
                begin
                  for (forvar3537 = (1'h0); (forvar3537 < (2'h3)); forvar3537 = (forvar3537 + (1'h1)))
                    begin
                      reg3538 <= $signed($signed(reg3446));
                      reg3539 <= reg3514;
                      reg3540 <= reg3440[(4'hc):(3'h4)];
                      reg3541 <= (&(^~(!(^(8'hb6)))));
                    end
                  if (reg3472)
                    begin
                      reg3542 <= ($signed((reg3489 <= (reg3504 * reg3491))) <= reg3510[(2'h3):(1'h1)]);
                      reg3543 <= (^{(reg3452 ^~ (~reg3475))});
                      reg3544 <= $unsigned({($signed((8'ha1)) <= {wire3525})});
                    end
                  else
                    begin
                      reg3542 <= $unsigned(($unsigned($unsigned(reg3538)) ?
                          ($signed(reg3513) >= {reg3530}) : (^~(reg3504 == reg3437))));
                      reg3543 <= reg3433[(2'h3):(1'h0)];
                      reg3544 <= reg3520;
                      reg3545 <= $signed($unsigned(reg3475[(4'h9):(4'h8)]));
                    end
                  if (reg3470)
                    begin
                      reg3546 <= {$unsigned((+{reg3440}))};
                      reg3547 <= ((^(reg3428 < reg3467)) << {wire3525});
                    end
                  else
                    begin
                      reg3546 <= {$unsigned(reg3504)};
                      reg3547 <= ((~^$unsigned($unsigned(reg3510))) >>> ($unsigned((&forvar3528)) ?
                          reg3491[(3'h4):(2'h3)] : ($signed(reg3456) >= (8'hb1))));
                    end
                  for (forvar3548 = (1'h0); (forvar3548 < (1'h0)); forvar3548 = (forvar3548 + (1'h1)))
                    begin
                      reg3549 <= (({reg3544} ?
                          (((8'ha6) ^ reg3457) ^~ (8'hb7)) : ($signed(reg3478) * (reg3490 > forvar3527))) <= reg3497);
                    end
                end
            end
          else
            begin
              if ($unsigned($unsigned({(reg3546 ? reg3443 : reg3428)})))
                begin
                  if (reg3498)
                    begin
                      reg3537 <= ((^$unsigned($signed((8'hb4)))) ?
                          forvar3548 : (8'hb9));
                      reg3538 <= ((((reg3481 ? reg3499 : reg3481) ?
                                  reg3539 : reg3465[(1'h0):(1'h0)]) ?
                              ((wire3422 ?
                                  reg3510 : reg3506) >>> $unsigned(reg3434)) : (8'ha4)) ?
                          ($signed(reg3482[(1'h1):(1'h0)]) << $signed((wire3522 | (8'ha5)))) : {reg3443});
                      reg3539 <= reg3443;
                      reg3540 <= reg3498;
                    end
                  else
                    begin
                      reg3537 <= ((~({reg3456} ?
                          (reg3466 ?
                              reg3456 : reg3437) : $signed(reg3431))) + (~|reg3492[(3'h6):(2'h2)]));
                      reg3538 <= $signed((reg3535[(1'h1):(1'h0)] ?
                          {(reg3465 ?
                                  reg3433 : (8'h9d))} : (~|((8'ha9) > wire3423))));
                    end
                  if ({(reg3444[(2'h2):(1'h0)] ?
                          $signed((reg3474 | reg3518)) : ((wire3425 ?
                                  reg3546 : (8'h9f)) ?
                              (+reg3461) : ((8'had) ? reg3467 : reg3462)))})
                    begin
                      reg3541 <= $signed(wire3523[(2'h3):(1'h0)]);
                      reg3542 <= $signed($signed(reg3459[(3'h7):(2'h3)]));
                      reg3543 <= $unsigned((((reg3494 && reg3492) ?
                          reg3507[(1'h1):(1'h0)] : $signed(reg3547)) && (~|$signed(reg3547))));
                    end
                  else
                    begin
                      reg3541 <= reg3489[(2'h3):(2'h2)];
                    end
                  reg3544 <= ($signed(({reg3470} ^~ $unsigned(reg3535))) >> ((reg3434[(1'h0):(1'h0)] << {reg3538}) ?
                      (-forvar3527) : ((&(8'ha6)) ~^ ((8'ha5) >= reg3477))));
                  reg3545 <= reg3504[(1'h1):(1'h0)];
                end
              else
                begin
                  if (reg3494[(1'h0):(1'h0)])
                    begin
                      reg3537 <= (+$unsigned(reg3509));
                      reg3538 <= $signed({reg3508});
                      reg3539 <= $signed(($unsigned({reg3488}) ?
                          ((8'haa) ?
                              (8'ha1) : $signed(reg3436)) : ($signed((8'hba)) || (reg3455 ?
                              reg3471 : reg3464))));
                      reg3540 <= reg3544;
                    end
                  else
                    begin
                      reg3537 <= ($unsigned($unsigned((reg3454 + (8'ha8)))) ?
                          reg3543 : $unsigned(((~^(8'ha4)) ?
                              $signed(reg3486) : (reg3510 ?
                                  (8'ha4) : (8'haf)))));
                      reg3538 <= reg3471;
                    end
                  for (forvar3541 = (1'h0); (forvar3541 < (2'h2)); forvar3541 = (forvar3541 + (1'h1)))
                    begin
                      reg3542 <= $signed(wire3423);
                      reg3543 <= ((+($unsigned(reg3500) && $unsigned(reg3492))) ?
                          reg3444 : reg3451[(1'h1):(1'h1)]);
                      reg3544 <= (($signed((8'hb1)) ?
                          reg3506 : $signed($signed(reg3538))) >= ($signed(reg3518[(3'h6):(2'h3)]) && ({reg3539} ~^ $signed(reg3472))));
                    end
                  if (($unsigned(forvar3548) ?
                      $unsigned((((8'hba) ? reg3533 : forvar3528) ?
                          reg3431 : reg3475)) : reg3500[(2'h3):(1'h1)]))
                    begin
                      reg3545 <= {(reg3506[(4'hf):(4'hd)] ?
                              (reg3444 << $signed(reg3544)) : $unsigned(reg3438))};
                    end
                  else
                    begin
                      reg3545 <= reg3518;
                      reg3546 <= ($unsigned((~(reg3482 ^~ reg3469))) ?
                          ((8'ha8) && reg3481) : (wire3425 + (wire3423[(3'h7):(3'h5)] ?
                              reg3468 : $unsigned((8'hb1)))));
                      reg3547 <= $signed(reg3546[(1'h1):(1'h1)]);
                      reg3548 <= ((|$signed((8'h9e))) - (reg3530[(3'h5):(1'h1)] ?
                          (reg3466[(2'h3):(2'h2)] ?
                              $unsigned(reg3447) : $signed(wire3424)) : $signed($signed(wire3424))));
                    end
                end
              if (($signed($unsigned(reg3439[(3'h4):(1'h1)])) ?
                  (&(((8'hb6) | (8'ha9)) && wire3524[(4'hb):(3'h7)])) : ((8'hb6) || reg3519[(2'h2):(1'h1)])))
                begin
                  for (forvar3549 = (1'h0); (forvar3549 < (2'h3)); forvar3549 = (forvar3549 + (1'h1)))
                    begin
                      reg3550 <= {((~$unsigned(reg3460)) ?
                              ($unsigned((8'hb7)) ^~ reg3474[(4'hf):(4'h8)]) : (~^reg3489))};
                    end
                  if ((-($signed((reg3441 ^~ reg3537)) + {(8'hab)})))
                    begin
                      reg3551 <= ((((+(8'haa)) ?
                          (~&reg3436) : (wire3425 - reg3489)) || ($signed(forvar3548) ?
                          $unsigned(wire3526) : reg3469[(3'h7):(1'h0)])) & reg3547);
                    end
                  else
                    begin
                      reg3551 <= {reg3543};
                    end
                end
              else
                begin
                  for (forvar3549 = (1'h0); (forvar3549 < (2'h2)); forvar3549 = (forvar3549 + (1'h1)))
                    begin
                      reg3550 <= $unsigned($signed((reg3492[(2'h3):(2'h3)] ?
                          $signed((8'ha2)) : reg3449)));
                    end
                  for (forvar3551 = (1'h0); (forvar3551 < (2'h2)); forvar3551 = (forvar3551 + (1'h1)))
                    begin
                      reg3552 <= ((+forvar3551[(2'h2):(1'h0)]) >>> {{(reg3483 ?
                                  reg3474 : reg3542)}});
                    end
                  for (forvar3553 = (1'h0); (forvar3553 < (1'h0)); forvar3553 = (forvar3553 + (1'h1)))
                    begin
                      reg3554 <= (|({(reg3450 ? reg3476 : (8'hb3))} ?
                          $unsigned(reg3477) : reg3471));
                      reg3555 <= $signed($signed(reg3453[(3'h6):(3'h4)]));
                    end
                  if ($unsigned((reg3512 ?
                      reg3520[(4'h8):(3'h4)] : $signed((~reg3554)))))
                    begin
                      reg3556 <= ($unsigned(((reg3543 ? (8'ha3) : (8'haf)) ?
                              (reg3532 ?
                                  reg3500 : reg3459) : $unsigned(reg3546))) ?
                          $signed({(~&reg3436)}) : reg3476[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg3556 <= (((^wire3526[(1'h1):(1'h0)]) >>> (((8'hba) ?
                              (8'h9e) : reg3537) ?
                          reg3547 : $unsigned(reg3475))) >>> (&($unsigned((8'had)) ?
                          reg3488 : reg3519[(2'h2):(2'h2)])));
                      reg3557 <= ((~|reg3543) ?
                          $unsigned((reg3517[(2'h3):(2'h3)] ?
                              $unsigned(reg3436) : reg3538)) : reg3442[(4'he):(4'hb)]);
                      reg3558 <= reg3507;
                      reg3559 <= $signed($unsigned(($signed(reg3497) + reg3488[(1'h0):(1'h0)])));
                    end
                end
            end
          for (forvar3560 = (1'h0); (forvar3560 < (2'h2)); forvar3560 = (forvar3560 + (1'h1)))
            begin
              if (reg3509[(2'h3):(2'h2)])
                begin
                  for (forvar3561 = (1'h0); (forvar3561 < (1'h1)); forvar3561 = (forvar3561 + (1'h1)))
                    begin
                      reg3562 <= (~(~($unsigned(reg3539) ?
                          (reg3543 ?
                              forvar3549 : reg3435) : $unsigned(reg3447))));
                      reg3563 <= reg3452[(2'h2):(2'h2)];
                      reg3564 <= $signed($unsigned(forvar3527));
                      reg3565 <= (&reg3451[(2'h2):(2'h2)]);
                    end
                  for (forvar3566 = (1'h0); (forvar3566 < (1'h0)); forvar3566 = (forvar3566 + (1'h1)))
                    begin
                      reg3567 <= $unsigned(((^$unsigned((8'ha1))) <= ((forvar3529 << reg3563) & {(8'hb3)})));
                    end
                  reg3568 <= reg3487[(4'h9):(4'h9)];
                end
              else
                begin
                  reg3561 <= $unsigned($unsigned($unsigned($signed(wire3526))));
                  reg3562 <= $signed((((-reg3488) ?
                      (8'hae) : reg3568) < $unsigned($unsigned(forvar3566))));
                  if ($signed($signed({{reg3548}})))
                    begin
                      reg3563 <= $signed($unsigned($signed((8'ha4))));
                      reg3564 <= (reg3534[(1'h0):(1'h0)] != $signed({forvar3527[(2'h3):(2'h2)]}));
                    end
                  else
                    begin
                      reg3563 <= ($unsigned($signed((reg3517 >> reg3557))) ?
                          {reg3451[(1'h1):(1'h0)]} : $unsigned($signed((reg3475 & reg3487))));
                      reg3564 <= reg3530;
                      reg3565 <= {((((8'ha8) ? reg3506 : reg3432) <= (wire3522 ?
                                  reg3475 : reg3510)) ?
                              ((~&wire3525) ?
                                  reg3487[(1'h0):(1'h0)] : {reg3429}) : ($signed(reg3564) < reg3538))};
                      reg3566 <= (|{(|(reg3456 ? reg3510 : reg3460))});
                    end
                  for (forvar3567 = (1'h0); (forvar3567 < (2'h2)); forvar3567 = (forvar3567 + (1'h1)))
                    begin
                      reg3568 <= (^~$unsigned((^(forvar3551 ?
                          (8'haf) : wire3526))));
                      reg3569 <= $unsigned($signed(forvar3567));
                      reg3570 <= ((reg3532[(1'h1):(1'h1)] != $unsigned(((8'ha5) ?
                              reg3472 : reg3449))) ?
                          $unsigned(((reg3565 >= reg3507) ?
                              reg3494[(1'h0):(1'h0)] : (-(8'ha5)))) : reg3508[(3'h7):(3'h6)]);
                    end
                end
              for (forvar3571 = (1'h0); (forvar3571 < (2'h3)); forvar3571 = (forvar3571 + (1'h1)))
                begin
                  if ((~|reg3562[(2'h3):(1'h0)]))
                    begin
                      reg3572 <= reg3452[(1'h0):(1'h0)];
                      reg3573 <= (reg3477[(2'h2):(1'h1)] && reg3572[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg3572 <= (&$signed($signed($signed(reg3490))));
                    end
                  for (forvar3574 = (1'h0); (forvar3574 < (2'h2)); forvar3574 = (forvar3574 + (1'h1)))
                    begin
                      reg3575 <= (^~{reg3521});
                      reg3576 <= $signed($unsigned((!reg3536)));
                    end
                end
            end
          for (forvar3577 = (1'h0); (forvar3577 < (2'h3)); forvar3577 = (forvar3577 + (1'h1)))
            begin
              if (((^~$signed({reg3493})) ?
                  (-reg3535) : (~&reg3492[(3'h6):(2'h2)])))
                begin
                  for (forvar3578 = (1'h0); (forvar3578 < (1'h1)); forvar3578 = (forvar3578 + (1'h1)))
                    begin
                      reg3579 <= forvar3574;
                    end
                  if ($unsigned((^$signed($unsigned(reg3492)))))
                    begin
                      reg3580 <= $signed($signed($signed($unsigned(reg3494))));
                      reg3581 <= $signed(($signed((reg3558 ?
                              (8'hb7) : (8'hb3))) ?
                          reg3432 : (reg3552 == forvar3537[(3'h5):(1'h1)])));
                      reg3582 <= reg3573[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg3580 <= reg3548;
                    end
                end
              else
                begin
                  reg3578 <= reg3467;
                end
              for (forvar3583 = (1'h0); (forvar3583 < (2'h2)); forvar3583 = (forvar3583 + (1'h1)))
                begin
                  if ($signed($unsigned(($signed(reg3446) ^ (reg3444 ?
                      reg3482 : reg3517)))))
                    begin
                      reg3584 <= ({{$unsigned((8'ha4))}} ? reg3555 : reg3441);
                      reg3585 <= (($signed(reg3435) < ({reg3552} ?
                              $signed((8'ha7)) : wire3422)) ?
                          ($unsigned($signed(reg3565)) ?
                              $signed((reg3449 + reg3442)) : reg3501[(2'h2):(1'h1)]) : reg3490);
                      reg3586 <= ($signed(($signed((8'haf)) ?
                              (reg3567 >>> reg3519) : (reg3559 ?
                                  reg3579 : reg3578))) ?
                          $signed(reg3472[(3'h6):(3'h4)]) : $unsigned((reg3568 ^~ (+wire3525))));
                      reg3587 <= reg3508[(4'ha):(1'h0)];
                    end
                  else
                    begin
                      reg3584 <= $unsigned($unsigned((reg3472 ?
                          (8'hac) : $signed(reg3555))));
                      reg3585 <= (reg3543[(1'h0):(1'h0)] ? reg3450 : reg3441);
                      reg3586 <= reg3557[(2'h3):(2'h3)];
                      reg3587 <= {((~&$unsigned(reg3521)) ?
                              (+$unsigned(wire3524)) : ((reg3504 ?
                                  reg3562 : reg3521) << (reg3475 || reg3581)))};
                    end
                  for (forvar3588 = (1'h0); (forvar3588 < (1'h1)); forvar3588 = (forvar3588 + (1'h1)))
                    begin
                      reg3589 <= (!{(reg3508 ? (8'hab) : reg3442)});
                      reg3590 <= $signed($unsigned((+(-reg3557))));
                      reg3591 <= ((forvar3560[(1'h0):(1'h0)] ?
                          reg3569 : ((8'h9e) & $unsigned(wire3426))) + {({reg3486} != (+reg3575))});
                      reg3592 <= ($signed(forvar3529) ?
                          ($unsigned(reg3439) ?
                              reg3460[(3'h4):(1'h0)] : (-reg3481)) : $signed((reg3428[(1'h0):(1'h0)] && reg3585)));
                    end
                  for (forvar3593 = (1'h0); (forvar3593 < (2'h2)); forvar3593 = (forvar3593 + (1'h1)))
                    begin
                      reg3594 <= (|($unsigned((|reg3456)) ?
                          $unsigned({wire3524}) : $signed($unsigned((8'hb6)))));
                      reg3595 <= {$signed((8'haf))};
                    end
                end
              if (($signed(reg3516[(4'ha):(2'h3)]) && $signed(((8'hba) ?
                  reg3455 : $unsigned(reg3451)))))
                begin
                  for (forvar3596 = (1'h0); (forvar3596 < (1'h0)); forvar3596 = (forvar3596 + (1'h1)))
                    begin
                      reg3597 <= reg3566;
                      reg3598 <= (^~(forvar3553[(2'h2):(1'h1)] && (^~(reg3545 ?
                          reg3587 : reg3438))));
                    end
                  for (forvar3599 = (1'h0); (forvar3599 < (1'h0)); forvar3599 = (forvar3599 + (1'h1)))
                    begin
                      reg3600 <= (reg3549 ? {$unsigned((!(8'ha6)))} : reg3440);
                      reg3601 <= reg3432;
                      reg3602 <= (^~{$signed({reg3531})});
                      reg3603 <= $unsigned(((8'hab) > $unsigned(reg3486[(1'h1):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar3596 = (1'h0); (forvar3596 < (1'h0)); forvar3596 = (forvar3596 + (1'h1)))
                    begin
                      reg3597 <= reg3437;
                      reg3598 <= $signed({$unsigned({reg3449})});
                    end
                  if ((~|(($unsigned(reg3581) ?
                          {forvar3599} : (forvar3596 < reg3569)) ?
                      $signed((reg3551 ?
                          forvar3560 : (8'ha4))) : (~|$signed(forvar3528)))))
                    begin
                      reg3599 <= reg3521[(4'hc):(4'hb)];
                      reg3600 <= (reg3556[(1'h1):(1'h1)] > (&wire3425));
                    end
                  else
                    begin
                      reg3599 <= $unsigned($unsigned(reg3466[(1'h1):(1'h1)]));
                      reg3600 <= ((|reg3550[(2'h3):(1'h0)]) ?
                          (($unsigned(reg3439) ?
                                  $unsigned(reg3504) : wire3525[(4'ha):(1'h0)]) ?
                              $signed(reg3507) : ($signed(reg3536) ?
                                  forvar3541 : $signed(reg3590))) : reg3467);
                      reg3601 <= ({$unsigned(reg3563[(2'h3):(2'h3)])} ?
                          $signed(({reg3508} ?
                              ((8'ha3) & reg3530) : (reg3452 >= reg3475))) : ({$unsigned((8'hb0))} ?
                              $signed($unsigned(forvar3593)) : ({reg3441} ?
                                  (+reg3503) : (reg3545 ^~ forvar3561))));
                    end
                end
            end
        end
      else
        begin
          for (forvar3527 = (1'h0); (forvar3527 < (1'h0)); forvar3527 = (forvar3527 + (1'h1)))
            begin
              if ($unsigned(($signed((wire3424 ^ reg3468)) ?
                  $unsigned((~^wire3522)) : (reg3448[(1'h0):(1'h0)] ^~ reg3561[(4'hb):(1'h0)]))))
                begin
                  if ($unsigned(reg3556))
                    begin
                      reg3528 <= reg3498[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg3528 <= wire3425[(4'ha):(4'ha)];
                      reg3529 <= (reg3590 > ({reg3542} ?
                          reg3481 : reg3459[(3'h5):(3'h4)]));
                      reg3530 <= ((~|$unsigned((forvar3567 ?
                          reg3557 : reg3434))) >= (~|($signed(reg3541) || (forvar3571 ?
                          reg3508 : (8'ha3)))));
                      reg3531 <= (~($unsigned((wire3523 < reg3461)) ^~ ((forvar3574 >>> (8'ha2)) ?
                          $unsigned(forvar3537) : wire3522)));
                    end
                  if ({(~&{reg3427[(3'h7):(1'h1)]})})
                    begin
                      reg3532 <= reg3599[(1'h1):(1'h0)];
                      reg3533 <= $signed(reg3549);
                      reg3534 <= $unsigned(((forvar3541 ?
                          reg3586[(2'h2):(1'h0)] : reg3536) || $unsigned(reg3476[(2'h3):(2'h3)])));
                      reg3535 <= (~|{{(reg3445 && forvar3548)}});
                    end
                  else
                    begin
                      reg3532 <= reg3457[(3'h6):(1'h0)];
                      reg3533 <= {$unsigned(((forvar3537 < reg3528) >>> $unsigned(reg3458)))};
                      reg3534 <= $signed($signed($signed((reg3491 & (8'hb1)))));
                      reg3535 <= $unsigned($signed(reg3504));
                    end
                end
              else
                begin
                  if (forvar3528[(2'h2):(1'h1)])
                    begin
                      reg3528 <= ($signed($signed({reg3506})) << (-reg3439[(1'h0):(1'h0)]));
                      reg3529 <= (|$signed((-$unsigned(forvar3553))));
                      reg3530 <= forvar3537[(1'h0):(1'h0)];
                      reg3531 <= (-(8'ha9));
                    end
                  else
                    begin
                      reg3528 <= wire3523;
                      reg3529 <= $signed((8'hb4));
                      reg3530 <= ($signed($signed($signed(reg3492))) ?
                          $signed(reg3498[(2'h2):(2'h2)]) : reg3450[(3'h7):(3'h4)]);
                      reg3531 <= {reg3465[(2'h3):(2'h2)]};
                    end
                  reg3532 <= ((~^$unsigned((reg3482 << reg3493))) & {$unsigned(reg3534[(2'h3):(2'h3)])});
                  reg3533 <= reg3484;
                end
              for (forvar3536 = (1'h0); (forvar3536 < (2'h2)); forvar3536 = (forvar3536 + (1'h1)))
                begin
                  reg3537 <= reg3535;
                  if (((+$unsigned(reg3457)) * forvar3529[(1'h1):(1'h1)]))
                    begin
                      reg3538 <= $signed((~|((reg3537 ?
                          reg3589 : reg3565) || reg3466)));
                      reg3539 <= ($signed(({reg3558} >= forvar3551[(2'h2):(1'h1)])) && ($unsigned(reg3484) ?
                          (reg3542 * reg3455[(4'h9):(1'h0)]) : reg3455[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg3538 <= ($signed(($signed(reg3440) >= ((8'hae) ?
                          wire3424 : (8'hba)))) & ((!(-reg3517)) && ((reg3436 ?
                          reg3533 : reg3533) ^~ $unsigned((8'hb3)))));
                    end
                end
            end
          if ($unsigned((reg3501[(2'h2):(2'h2)] ?
              $unsigned((reg3562 ?
                  reg3463 : reg3569)) : reg3595[(1'h1):(1'h0)])))
            begin
              for (forvar3540 = (1'h0); (forvar3540 < (2'h2)); forvar3540 = (forvar3540 + (1'h1)))
                begin
                  if ((~^(((reg3492 == reg3603) < (~^reg3572)) ?
                      (^((8'hb7) ?
                          (8'hb3) : reg3563)) : $unsigned($unsigned(reg3541)))))
                    begin
                      reg3541 <= $unsigned((reg3433[(4'ha):(4'h8)] ?
                          ($unsigned(reg3507) ?
                              $signed(reg3552) : {reg3602}) : {$signed(reg3436)}));
                    end
                  else
                    begin
                      reg3541 <= ($signed(reg3498) < (forvar3588 == $signed((~|reg3578))));
                      reg3542 <= reg3544;
                      reg3543 <= (({wire3423} ?
                          reg3518 : ($unsigned(reg3576) >>> {reg3429})) & (~|((reg3510 < reg3601) ?
                          ((8'h9d) ? (8'haf) : reg3429) : {forvar3528})));
                    end
                  reg3544 <= (reg3575 ^ (reg3483[(1'h0):(1'h0)] >> $signed($unsigned(reg3475))));
                  for (forvar3545 = (1'h0); (forvar3545 < (2'h3)); forvar3545 = (forvar3545 + (1'h1)))
                    begin
                      reg3546 <= $unsigned($signed((8'hb6)));
                    end
                end
              if (((|$signed((reg3441 == reg3549))) >= {($unsigned(reg3594) || $unsigned(reg3562))}))
                begin
                  if ($signed((~reg3533)))
                    begin
                      reg3547 <= (|(((&reg3451) - (reg3482 ^ reg3556)) & $signed({(8'hb6)})));
                    end
                  else
                    begin
                      reg3547 <= {((^reg3592) & ((reg3545 ?
                              (8'hb1) : reg3556) || $unsigned(reg3548)))};
                      reg3548 <= ($unsigned($unsigned(reg3453[(4'hc):(4'h8)])) - reg3455[(3'h7):(1'h1)]);
                      reg3549 <= (((reg3468 & $unsigned(reg3501)) ?
                          {(wire3522 <= reg3554)} : $signed((reg3536 << reg3557))) * {reg3516});
                    end
                end
              else
                begin
                  if (reg3435)
                    begin
                      reg3547 <= reg3565;
                      reg3548 <= $signed({(~|$signed((8'hb4)))});
                    end
                  else
                    begin
                      reg3547 <= $unsigned(wire3425);
                      reg3548 <= $signed(((&{(8'hba)}) ?
                          ({(8'ha6)} ?
                              (forvar3541 || reg3589) : (reg3456 ^~ reg3532)) : (8'h9e)));
                      reg3549 <= $signed((($unsigned(reg3520) ?
                          (~reg3447) : $unsigned(reg3510)) <<< $unsigned($signed(reg3438))));
                    end
                  reg3550 <= $signed(reg3579);
                  for (forvar3551 = (1'h0); (forvar3551 < (1'h1)); forvar3551 = (forvar3551 + (1'h1)))
                    begin
                      reg3552 <= $signed(($unsigned((+reg3513)) || $unsigned($signed(reg3494))));
                      reg3553 <= (((+reg3469) ?
                          ({reg3456} ?
                              $signed((8'hb2)) : reg3455) : reg3482) && reg3512);
                      reg3554 <= $unsigned($signed((^$unsigned((8'hb4)))));
                    end
                end
              for (forvar3555 = (1'h0); (forvar3555 < (2'h2)); forvar3555 = (forvar3555 + (1'h1)))
                begin
                  if ((~&reg3544))
                    begin
                      reg3556 <= $unsigned((reg3428[(3'h5):(2'h3)] ?
                          ($unsigned(reg3507) ?
                              (reg3512 ?
                                  (8'had) : reg3544) : forvar3548[(1'h1):(1'h0)]) : reg3572[(3'h5):(3'h5)]));
                      reg3557 <= $signed((forvar3571[(2'h3):(1'h0)] ?
                          reg3497[(3'h4):(2'h3)] : reg3567[(2'h3):(2'h3)]));
                      reg3558 <= reg3494;
                      reg3559 <= (~^reg3540[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg3556 <= reg3508[(3'h4):(1'h0)];
                      reg3557 <= (~|{(^reg3470)});
                    end
                end
            end
          else
            begin
              if ((8'hb6))
                begin
                  for (forvar3540 = (1'h0); (forvar3540 < (1'h0)); forvar3540 = (forvar3540 + (1'h1)))
                    begin
                      reg3541 <= {(reg3475 ?
                              {reg3460[(1'h1):(1'h1)]} : (reg3534[(4'h8):(4'h8)] ?
                                  (reg3545 ?
                                      reg3453 : reg3550) : $unsigned(reg3444)))};
                      reg3542 <= ($unsigned({(reg3458 ?
                              (8'ha5) : (8'hb9))}) | ($unsigned((^reg3555)) >= ((8'ha1) ?
                          $signed(reg3433) : (reg3468 ? reg3540 : reg3512))));
                      reg3543 <= (~^(($signed(reg3431) ?
                              (^~forvar3548) : $unsigned((8'hba))) ?
                          $signed(reg3489[(2'h2):(1'h0)]) : {reg3568[(3'h6):(3'h5)]}));
                    end
                  for (forvar3544 = (1'h0); (forvar3544 < (2'h3)); forvar3544 = (forvar3544 + (1'h1)))
                    begin
                      reg3545 <= ({reg3446[(1'h0):(1'h0)]} ?
                          $signed((^~((8'hb8) ?
                              reg3528 : (8'ha3)))) : $signed($unsigned((reg3582 ^ reg3549))));
                      reg3546 <= (8'h9c);
                    end
                  reg3547 <= reg3555;
                end
              else
                begin
                  for (forvar3540 = (1'h0); (forvar3540 < (2'h3)); forvar3540 = (forvar3540 + (1'h1)))
                    begin
                      reg3541 <= (((+{forvar3596}) ?
                          reg3455[(1'h1):(1'h0)] : reg3557[(3'h5):(2'h3)]) * $signed(reg3468));
                      reg3542 <= $signed(({(!forvar3567)} ?
                          ((forvar3529 ? reg3555 : reg3499) ?
                              ((8'hac) ?
                                  (8'ha6) : reg3514) : forvar3537) : reg3602[(4'h8):(3'h6)]));
                      reg3543 <= (((~|(&reg3543)) ?
                          (-(forvar3540 < reg3541)) : ($unsigned((8'haf)) ?
                              (^reg3584) : wire3522)) > (~^$signed(reg3584)));
                      reg3544 <= $signed((8'hac));
                    end
                end
            end
          for (forvar3560 = (1'h0); (forvar3560 < (1'h0)); forvar3560 = (forvar3560 + (1'h1)))
            begin
              for (forvar3561 = (1'h0); (forvar3561 < (1'h0)); forvar3561 = (forvar3561 + (1'h1)))
                begin
                  if (((~((reg3469 ? reg3427 : (8'haf)) ?
                          (forvar3567 ? (8'hb8) : (8'hb0)) : (reg3482 ?
                              forvar3560 : reg3554))) ?
                      $unsigned({(~^(8'had))}) : $signed((~^$unsigned(wire3426)))))
                    begin
                      reg3562 <= {{reg3475}};
                      reg3563 <= wire3522;
                      reg3564 <= (forvar3541 ?
                          ((reg3445 ?
                                  (reg3508 ?
                                      (8'hb7) : reg3511) : (reg3477 > reg3548)) ?
                              reg3446 : $signed($signed(reg3599))) : (^$signed((forvar3561 ?
                              reg3460 : (8'ha7)))));
                    end
                  else
                    begin
                      reg3562 <= (~&($unsigned($unsigned(reg3511)) + $signed((+reg3553))));
                      reg3563 <= (8'hab);
                    end
                  if ((reg3566[(2'h2):(1'h1)] ?
                      (reg3592[(1'h0):(1'h0)] ?
                          forvar3555[(2'h2):(2'h2)] : reg3483[(4'h9):(1'h1)]) : ($signed((forvar3528 && reg3467)) | $signed((reg3507 ?
                          reg3494 : reg3438)))))
                    begin
                      reg3565 <= {(((forvar3571 * (8'ha9)) ?
                                  $unsigned((8'hb4)) : (reg3564 ?
                                      reg3592 : reg3536)) ?
                              $unsigned($signed(reg3437)) : (8'hb1))};
                      reg3566 <= (reg3580[(2'h3):(1'h0)] ? reg3549 : reg3594);
                      reg3567 <= reg3458;
                    end
                  else
                    begin
                      reg3565 <= {(($signed(wire3525) == reg3545[(2'h3):(2'h3)]) - (reg3444 == reg3564))};
                      reg3566 <= (!(&reg3472[(4'h9):(4'h9)]));
                    end
                  for (forvar3568 = (1'h0); (forvar3568 < (2'h3)); forvar3568 = (forvar3568 + (1'h1)))
                    begin
                      reg3569 <= (&(($signed(reg3595) ?
                          reg3536 : (8'had)) <= reg3530[(1'h0):(1'h0)]));
                      reg3570 <= $unsigned(reg3450[(1'h0):(1'h0)]);
                      reg3571 <= $unsigned((~|$signed({reg3550})));
                    end
                  if ((reg3600[(4'hb):(3'h4)] ?
                      ($unsigned($signed((8'hab))) ?
                          (^forvar3545[(2'h3):(2'h2)]) : (!{reg3536})) : reg3455))
                    begin
                      reg3572 <= (($unsigned($unsigned(reg3428)) >= reg3489) ?
                          (&(((8'ha2) >> forvar3593) ?
                              (^~reg3484) : ((8'ha5) ^~ reg3544))) : $unsigned(forvar3561[(4'hc):(4'h9)]));
                      reg3573 <= $signed((+{$signed(reg3484)}));
                    end
                  else
                    begin
                      reg3572 <= $unsigned($unsigned({reg3545[(1'h1):(1'h1)]}));
                      reg3573 <= $unsigned(((((8'ha4) ? reg3546 : reg3487) ?
                              reg3487 : (reg3564 * reg3580)) ?
                          (^(~&wire3425)) : ($unsigned(reg3551) ?
                              (-reg3513) : $unsigned(reg3531))));
                      reg3574 <= reg3569[(4'hd):(3'h4)];
                      reg3575 <= $unsigned({reg3467});
                    end
                end
              reg3576 <= reg3512[(3'h4):(1'h1)];
              for (forvar3577 = (1'h0); (forvar3577 < (1'h1)); forvar3577 = (forvar3577 + (1'h1)))
                begin
                  if ((~^$signed((~(reg3450 > reg3558)))))
                    begin
                      reg3578 <= {$unsigned(reg3499)};
                      reg3579 <= ($unsigned(reg3517) >> reg3574[(1'h0):(1'h0)]);
                      reg3580 <= (($unsigned($signed((8'ha7))) << {(|reg3571)}) ?
                          (~|$signed(forvar3588)) : $unsigned(((~&reg3465) ?
                              $unsigned(reg3530) : (reg3506 > (8'ha3)))));
                    end
                  else
                    begin
                      reg3578 <= reg3490[(2'h2):(2'h2)];
                    end
                  for (forvar3581 = (1'h0); (forvar3581 < (1'h1)); forvar3581 = (forvar3581 + (1'h1)))
                    begin
                      reg3582 <= $unsigned(forvar3551[(2'h2):(2'h2)]);
                      reg3583 <= (forvar3568 ?
                          ((+(reg3539 + (8'hae))) <= $unsigned($signed(forvar3540))) : $unsigned((^~$signed(reg3456))));
                      reg3584 <= ($signed(((&reg3468) ?
                          (+wire3525) : reg3432[(3'h7):(3'h6)])) != $signed((&(reg3547 > (8'hb4)))));
                    end
                  for (forvar3585 = (1'h0); (forvar3585 < (1'h0)); forvar3585 = (forvar3585 + (1'h1)))
                    begin
                      reg3586 <= reg3461;
                    end
                end
              reg3587 <= ($signed(reg3466) | reg3457[(2'h3):(1'h1)]);
            end
        end
      if (reg3441)
        begin
          reg3604 <= (~(^reg3448));
        end
      else
        begin
          for (forvar3604 = (1'h0); (forvar3604 < (2'h3)); forvar3604 = (forvar3604 + (1'h1)))
            begin
              reg3605 <= (reg3491[(3'h4):(2'h3)] ?
                  {(&(-reg3438))} : $unsigned($unsigned($signed(forvar3540))));
              for (forvar3606 = (1'h0); (forvar3606 < (1'h0)); forvar3606 = (forvar3606 + (1'h1)))
                begin
                  for (forvar3607 = (1'h0); (forvar3607 < (1'h1)); forvar3607 = (forvar3607 + (1'h1)))
                    begin
                      reg3608 <= $signed(($unsigned({forvar3537}) && forvar3585[(4'h9):(4'h9)]));
                      reg3609 <= (8'ha2);
                      reg3610 <= (!reg3555);
                    end
                end
              if (reg3489[(1'h0):(1'h0)])
                begin
                  for (forvar3611 = (1'h0); (forvar3611 < (1'h1)); forvar3611 = (forvar3611 + (1'h1)))
                    begin
                      reg3612 <= $signed(($unsigned(reg3435[(4'ha):(2'h2)]) ?
                          reg3451 : reg3600[(1'h1):(1'h1)]));
                      reg3613 <= $signed((((reg3431 ? reg3500 : reg3451) ?
                              $unsigned(reg3567) : forvar3560[(3'h4):(2'h2)]) ?
                          {(~(8'hb1))} : $unsigned((reg3579 ?
                              reg3475 : forvar3607))));
                      reg3614 <= reg3548[(3'h5):(3'h5)];
                    end
                  if ((~&($unsigned($signed(reg3545)) >>> ((reg3533 ?
                          reg3521 : forvar3568) ?
                      {reg3572} : reg3462[(2'h2):(2'h2)]))))
                    begin
                      reg3615 <= (forvar3588[(1'h1):(1'h0)] ~^ (forvar3607 ?
                          (~reg3592[(3'h4):(1'h0)]) : $signed(reg3601[(3'h4):(1'h0)])));
                    end
                  else
                    begin
                      reg3615 <= ({(reg3490 ^ $signed(reg3544))} ~^ $signed(reg3449[(4'hc):(2'h3)]));
                      reg3616 <= ($signed(((reg3595 << (8'hb5)) ?
                              {(8'haf)} : forvar3578[(3'h7):(2'h2)])) ?
                          (reg3564[(1'h1):(1'h0)] >>> (8'hb9)) : reg3539[(3'h5):(1'h1)]);
                      reg3617 <= ((!((~|reg3453) ?
                          reg3427 : reg3468)) >> reg3429[(3'h4):(2'h3)]);
                      reg3618 <= reg3539[(2'h2):(2'h2)];
                    end
                end
              else
                begin
                  if ($signed(($unsigned((^reg3581)) ?
                      reg3567[(3'h7):(1'h1)] : ((forvar3560 >= reg3550) >> forvar3578))))
                    begin
                      reg3611 <= ($signed($unsigned(reg3570)) ?
                          (reg3439[(2'h3):(1'h1)] ?
                              {$unsigned(wire3526)} : $signed($signed(wire3523))) : (^~{$unsigned(reg3546)}));
                    end
                  else
                    begin
                      reg3611 <= ($signed((reg3509 ?
                              $signed(forvar3528) : reg3550[(4'ha):(3'h7)])) ?
                          $signed(reg3581[(4'ha):(2'h2)]) : ($signed((~|forvar3537)) ?
                              (~|{reg3486}) : $unsigned((~|reg3458))));
                      reg3612 <= reg3476[(2'h2):(1'h0)];
                      reg3613 <= $unsigned({(^$unsigned(forvar3555))});
                      reg3614 <= (^~($signed(reg3571) ?
                          ((wire3523 ?
                              forvar3544 : (8'h9f)) <<< $signed(wire3526)) : $unsigned((8'hb0))));
                    end
                  if ((8'hb1))
                    begin
                      reg3615 <= (reg3618[(4'h8):(2'h3)] << (-reg3487));
                    end
                  else
                    begin
                      reg3615 <= $signed($signed($unsigned(reg3510[(3'h4):(2'h3)])));
                      reg3616 <= ($signed((reg3598 ?
                              reg3530[(3'h5):(1'h0)] : reg3465[(1'h0):(1'h0)])) ?
                          ($unsigned($signed(reg3458)) - reg3461[(3'h6):(3'h5)]) : {({(8'h9c)} ?
                                  reg3538[(2'h3):(2'h2)] : {reg3476})});
                    end
                  reg3617 <= $unsigned(reg3461);
                  reg3618 <= (+($unsigned(reg3428[(4'ha):(3'h5)]) >>> ((~forvar3549) <<< reg3481[(3'h4):(3'h4)])));
                end
            end
          reg3619 <= reg3452;
        end
      for (forvar3620 = (1'h0); (forvar3620 < (2'h2)); forvar3620 = (forvar3620 + (1'h1)))
        begin
          for (forvar3621 = (1'h0); (forvar3621 < (1'h0)); forvar3621 = (forvar3621 + (1'h1)))
            begin
              if ($signed(forvar3578))
                begin
                  for (forvar3622 = (1'h0); (forvar3622 < (1'h0)); forvar3622 = (forvar3622 + (1'h1)))
                    begin
                      reg3623 <= {(&reg3595[(1'h1):(1'h0)])};
                    end
                  for (forvar3624 = (1'h0); (forvar3624 < (2'h3)); forvar3624 = (forvar3624 + (1'h1)))
                    begin
                      reg3625 <= wire3526[(3'h4):(2'h3)];
                      reg3626 <= forvar3585[(4'h8):(4'h8)];
                      reg3627 <= wire3424[(3'h6):(1'h0)];
                    end
                  reg3628 <= (8'hb8);
                end
              else
                begin
                  for (forvar3622 = (1'h0); (forvar3622 < (1'h0)); forvar3622 = (forvar3622 + (1'h1)))
                    begin
                      reg3623 <= (wire3524[(2'h2):(1'h1)] > ((((8'hba) ?
                              (8'h9e) : reg3563) && $signed((8'ha3))) ?
                          (reg3535[(1'h0):(1'h0)] + reg3489[(1'h1):(1'h1)]) : reg3550[(3'h7):(2'h3)]));
                      reg3624 <= reg3461;
                    end
                  reg3625 <= (reg3610[(2'h2):(1'h0)] ?
                      reg3616[(3'h5):(2'h3)] : ((^$unsigned(reg3512)) + reg3514));
                end
              for (forvar3629 = (1'h0); (forvar3629 < (2'h3)); forvar3629 = (forvar3629 + (1'h1)))
                begin
                  if ((reg3569[(4'he):(1'h1)] ?
                      forvar3561 : $unsigned(reg3458)))
                    begin
                      reg3630 <= (({(reg3499 ?
                              reg3561 : forvar3585)} ^ $signed(reg3582[(2'h3):(2'h3)])) * $unsigned({$signed(reg3627)}));
                      reg3631 <= $unsigned((reg3614 ?
                          reg3499[(3'h4):(1'h1)] : forvar3555[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg3630 <= $signed($unsigned($signed($signed((8'hab)))));
                      reg3631 <= $signed($unsigned(((reg3619 ^ reg3461) ^ $signed((8'h9d)))));
                      reg3632 <= (reg3566[(1'h0):(1'h0)] ?
                          {(|reg3447)} : (reg3444 <<< (+{reg3550})));
                      reg3633 <= (~^(reg3579[(2'h2):(1'h0)] ?
                          $unsigned((8'ha0)) : reg3580[(2'h3):(1'h1)]));
                    end
                end
            end
          reg3634 <= (8'had);
        end
      if (reg3633[(3'h5):(3'h5)])
        begin
          if ((^$unsigned(((reg3478 ? wire3422 : (8'hb2)) ?
              $unsigned(reg3580) : $signed(reg3615)))))
            begin
              for (forvar3635 = (1'h0); (forvar3635 < (2'h2)); forvar3635 = (forvar3635 + (1'h1)))
                begin
                  for (forvar3636 = (1'h0); (forvar3636 < (2'h3)); forvar3636 = (forvar3636 + (1'h1)))
                    begin
                      reg3637 <= (reg3477[(2'h2):(1'h1)] - $unsigned($signed(reg3594)));
                      reg3638 <= ({{reg3576}} ?
                          (forvar3620[(5'h10):(3'h6)] ~^ ($unsigned((8'ha5)) ?
                              {forvar3527} : $signed(reg3632))) : (+(!$unsigned(reg3594))));
                    end
                  if ((-((|(8'h9c)) ?
                      forvar3560 : ((^reg3446) ? {(8'ha1)} : {reg3501}))))
                    begin
                      reg3639 <= (~($unsigned(reg3448[(1'h0):(1'h0)]) ?
                          reg3451[(1'h0):(1'h0)] : reg3599[(3'h7):(2'h3)]));
                      reg3640 <= $signed((^~(((8'hab) - reg3508) << ((8'hb7) >= reg3429))));
                    end
                  else
                    begin
                      reg3639 <= $signed({reg3591[(2'h3):(1'h1)]});
                      reg3640 <= (~reg3632[(3'h4):(1'h0)]);
                    end
                end
              if ((|forvar3545))
                begin
                  for (forvar3641 = (1'h0); (forvar3641 < (1'h1)); forvar3641 = (forvar3641 + (1'h1)))
                    begin
                      reg3642 <= (8'hb6);
                      reg3643 <= {$unsigned(({reg3575} >>> (!reg3531)))};
                    end
                  reg3644 <= reg3508;
                  if ($unsigned(((^~(&reg3478)) ?
                      wire3423 : (~|$signed(reg3634)))))
                    begin
                      reg3645 <= reg3492[(1'h1):(1'h1)];
                      reg3646 <= $unsigned($unsigned($unsigned($signed(reg3630))));
                    end
                  else
                    begin
                      reg3645 <= (~&reg3491[(1'h0):(1'h0)]);
                      reg3646 <= $unsigned(reg3457);
                      reg3647 <= reg3488;
                      reg3648 <= $unsigned($unsigned(((8'hb2) & reg3448)));
                    end
                  for (forvar3649 = (1'h0); (forvar3649 < (1'h1)); forvar3649 = (forvar3649 + (1'h1)))
                    begin
                      reg3650 <= ((-((forvar3536 ?
                              reg3467 : reg3501) <<< ((8'hb7) | reg3566))) ?
                          (((reg3446 ? reg3433 : reg3645) ?
                                  forvar3607 : (reg3643 > reg3573)) ?
                              ((!forvar3588) || reg3456[(3'h4):(1'h0)]) : wire3522[(4'hd):(1'h0)]) : {$signed((!reg3542))});
                    end
                end
              else
                begin
                  if ($signed($unsigned((~^reg3512))))
                    begin
                      reg3641 <= $unsigned((reg3537[(2'h2):(1'h1)] >>> reg3468));
                      reg3642 <= $signed((($unsigned(forvar3599) != $unsigned(reg3447)) >= $unsigned((^~(8'ha1)))));
                    end
                  else
                    begin
                      reg3641 <= {$signed($signed((-(8'ha7))))};
                      reg3642 <= (~|($unsigned(reg3483[(3'h5):(3'h4)]) + forvar3606));
                    end
                  reg3643 <= reg3439;
                  reg3644 <= reg3494[(1'h0):(1'h0)];
                end
            end
          else
            begin
              if ((~(^$signed(forvar3599))))
                begin
                  for (forvar3635 = (1'h0); (forvar3635 < (1'h0)); forvar3635 = (forvar3635 + (1'h1)))
                    begin
                      reg3636 <= reg3475[(1'h1):(1'h1)];
                      reg3637 <= (($signed((~&reg3556)) ?
                          ((wire3422 >> reg3442) + reg3459[(3'h5):(1'h1)]) : ((reg3570 ?
                              (8'haf) : forvar3596) | (reg3472 ?
                              (8'hac) : forvar3527))) && $signed(reg3551));
                      reg3638 <= forvar3636;
                      reg3639 <= (&($unsigned((^forvar3566)) && (((8'hba) ?
                          wire3423 : reg3442) < $unsigned(reg3516))));
                    end
                  if (reg3594)
                    begin
                      reg3640 <= ($unsigned({reg3549}) ?
                          $unsigned(reg3486) : reg3632);
                      reg3641 <= ($unsigned(reg3616[(3'h5):(3'h5)]) ?
                          (({(8'h9e)} ?
                                  (~^forvar3611) : (reg3535 <<< reg3438)) ?
                              ($unsigned(reg3439) > $unsigned(reg3454)) : {$signed(reg3477)}) : ($unsigned($signed(reg3613)) + $signed((&reg3536))));
                      reg3642 <= $unsigned((reg3516[(3'h5):(1'h1)] != $signed(reg3552[(1'h0):(1'h0)])));
                      reg3643 <= reg3482[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3640 <= (forvar3596[(2'h3):(1'h1)] ?
                          $signed({$signed(reg3636)}) : $signed(reg3552));
                      reg3641 <= ($signed(forvar3574) ~^ reg3545[(2'h3):(2'h2)]);
                      reg3642 <= $signed(reg3624);
                    end
                  reg3644 <= $unsigned((((8'hb9) + forvar3606) && ((~^reg3601) ?
                      (reg3645 ? reg3633 : (8'hb8)) : $signed(reg3497))));
                  for (forvar3645 = (1'h0); (forvar3645 < (2'h2)); forvar3645 = (forvar3645 + (1'h1)))
                    begin
                      reg3646 <= ($signed(((+reg3437) - ((8'had) + reg3569))) ?
                          $signed(($unsigned(reg3428) - reg3431[(4'hc):(4'h8)])) : $signed($signed($unsigned(reg3470))));
                      reg3647 <= $signed(reg3638);
                      reg3648 <= ((~|($signed((8'ha3)) ~^ (8'ha1))) == $unsigned(((forvar3588 ?
                              reg3462 : reg3548) ?
                          {reg3639} : ((8'haa) ^~ reg3637))));
                      reg3649 <= (-reg3615[(3'h7):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar3635 = (1'h0); (forvar3635 < (1'h0)); forvar3635 = (forvar3635 + (1'h1)))
                    begin
                      reg3636 <= (reg3546 ?
                          reg3487 : $unsigned(((reg3555 == reg3575) ?
                              (-reg3648) : (reg3437 + reg3529))));
                      reg3637 <= reg3639;
                    end
                  for (forvar3638 = (1'h0); (forvar3638 < (2'h2)); forvar3638 = (forvar3638 + (1'h1)))
                    begin
                      reg3639 <= (~^{forvar3622});
                      reg3640 <= reg3643[(3'h7):(3'h7)];
                      reg3641 <= (&$unsigned((forvar3593[(1'h0):(1'h0)] != (reg3544 ?
                          (8'hac) : reg3591))));
                    end
                  for (forvar3642 = (1'h0); (forvar3642 < (2'h3)); forvar3642 = (forvar3642 + (1'h1)))
                    begin
                      reg3643 <= $unsigned((((forvar3629 >= (8'hb3)) & reg3550[(4'hf):(3'h7)]) < (|forvar3571)));
                      reg3644 <= ((^(reg3592[(3'h5):(3'h5)] + reg3439)) ?
                          reg3597 : $signed(((reg3640 ?
                              forvar3649 : reg3507) ~^ (reg3608 ?
                              (8'ha1) : reg3517))));
                      reg3645 <= $unsigned((((forvar3574 <= reg3643) ?
                              (forvar3560 & forvar3551) : reg3630[(3'h5):(2'h3)]) ?
                          reg3514 : (forvar3638 ?
                              (reg3552 <<< reg3481) : reg3614[(4'h8):(4'h8)])));
                    end
                end
              for (forvar3650 = (1'h0); (forvar3650 < (1'h1)); forvar3650 = (forvar3650 + (1'h1)))
                begin
                  if ($signed(($signed(forvar3528) ^ forvar3620)))
                    begin
                      reg3651 <= reg3597[(1'h1):(1'h0)];
                      reg3652 <= (forvar3536[(2'h3):(2'h2)] ?
                          ($unsigned($signed(reg3649)) ?
                              $signed((^~reg3492)) : $signed($unsigned(reg3439))) : forvar3555);
                      reg3653 <= ((!$signed($unsigned(reg3529))) << reg3568[(3'h6):(2'h3)]);
                    end
                  else
                    begin
                      reg3651 <= (-(|($signed(reg3499) >> reg3506[(4'h9):(3'h6)])));
                    end
                  if (($unsigned(reg3632[(4'h9):(1'h0)]) <= ({$unsigned(reg3456)} >>> reg3564)))
                    begin
                      reg3654 <= ((reg3442[(3'h6):(2'h3)] ~^ $unsigned($unsigned(forvar3621))) < ($unsigned(wire3424) ?
                          ((^reg3580) ?
                              reg3538 : (reg3462 ?
                                  reg3431 : reg3585)) : ($signed(forvar3629) ?
                              (~|reg3430) : (forvar3553 >> reg3517))));
                      reg3655 <= $signed({(8'ha2)});
                      reg3656 <= (~&(^((reg3493 ? reg3533 : reg3605) ?
                          reg3507 : $signed(reg3652))));
                      reg3657 <= $unsigned($signed(((~|(8'hb6)) ?
                          (|(8'ha5)) : (reg3491 ? reg3600 : reg3436))));
                    end
                  else
                    begin
                      reg3654 <= {reg3557};
                      reg3655 <= ({(!(8'ha3))} ?
                          ($signed($signed(reg3540)) ?
                              reg3602 : {(+reg3536)}) : $signed(reg3603));
                      reg3656 <= reg3582;
                      reg3657 <= ((~&reg3429) < forvar3536);
                    end
                  for (forvar3658 = (1'h0); (forvar3658 < (2'h3)); forvar3658 = (forvar3658 + (1'h1)))
                    begin
                      reg3659 <= (8'hb2);
                    end
                end
            end
          if (reg3544[(4'hb):(3'h4)])
            begin
              for (forvar3660 = (1'h0); (forvar3660 < (1'h0)); forvar3660 = (forvar3660 + (1'h1)))
                begin
                  if ($signed((reg3517 ?
                      $signed((forvar3660 ? reg3563 : reg3478)) : ((reg3630 ?
                              reg3605 : reg3569) ?
                          $unsigned(forvar3537) : (reg3438 >> reg3558)))))
                    begin
                      reg3661 <= ((8'ha8) < $unsigned(reg3649));
                    end
                  else
                    begin
                      reg3661 <= ((~|$signed($signed((8'hb2)))) >= $unsigned(((~|reg3630) ?
                          $unsigned(reg3642) : {reg3501})));
                    end
                end
              for (forvar3662 = (1'h0); (forvar3662 < (2'h2)); forvar3662 = (forvar3662 + (1'h1)))
                begin
                  for (forvar3663 = (1'h0); (forvar3663 < (1'h1)); forvar3663 = (forvar3663 + (1'h1)))
                    begin
                      reg3664 <= (~^(((~reg3481) ^~ forvar3536[(2'h2):(1'h0)]) & $signed($signed((8'hb5)))));
                      reg3665 <= reg3559;
                    end
                  for (forvar3666 = (1'h0); (forvar3666 < (1'h0)); forvar3666 = (forvar3666 + (1'h1)))
                    begin
                      reg3667 <= reg3601;
                      reg3668 <= forvar3548;
                      reg3669 <= {(~&($signed(reg3618) ?
                              $unsigned(reg3536) : $unsigned(reg3470)))};
                    end
                  for (forvar3670 = (1'h0); (forvar3670 < (2'h3)); forvar3670 = (forvar3670 + (1'h1)))
                    begin
                      reg3671 <= ($unsigned(reg3434[(1'h1):(1'h0)]) ?
                          reg3618 : reg3625);
                      reg3672 <= ((((forvar3536 <= forvar3553) <<< reg3472) ^ $signed({forvar3566})) + reg3585[(3'h4):(1'h1)]);
                      reg3673 <= (((&(reg3457 + reg3569)) >= (|$unsigned(reg3581))) ?
                          wire3425[(4'h9):(4'h9)] : ({{reg3463}} || reg3602[(3'h7):(2'h3)]));
                    end
                  for (forvar3674 = (1'h0); (forvar3674 < (1'h1)); forvar3674 = (forvar3674 + (1'h1)))
                    begin
                      reg3675 <= ((8'h9d) == ($signed($unsigned(reg3667)) ~^ (-(reg3656 ?
                          reg3428 : reg3548))));
                    end
                end
            end
          else
            begin
              if (({reg3571[(3'h4):(3'h4)]} & reg3639[(2'h2):(1'h0)]))
                begin
                  for (forvar3660 = (1'h0); (forvar3660 < (2'h3)); forvar3660 = (forvar3660 + (1'h1)))
                    begin
                      reg3661 <= ((((^forvar3650) ? reg3634 : forvar3537) ?
                          reg3570 : ((&(8'hae)) | {reg3580})) || ($unsigned($signed(reg3517)) ~^ (^(reg3452 ?
                          reg3491 : (8'ha4)))));
                      reg3662 <= (~^{reg3562});
                      reg3663 <= (~^$signed(reg3605));
                    end
                  if (reg3461)
                    begin
                      reg3664 <= reg3665[(4'h9):(3'h4)];
                      reg3665 <= ({{$unsigned((8'hb1))}} ?
                          (-$unsigned($signed(wire3423))) : ($unsigned((8'ha0)) ?
                              reg3556[(2'h2):(1'h1)] : wire3526));
                      reg3666 <= $unsigned(((~|reg3630) ?
                          ({reg3543} ?
                              $signed(forvar3544) : (reg3519 + reg3583)) : $signed(reg3584[(3'h6):(3'h4)])));
                    end
                  else
                    begin
                      reg3664 <= (^$unsigned((reg3537 & $signed(reg3506))));
                      reg3665 <= ((&$unsigned(reg3673[(4'h9):(2'h2)])) ?
                          ($signed(reg3542[(1'h0):(1'h0)]) ^ $unsigned((reg3440 || reg3598))) : forvar3642[(3'h4):(1'h0)]);
                      reg3666 <= reg3576;
                    end
                end
              else
                begin
                  if ($signed(((((8'ha9) <<< (8'ha1)) <<< reg3582) ?
                      $unsigned((8'ha7)) : ({(8'hb3)} >> reg3557[(1'h1):(1'h0)]))))
                    begin
                      reg3660 <= $signed(forvar3666[(4'hf):(2'h2)]);
                    end
                  else
                    begin
                      reg3660 <= (~(~$unsigned((reg3439 ?
                          reg3487 : forvar3545))));
                      reg3661 <= $unsigned($unsigned({(reg3556 >= forvar3641)}));
                      reg3662 <= reg3448[(1'h0):(1'h0)];
                    end
                  for (forvar3663 = (1'h0); (forvar3663 < (2'h2)); forvar3663 = (forvar3663 + (1'h1)))
                    begin
                      reg3664 <= (reg3645[(1'h0):(1'h0)] ^~ reg3673);
                    end
                  for (forvar3665 = (1'h0); (forvar3665 < (1'h0)); forvar3665 = (forvar3665 + (1'h1)))
                    begin
                      reg3666 <= (wire3522[(1'h0):(1'h0)] & ($unsigned(reg3633) & reg3520));
                      reg3667 <= ($signed(($unsigned(reg3576) | reg3544)) ?
                          (reg3469[(4'ha):(4'h8)] | (reg3509 - (~&reg3613))) : (^~((-forvar3571) ?
                              (~&reg3611) : reg3489[(2'h2):(1'h0)])));
                    end
                  for (forvar3668 = (1'h0); (forvar3668 < (1'h1)); forvar3668 = (forvar3668 + (1'h1)))
                    begin
                      reg3669 <= (|(forvar3548[(2'h2):(1'h1)] <= (reg3475[(2'h3):(1'h1)] >= forvar3665[(3'h6):(2'h2)])));
                      reg3670 <= {$unsigned($unsigned((reg3499 <= reg3431)))};
                    end
                end
              for (forvar3671 = (1'h0); (forvar3671 < (1'h1)); forvar3671 = (forvar3671 + (1'h1)))
                begin
                  for (forvar3672 = (1'h0); (forvar3672 < (2'h3)); forvar3672 = (forvar3672 + (1'h1)))
                    begin
                      reg3673 <= (((8'hb0) ~^ $signed($unsigned(reg3634))) ?
                          $signed($signed($unsigned(reg3506))) : (reg3438 & reg3492));
                      reg3674 <= forvar3541[(3'h4):(1'h0)];
                      reg3675 <= $signed(forvar3672);
                      reg3676 <= $signed($signed(((&forvar3641) <<< (forvar3560 ?
                          reg3510 : reg3617))));
                    end
                  for (forvar3677 = (1'h0); (forvar3677 < (1'h0)); forvar3677 = (forvar3677 + (1'h1)))
                    begin
                      reg3678 <= (((|(reg3468 & reg3519)) ?
                              ((reg3669 >= reg3500) ?
                                  (!reg3462) : ((8'h9e) || reg3434)) : $unsigned($unsigned(reg3562))) ?
                          (($unsigned(reg3516) ?
                                  $signed(reg3444) : (reg3466 + reg3672)) ?
                              reg3458[(1'h0):(1'h0)] : (^(reg3565 & reg3476))) : ((!(forvar3629 ?
                                  reg3535 : (8'hac))) ?
                              $unsigned((forvar3604 ?
                                  forvar3622 : forvar3537)) : (reg3594 - (8'hb3))));
                      reg3679 <= ((reg3568 <<< (|(reg3510 >> reg3467))) ?
                          forvar3560 : ($unsigned(reg3572[(4'hc):(4'h8)]) ?
                              (forvar3537[(3'h7):(3'h7)] ?
                                  (~^reg3615) : (8'ha7)) : ($signed(reg3589) > reg3464[(1'h1):(1'h0)])));
                      reg3680 <= reg3627;
                    end
                end
              if ($signed(reg3679[(3'h5):(1'h1)]))
                begin
                  for (forvar3681 = (1'h0); (forvar3681 < (1'h1)); forvar3681 = (forvar3681 + (1'h1)))
                    begin
                      reg3682 <= (({$signed(reg3648)} ?
                          ((reg3487 && reg3675) || (reg3488 ?
                              reg3556 : forvar3555)) : forvar3662) << (~&($unsigned((8'h9d)) ?
                          (~|reg3540) : reg3507[(1'h1):(1'h0)])));
                      reg3683 <= (+reg3511[(1'h1):(1'h1)]);
                    end
                  for (forvar3684 = (1'h0); (forvar3684 < (1'h0)); forvar3684 = (forvar3684 + (1'h1)))
                    begin
                      reg3685 <= reg3511[(1'h0):(1'h0)];
                      reg3686 <= (reg3554[(4'ha):(3'h7)] >>> (($signed(reg3548) || $signed(reg3633)) ?
                          $unsigned((reg3451 * reg3591)) : {reg3623[(1'h1):(1'h1)]}));
                    end
                  reg3687 <= $signed($signed((((8'ha5) ?
                          forvar3581 : forvar3577) ?
                      {reg3680} : (&reg3472))));
                end
              else
                begin
                  if ($unsigned((reg3487[(4'hd):(4'hd)] - (8'hba))))
                    begin
                      reg3681 <= $signed(reg3450[(3'h7):(3'h6)]);
                      reg3682 <= reg3662[(3'h4):(2'h3)];
                      reg3683 <= reg3652;
                      reg3684 <= $signed((8'hb5));
                    end
                  else
                    begin
                      reg3681 <= $signed((($unsigned(forvar3635) ?
                          {forvar3642} : reg3490[(1'h0):(1'h0)]) ~^ ({reg3513} ?
                          forvar3571[(3'h4):(2'h2)] : {forvar3599})));
                      reg3682 <= forvar3596;
                    end
                  for (forvar3685 = (1'h0); (forvar3685 < (1'h1)); forvar3685 = (forvar3685 + (1'h1)))
                    begin
                      reg3686 <= {forvar3536};
                      reg3687 <= $signed((&reg3616));
                      reg3688 <= (8'h9e);
                    end
                  if (((((reg3531 ? reg3514 : forvar3622) & (reg3562 ?
                              forvar3636 : reg3565)) ?
                          $unsigned($signed(reg3464)) : (wire3526 ?
                              reg3626[(1'h1):(1'h0)] : $unsigned(forvar3604))) ?
                      $unsigned($signed((reg3634 - forvar3681))) : {(|reg3580)}))
                    begin
                      reg3689 <= (~|({$signed(reg3628)} ?
                          {$unsigned(reg3669)} : reg3688));
                      reg3690 <= reg3547[(3'h4):(2'h3)];
                      reg3691 <= $unsigned(reg3455);
                    end
                  else
                    begin
                      reg3689 <= {(!$unsigned($signed(forvar3548)))};
                    end
                  reg3692 <= (~|(reg3558[(4'hd):(3'h6)] ?
                      reg3558[(3'h7):(2'h2)] : (((8'ha2) >= reg3683) != $signed(reg3490))));
                end
            end
          reg3693 <= reg3465;
          for (forvar3694 = (1'h0); (forvar3694 < (1'h0)); forvar3694 = (forvar3694 + (1'h1)))
            begin
              for (forvar3695 = (1'h0); (forvar3695 < (2'h3)); forvar3695 = (forvar3695 + (1'h1)))
                begin
                  for (forvar3696 = (1'h0); (forvar3696 < (1'h0)); forvar3696 = (forvar3696 + (1'h1)))
                    begin
                      reg3697 <= reg3657[(1'h0):(1'h0)];
                      reg3698 <= (|{reg3664});
                      reg3699 <= reg3474;
                      reg3700 <= forvar3641[(3'h6):(1'h1)];
                    end
                  if ($signed($unsigned(reg3447[(2'h2):(1'h0)])))
                    begin
                      reg3701 <= reg3466[(1'h1):(1'h1)];
                      reg3702 <= $signed({(&(&wire3525))});
                      reg3703 <= ((~{reg3557[(3'h6):(3'h4)]}) > reg3602[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg3701 <= ((8'ha0) ?
                          $signed($unsigned((forvar3694 ~^ reg3549))) : reg3462[(3'h7):(2'h3)]);
                      reg3702 <= {$signed(((8'ha3) ?
                              ((8'hb5) ?
                                  reg3597 : reg3546) : $unsigned(forvar3611)))};
                    end
                end
              if ({$signed(reg3623[(3'h6):(3'h4)])})
                begin
                  for (forvar3704 = (1'h0); (forvar3704 < (2'h2)); forvar3704 = (forvar3704 + (1'h1)))
                    begin
                      reg3705 <= ({(-{reg3470})} <= (reg3651[(3'h7):(1'h0)] - (reg3610[(1'h0):(1'h0)] ?
                          $signed((8'h9c)) : (forvar3567 ?
                              reg3689 : forvar3624))));
                      reg3706 <= (reg3681[(3'h5):(3'h4)] ?
                          $unsigned((8'hb6)) : (((forvar3629 ?
                                      forvar3599 : reg3644) ?
                                  reg3476 : (reg3570 ? reg3546 : (8'hb4))) ?
                              forvar3611[(1'h1):(1'h0)] : ({reg3634} ?
                                  reg3705[(4'h9):(3'h5)] : ((8'h9d) >> forvar3585))));
                      reg3707 <= $unsigned(($unsigned({reg3599}) ?
                          $unsigned({reg3666}) : ($signed(reg3432) ?
                              $unsigned(reg3481) : reg3434[(2'h2):(1'h1)])));
                    end
                  for (forvar3708 = (1'h0); (forvar3708 < (1'h0)); forvar3708 = (forvar3708 + (1'h1)))
                    begin
                      reg3709 <= $unsigned((8'hb7));
                      reg3710 <= ((reg3431 ^~ (reg3564 ?
                          forvar3577 : (reg3569 ?
                              forvar3668 : reg3636))) * (((8'hae) >> (reg3581 ^~ reg3661)) ?
                          (!(8'hb0)) : reg3539));
                    end
                  reg3711 <= $unsigned(((reg3531 ?
                          {reg3439} : (wire3425 ^~ (8'ha0))) ?
                      ($signed(reg3707) || $signed(reg3488)) : (^~(8'hb6))));
                end
              else
                begin
                  if ((forvar3528[(1'h1):(1'h0)] ?
                      ({forvar3704} ?
                          $signed((8'ha7)) : wire3425[(4'h8):(3'h7)]) : $signed($signed(forvar3695))))
                    begin
                      reg3704 <= (~&reg3674);
                      reg3705 <= forvar3599[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg3704 <= $unsigned((((reg3610 ?
                                  forvar3677 : forvar3695) ?
                              (forvar3528 > reg3445) : (&reg3616)) ?
                          ($signed((8'hb2)) ?
                              forvar3704[(1'h1):(1'h0)] : $unsigned(wire3422)) : reg3640[(1'h1):(1'h1)]));
                    end
                  if ({$signed($unsigned(forvar3541[(2'h2):(1'h0)]))})
                    begin
                      reg3706 <= $signed($signed($unsigned((8'h9e))));
                      reg3707 <= (-{((reg3646 - reg3442) ?
                              (~&reg3665) : $signed(forvar3574))});
                      reg3708 <= ($unsigned(($unsigned(reg3511) & (reg3592 >= reg3563))) ?
                          (!(~^{forvar3681})) : $unsigned((!forvar3578)));
                    end
                  else
                    begin
                      reg3706 <= (forvar3581 ?
                          {reg3608[(4'h9):(3'h6)]} : (reg3663[(4'ha):(3'h4)] ?
                              $signed(reg3589) : $signed((~|(8'ha1)))));
                    end
                end
              reg3712 <= (~|$signed(reg3442[(4'hf):(4'h8)]));
            end
        end
      else
        begin
          reg3635 <= $signed((reg3655 ^~ ($signed(forvar3545) >> reg3499)));
        end
    end
  assign wire3713 = reg3555;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3936  (y, clk, wire3941, wire3940, wire3939, wire3938, wire3937);
  output wire [(32'hc39):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire3941;
  input wire [(2'h2):(1'h0)] wire3940;
  input wire signed [(3'h6):(1'h0)] wire3939;
  input wire [(3'h4):(1'h0)] wire3938;
  input wire signed [(3'h7):(1'h0)] wire3937;
  wire signed [(2'h2):(1'h0)] wire4538;
  wire signed [(4'hb):(1'h0)] wire4537;
  wire [(4'he):(1'h0)] wire4536;
  wire signed [(5'h10):(1'h0)] wire4535;
  wire signed [(4'hf):(1'h0)] wire4533;
  wire signed [(2'h3):(1'h0)] wire4213;
  wire signed [(3'h4):(1'h0)] wire4212;
  wire signed [(3'h4):(1'h0)] wire3944;
  wire signed [(3'h5):(1'h0)] wire3943;
  wire [(4'he):(1'h0)] wire3942;
  reg signed [(5'h10):(1'h0)] reg4126 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4211 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4210 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4208 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4207 = (1'h0);
  reg [(2'h2):(1'h0)] reg4205 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4206 = (1'h0);
  reg [(4'hb):(1'h0)] reg4204 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4203 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4202 = (1'h0);
  reg [(4'h9):(1'h0)] reg4200 = (1'h0);
  reg [(2'h3):(1'h0)] reg4199 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4198 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4194 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4196 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4195 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4193 = (1'h0);
  reg [(4'h9):(1'h0)] reg4153 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4148 = (1'h0);
  reg [(2'h3):(1'h0)] reg4191 = (1'h0);
  reg [(4'hf):(1'h0)] reg4190 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4189 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4188 = (1'h0);
  reg [(3'h7):(1'h0)] reg4187 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4185 = (1'h0);
  reg [(4'h9):(1'h0)] reg4184 = (1'h0);
  reg [(4'he):(1'h0)] reg4183 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4182 = (1'h0);
  reg [(4'hf):(1'h0)] reg4181 = (1'h0);
  reg [(4'ha):(1'h0)] reg4180 = (1'h0);
  reg [(4'hf):(1'h0)] reg4178 = (1'h0);
  reg [(4'hb):(1'h0)] reg4177 = (1'h0);
  reg [(4'hf):(1'h0)] reg4176 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4175 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4174 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4172 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4169 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4167 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4166 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4165 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4164 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4158 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4163 = (1'h0);
  reg [(3'h7):(1'h0)] reg4162 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4161 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4160 = (1'h0);
  reg [(4'ha):(1'h0)] reg4159 = (1'h0);
  reg [(2'h2):(1'h0)] reg4157 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4156 = (1'h0);
  reg [(4'h9):(1'h0)] reg4155 = (1'h0);
  reg [(4'hd):(1'h0)] reg4154 = (1'h0);
  reg [(4'hb):(1'h0)] reg4152 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4151 = (1'h0);
  reg [(4'h9):(1'h0)] reg4150 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4149 = (1'h0);
  reg [(3'h4):(1'h0)] reg4147 = (1'h0);
  reg [(3'h4):(1'h0)] reg4144 = (1'h0);
  reg [(4'h9):(1'h0)] reg4146 = (1'h0);
  reg [(3'h6):(1'h0)] reg4145 = (1'h0);
  reg [(3'h6):(1'h0)] reg4143 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4141 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4133 = (1'h0);
  reg [(3'h4):(1'h0)] reg4128 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4139 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4137 = (1'h0);
  reg [(4'he):(1'h0)] reg4136 = (1'h0);
  reg [(2'h2):(1'h0)] reg4135 = (1'h0);
  reg [(2'h3):(1'h0)] reg4134 = (1'h0);
  reg [(5'h10):(1'h0)] reg4132 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4131 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4130 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4129 = (1'h0);
  reg [(3'h4):(1'h0)] reg4127 = (1'h0);
  reg [(3'h7):(1'h0)] reg4125 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4100 = (1'h0);
  reg [(4'hf):(1'h0)] reg4108 = (1'h0);
  reg [(4'ha):(1'h0)] reg4104 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4103 = (1'h0);
  reg [(4'hd):(1'h0)] reg4097 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4124 = (1'h0);
  reg [(4'ha):(1'h0)] reg4123 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4122 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4120 = (1'h0);
  reg [(3'h6):(1'h0)] reg4119 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4118 = (1'h0);
  reg [(4'hd):(1'h0)] reg4117 = (1'h0);
  reg [(3'h4):(1'h0)] reg4116 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4109 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4115 = (1'h0);
  reg [(2'h3):(1'h0)] reg4114 = (1'h0);
  reg [(4'hb):(1'h0)] reg4113 = (1'h0);
  reg [(4'he):(1'h0)] reg4112 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4111 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4110 = (1'h0);
  reg [(4'h8):(1'h0)] reg4107 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4106 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4105 = (1'h0);
  reg [(2'h2):(1'h0)] reg4102 = (1'h0);
  reg [(5'h10):(1'h0)] reg4101 = (1'h0);
  reg [(4'h8):(1'h0)] reg4099 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4051 = (1'h0);
  reg [(2'h3):(1'h0)] reg4050 = (1'h0);
  reg [(3'h4):(1'h0)] reg4038 = (1'h0);
  reg [(4'h8):(1'h0)] reg4027 = (1'h0);
  reg [(4'h8):(1'h0)] reg4023 = (1'h0);
  reg [(3'h5):(1'h0)] reg4003 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4002 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3985 = (1'h0);
  reg [(4'hd):(1'h0)] reg3986 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3983 = (1'h0);
  reg [(4'h8):(1'h0)] reg3982 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3981 = (1'h0);
  reg [(3'h4):(1'h0)] reg4096 = (1'h0);
  reg [(3'h6):(1'h0)] reg4091 = (1'h0);
  reg [(4'h9):(1'h0)] reg4095 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4094 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4093 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4092 = (1'h0);
  reg [(4'h9):(1'h0)] reg4090 = (1'h0);
  reg [(4'hf):(1'h0)] reg4089 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4088 = (1'h0);
  reg [(4'hb):(1'h0)] reg4087 = (1'h0);
  reg [(4'hf):(1'h0)] reg4086 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4085 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4084 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4083 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4082 = (1'h0);
  reg [(5'h10):(1'h0)] reg4076 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4081 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4080 = (1'h0);
  reg [(3'h4):(1'h0)] reg4079 = (1'h0);
  reg [(3'h4):(1'h0)] reg4078 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4077 = (1'h0);
  reg [(4'he):(1'h0)] reg4075 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4074 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4073 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4071 = (1'h0);
  reg [(2'h2):(1'h0)] reg4070 = (1'h0);
  reg [(3'h4):(1'h0)] reg4069 = (1'h0);
  reg [(3'h5):(1'h0)] reg4068 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4067 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4066 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4065 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4064 = (1'h0);
  reg [(4'hd):(1'h0)] reg4063 = (1'h0);
  reg [(2'h3):(1'h0)] reg4062 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4061 = (1'h0);
  reg [(4'hd):(1'h0)] reg4060 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4059 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4058 = (1'h0);
  reg [(3'h6):(1'h0)] reg4057 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4056 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4055 = (1'h0);
  reg [(2'h2):(1'h0)] reg4054 = (1'h0);
  reg [(4'hc):(1'h0)] reg4053 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4052 = (1'h0);
  reg [(3'h6):(1'h0)] reg4049 = (1'h0);
  reg [(4'hc):(1'h0)] reg4048 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4044 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4040 = (1'h0);
  reg [(3'h4):(1'h0)] reg4047 = (1'h0);
  reg [(3'h7):(1'h0)] reg4046 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4045 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4043 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4042 = (1'h0);
  reg [(5'h10):(1'h0)] reg4041 = (1'h0);
  reg [(4'ha):(1'h0)] reg4039 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4037 = (1'h0);
  reg [(4'he):(1'h0)] reg4034 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4031 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4036 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4035 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4033 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4032 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4030 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4029 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4028 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4015 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4026 = (1'h0);
  reg [(4'hf):(1'h0)] reg4025 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4024 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4022 = (1'h0);
  reg [(2'h3):(1'h0)] reg4021 = (1'h0);
  reg [(3'h4):(1'h0)] reg4019 = (1'h0);
  reg [(4'hf):(1'h0)] reg4018 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4016 = (1'h0);
  reg [(5'h10):(1'h0)] reg4014 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4012 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4011 = (1'h0);
  reg [(4'h9):(1'h0)] reg4010 = (1'h0);
  reg [(4'hb):(1'h0)] reg4009 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4008 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4007 = (1'h0);
  reg [(2'h2):(1'h0)] reg4006 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4004 = (1'h0);
  reg [(4'h8):(1'h0)] reg4001 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4000 = (1'h0);
  reg [(5'h10):(1'h0)] reg3999 = (1'h0);
  reg [(5'h10):(1'h0)] reg3998 = (1'h0);
  reg [(2'h2):(1'h0)] reg3997 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3996 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3995 = (1'h0);
  reg [(2'h3):(1'h0)] reg3994 = (1'h0);
  reg [(2'h2):(1'h0)] reg3992 = (1'h0);
  reg [(4'ha):(1'h0)] reg3991 = (1'h0);
  reg [(5'h10):(1'h0)] reg3990 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3989 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3988 = (1'h0);
  reg [(5'h10):(1'h0)] reg3987 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3984 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3980 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3979 = (1'h0);
  reg [(4'hd):(1'h0)] reg3978 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3977 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3976 = (1'h0);
  reg [(4'hc):(1'h0)] reg3975 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3974 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3973 = (1'h0);
  reg [(4'ha):(1'h0)] reg3971 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3970 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3969 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3968 = (1'h0);
  reg [(2'h2):(1'h0)] reg3966 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3965 = (1'h0);
  reg [(5'h10):(1'h0)] reg3964 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3963 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3961 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3960 = (1'h0);
  reg [(4'h8):(1'h0)] reg3958 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3957 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3956 = (1'h0);
  reg [(3'h7):(1'h0)] reg3952 = (1'h0);
  reg [(4'h8):(1'h0)] reg3949 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3955 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3954 = (1'h0);
  reg [(2'h2):(1'h0)] reg3953 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3951 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3950 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3948 = (1'h0);
  reg [(2'h2):(1'h0)] reg3947 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3946 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3945 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4209 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4204 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4205 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4201 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4197 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4194 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4192 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4160 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4152 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4186 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4179 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4173 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4171 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4170 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4168 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4157 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4158 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4153 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4148 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4144 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4142 = (1'h0);
  reg [(4'he):(1'h0)] forvar4140 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4135 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4134 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4129 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4127 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4138 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4133 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4128 = (1'h0);
  reg [(4'he):(1'h0)] forvar4126 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4107 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4102 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4121 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4109 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4108 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4104 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4103 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4100 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4098 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4097 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4058 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4075 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4069 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4060 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4059 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4054 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4047 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4046 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4037 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4036 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4029 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4024 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4004 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4091 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4078 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4071 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4076 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4072 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4051 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4050 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4044 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4040 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4038 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4035 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4033 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4028 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4034 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4031 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4027 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4023 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4020 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4017 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4015 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4013 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4005 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4003 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4002 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3993 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3986 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3985 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3983 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3982 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3981 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3968 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3975 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3972 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3967 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3948 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3962 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3959 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3954 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3950 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3952 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3949 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3945 = (1'h0);
  assign y = {wire4538,
                 wire4537,
                 wire4536,
                 wire4535,
                 wire4533,
                 wire4213,
                 wire4212,
                 wire3944,
                 wire3943,
                 wire3942,
                 reg4126,
                 reg4211,
                 reg4210,
                 reg4208,
                 reg4207,
                 reg4205,
                 reg4206,
                 reg4204,
                 reg4203,
                 reg4202,
                 reg4200,
                 reg4199,
                 reg4198,
                 reg4194,
                 reg4196,
                 reg4195,
                 reg4193,
                 reg4153,
                 reg4148,
                 reg4191,
                 reg4190,
                 reg4189,
                 reg4188,
                 reg4187,
                 reg4185,
                 reg4184,
                 reg4183,
                 reg4182,
                 reg4181,
                 reg4180,
                 reg4178,
                 reg4177,
                 reg4176,
                 reg4175,
                 reg4174,
                 reg4172,
                 reg4169,
                 reg4167,
                 reg4166,
                 reg4165,
                 reg4164,
                 reg4158,
                 reg4163,
                 reg4162,
                 reg4161,
                 reg4160,
                 reg4159,
                 reg4157,
                 reg4156,
                 reg4155,
                 reg4154,
                 reg4152,
                 reg4151,
                 reg4150,
                 reg4149,
                 reg4147,
                 reg4144,
                 reg4146,
                 reg4145,
                 reg4143,
                 reg4141,
                 reg4133,
                 reg4128,
                 reg4139,
                 reg4137,
                 reg4136,
                 reg4135,
                 reg4134,
                 reg4132,
                 reg4131,
                 reg4130,
                 reg4129,
                 reg4127,
                 reg4125,
                 reg4100,
                 reg4108,
                 reg4104,
                 reg4103,
                 reg4097,
                 reg4124,
                 reg4123,
                 reg4122,
                 reg4120,
                 reg4119,
                 reg4118,
                 reg4117,
                 reg4116,
                 reg4109,
                 reg4115,
                 reg4114,
                 reg4113,
                 reg4112,
                 reg4111,
                 reg4110,
                 reg4107,
                 reg4106,
                 reg4105,
                 reg4102,
                 reg4101,
                 reg4099,
                 reg4051,
                 reg4050,
                 reg4038,
                 reg4027,
                 reg4023,
                 reg4003,
                 reg4002,
                 reg3985,
                 reg3986,
                 reg3983,
                 reg3982,
                 reg3981,
                 reg4096,
                 reg4091,
                 reg4095,
                 reg4094,
                 reg4093,
                 reg4092,
                 reg4090,
                 reg4089,
                 reg4088,
                 reg4087,
                 reg4086,
                 reg4085,
                 reg4084,
                 reg4083,
                 reg4082,
                 reg4076,
                 reg4081,
                 reg4080,
                 reg4079,
                 reg4078,
                 reg4077,
                 reg4075,
                 reg4074,
                 reg4073,
                 reg4071,
                 reg4070,
                 reg4069,
                 reg4068,
                 reg4067,
                 reg4066,
                 reg4065,
                 reg4064,
                 reg4063,
                 reg4062,
                 reg4061,
                 reg4060,
                 reg4059,
                 reg4058,
                 reg4057,
                 reg4056,
                 reg4055,
                 reg4054,
                 reg4053,
                 reg4052,
                 reg4049,
                 reg4048,
                 reg4044,
                 reg4040,
                 reg4047,
                 reg4046,
                 reg4045,
                 reg4043,
                 reg4042,
                 reg4041,
                 reg4039,
                 reg4037,
                 reg4034,
                 reg4031,
                 reg4036,
                 reg4035,
                 reg4033,
                 reg4032,
                 reg4030,
                 reg4029,
                 reg4028,
                 reg4015,
                 reg4026,
                 reg4025,
                 reg4024,
                 reg4022,
                 reg4021,
                 reg4019,
                 reg4018,
                 reg4016,
                 reg4014,
                 reg4012,
                 reg4011,
                 reg4010,
                 reg4009,
                 reg4008,
                 reg4007,
                 reg4006,
                 reg4004,
                 reg4001,
                 reg4000,
                 reg3999,
                 reg3998,
                 reg3997,
                 reg3996,
                 reg3995,
                 reg3994,
                 reg3992,
                 reg3991,
                 reg3990,
                 reg3989,
                 reg3988,
                 reg3987,
                 reg3984,
                 reg3980,
                 reg3979,
                 reg3978,
                 reg3977,
                 reg3976,
                 reg3975,
                 reg3974,
                 reg3973,
                 reg3971,
                 reg3970,
                 reg3969,
                 reg3968,
                 reg3966,
                 reg3965,
                 reg3964,
                 reg3963,
                 reg3961,
                 reg3960,
                 reg3958,
                 reg3957,
                 reg3956,
                 reg3952,
                 reg3949,
                 reg3955,
                 reg3954,
                 reg3953,
                 reg3951,
                 reg3950,
                 reg3948,
                 reg3947,
                 reg3946,
                 reg3945,
                 forvar4209,
                 forvar4204,
                 forvar4205,
                 forvar4201,
                 forvar4197,
                 forvar4194,
                 forvar4192,
                 forvar4160,
                 forvar4152,
                 forvar4186,
                 forvar4179,
                 forvar4173,
                 forvar4171,
                 forvar4170,
                 forvar4168,
                 forvar4157,
                 forvar4158,
                 forvar4153,
                 forvar4148,
                 forvar4144,
                 forvar4142,
                 forvar4140,
                 forvar4135,
                 forvar4134,
                 forvar4129,
                 forvar4127,
                 forvar4138,
                 forvar4133,
                 forvar4128,
                 forvar4126,
                 forvar4107,
                 forvar4102,
                 forvar4121,
                 forvar4109,
                 forvar4108,
                 forvar4104,
                 forvar4103,
                 forvar4100,
                 forvar4098,
                 forvar4097,
                 forvar4058,
                 forvar4075,
                 forvar4069,
                 forvar4060,
                 forvar4059,
                 forvar4054,
                 forvar4047,
                 forvar4046,
                 forvar4037,
                 forvar4036,
                 forvar4029,
                 forvar4024,
                 forvar4004,
                 forvar4091,
                 forvar4078,
                 forvar4071,
                 forvar4076,
                 forvar4072,
                 forvar4051,
                 forvar4050,
                 forvar4044,
                 forvar4040,
                 forvar4038,
                 forvar4035,
                 forvar4033,
                 forvar4028,
                 forvar4034,
                 forvar4031,
                 forvar4027,
                 forvar4023,
                 forvar4020,
                 forvar4017,
                 forvar4015,
                 forvar4013,
                 forvar4005,
                 forvar4003,
                 forvar4002,
                 forvar3993,
                 forvar3986,
                 forvar3985,
                 forvar3983,
                 forvar3982,
                 forvar3981,
                 forvar3968,
                 forvar3975,
                 forvar3972,
                 forvar3967,
                 forvar3948,
                 forvar3962,
                 forvar3959,
                 forvar3954,
                 forvar3950,
                 forvar3952,
                 forvar3949,
                 forvar3945,
                 (1'h0)};
  assign wire3942 = (~&((8'haf) ?
                        ((^~(8'h9d)) | wire3937) : ((wire3940 ?
                                wire3941 : wire3938) ?
                            $signed((8'hb5)) : $unsigned((8'ha8)))));
  assign wire3943 = $unsigned(wire3940);
  assign wire3944 = ($signed($signed(((8'ha4) ?
                        (8'had) : wire3942))) <= wire3937[(2'h2):(1'h1)]);
  always
    @(posedge clk) begin
      if (((~wire3944[(2'h3):(2'h3)]) <<< wire3944))
        begin
          if ((^$signed(((wire3944 ? wire3943 : wire3940) ?
              (wire3937 << (8'hb9)) : wire3944[(2'h2):(2'h2)]))))
            begin
              if ((!{$signed(wire3942)}))
                begin
                  reg3945 <= (wire3939[(3'h4):(1'h0)] << wire3938);
                end
              else
                begin
                  for (forvar3945 = (1'h0); (forvar3945 < (2'h2)); forvar3945 = (forvar3945 + (1'h1)))
                    begin
                      reg3946 <= reg3945;
                      reg3947 <= $unsigned(wire3943);
                    end
                  reg3948 <= reg3947[(1'h1):(1'h1)];
                end
              for (forvar3949 = (1'h0); (forvar3949 < (1'h1)); forvar3949 = (forvar3949 + (1'h1)))
                begin
                  reg3950 <= (8'ha7);
                  reg3951 <= $signed(wire3941);
                end
              for (forvar3952 = (1'h0); (forvar3952 < (1'h1)); forvar3952 = (forvar3952 + (1'h1)))
                begin
                  if (($signed(reg3948) ?
                      ((8'ha1) ?
                          (wire3939 || (-forvar3952)) : ((reg3945 ?
                                  forvar3945 : (8'haf)) ?
                              wire3940 : $signed(wire3941))) : $unsigned($signed(forvar3945[(2'h2):(2'h2)]))))
                    begin
                      reg3953 <= (8'ha3);
                    end
                  else
                    begin
                      reg3953 <= reg3946[(3'h4):(2'h3)];
                      reg3954 <= $unsigned(($signed($unsigned(wire3937)) ?
                          reg3953[(1'h1):(1'h1)] : (!$unsigned(reg3950))));
                      reg3955 <= $unsigned(wire3941[(3'h7):(2'h3)]);
                    end
                end
            end
          else
            begin
              for (forvar3945 = (1'h0); (forvar3945 < (2'h2)); forvar3945 = (forvar3945 + (1'h1)))
                begin
                  if ({((wire3938[(3'h4):(3'h4)] ?
                          (reg3955 == wire3942) : (^~wire3944)) != $signed((wire3942 ?
                          forvar3952 : reg3953)))})
                    begin
                      reg3946 <= $signed((^wire3937));
                      reg3947 <= wire3943[(3'h4):(3'h4)];
                      reg3948 <= {wire3939};
                      reg3949 <= $signed((((wire3937 ?
                              reg3950 : (8'h9d)) && ((8'h9c) ?
                              forvar3952 : wire3941)) ?
                          (reg3951 < reg3955) : (!$signed(wire3939))));
                    end
                  else
                    begin
                      reg3946 <= ((|$signed((reg3949 - wire3941))) != (reg3953[(1'h1):(1'h0)] ?
                          ((reg3951 || (8'h9f)) ?
                              reg3947[(2'h2):(2'h2)] : (wire3944 >>> wire3942)) : ($signed(reg3953) == (forvar3949 & reg3949))));
                      reg3947 <= (wire3938[(1'h0):(1'h0)] != {((~wire3937) ?
                              (reg3949 ? reg3954 : (8'hb6)) : wire3940)});
                    end
                end
            end
        end
      else
        begin
          if ((~(forvar3952[(3'h7):(2'h2)] || reg3946)))
            begin
              if ({{wire3939[(2'h2):(2'h2)]}})
                begin
                  reg3945 <= ((^forvar3945[(3'h4):(1'h1)]) ?
                      (~(-$unsigned((8'hac)))) : wire3943[(1'h1):(1'h1)]);
                end
              else
                begin
                  for (forvar3945 = (1'h0); (forvar3945 < (1'h1)); forvar3945 = (forvar3945 + (1'h1)))
                    begin
                      reg3946 <= $unsigned($signed(($signed(forvar3945) + $unsigned(wire3940))));
                      reg3947 <= ({reg3945} < ((reg3949 < wire3939[(1'h1):(1'h0)]) || $signed((~|reg3949))));
                      reg3948 <= wire3944;
                      reg3949 <= $signed($signed(reg3946[(3'h4):(1'h1)]));
                    end
                  for (forvar3950 = (1'h0); (forvar3950 < (1'h0)); forvar3950 = (forvar3950 + (1'h1)))
                    begin
                      reg3951 <= (-(reg3950[(2'h3):(1'h1)] << ((wire3937 ?
                          reg3949 : forvar3952) * (|forvar3949))));
                      reg3952 <= $signed(($signed((&wire3944)) ^ {reg3949}));
                      reg3953 <= $signed(wire3941[(4'hc):(4'h9)]);
                    end
                  for (forvar3954 = (1'h0); (forvar3954 < (2'h2)); forvar3954 = (forvar3954 + (1'h1)))
                    begin
                      reg3955 <= wire3939;
                      reg3956 <= (8'ha0);
                      reg3957 <= $unsigned((&(|{forvar3949})));
                      reg3958 <= (~(reg3946 == $unsigned($unsigned(reg3953))));
                    end
                  for (forvar3959 = (1'h0); (forvar3959 < (2'h2)); forvar3959 = (forvar3959 + (1'h1)))
                    begin
                      reg3960 <= forvar3954;
                      reg3961 <= ($unsigned($signed({forvar3952})) | (forvar3949 ?
                          reg3949[(3'h5):(3'h4)] : $signed((|(8'hac)))));
                    end
                end
              for (forvar3962 = (1'h0); (forvar3962 < (1'h0)); forvar3962 = (forvar3962 + (1'h1)))
                begin
                  if ($unsigned($signed((~reg3957))))
                    begin
                      reg3963 <= (({$unsigned(reg3949)} || reg3951[(2'h2):(1'h1)]) <= (((8'haa) << (wire3943 >> reg3958)) ^ $signed((^~wire3943))));
                      reg3964 <= $signed(forvar3949[(3'h7):(2'h3)]);
                      reg3965 <= {(wire3940[(1'h0):(1'h0)] & {{reg3961}})};
                      reg3966 <= forvar3945[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3963 <= {$unsigned(($unsigned(wire3942) ~^ (reg3949 ^~ reg3961)))};
                    end
                end
            end
          else
            begin
              for (forvar3945 = (1'h0); (forvar3945 < (1'h1)); forvar3945 = (forvar3945 + (1'h1)))
                begin
                  if ($signed((reg3966[(1'h1):(1'h0)] ?
                      $signed((&reg3957)) : $unsigned((~^(8'had))))))
                    begin
                      reg3946 <= ((((reg3946 ?
                              wire3942 : reg3953) + (8'hb9)) >>> (^~wire3944[(3'h4):(1'h1)])) ?
                          reg3966 : $unsigned(wire3939));
                    end
                  else
                    begin
                      reg3946 <= (^~$signed({$unsigned(reg3945)}));
                      reg3947 <= wire3944;
                    end
                end
              for (forvar3948 = (1'h0); (forvar3948 < (2'h3)); forvar3948 = (forvar3948 + (1'h1)))
                begin
                  for (forvar3949 = (1'h0); (forvar3949 < (2'h3)); forvar3949 = (forvar3949 + (1'h1)))
                    begin
                      reg3950 <= $signed($unsigned(((reg3950 ?
                              reg3954 : reg3958) ?
                          ((8'ha7) ? forvar3959 : forvar3950) : (~|wire3940))));
                      reg3951 <= wire3940;
                      reg3952 <= ($signed(reg3955) < reg3952);
                    end
                  if (((~^reg3953[(1'h1):(1'h0)]) ?
                      ($unsigned((wire3938 ?
                          (8'ha0) : reg3958)) ^~ {(~^forvar3945)}) : ({(reg3953 ?
                              (8'ha5) : reg3961)} && wire3937)))
                    begin
                      reg3953 <= wire3943;
                    end
                  else
                    begin
                      reg3953 <= ((((reg3960 ?
                              forvar3952 : reg3964) >> (reg3955 >= (8'hb4))) ~^ $unsigned(reg3966)) ?
                          (reg3946[(1'h1):(1'h1)] ?
                              $signed({wire3943}) : $unsigned($unsigned(wire3941))) : ((((8'hae) > reg3957) << (^~reg3956)) ?
                              $signed(((8'hb0) ^ reg3958)) : $unsigned(reg3963[(1'h0):(1'h0)])));
                      reg3954 <= $unsigned(({$signed(wire3943)} ?
                          (8'ha1) : reg3965[(3'h5):(1'h0)]));
                      reg3955 <= reg3951;
                      reg3956 <= (forvar3950 ?
                          wire3943[(2'h3):(2'h3)] : $unsigned(reg3960));
                    end
                end
            end
          if ((wire3937 ?
              (-$unsigned((forvar3959 || forvar3962))) : {$signed((forvar3948 || reg3950))}))
            begin
              if (($unsigned($unsigned((8'ha9))) ~^ (($unsigned(reg3960) ?
                  $unsigned(reg3966) : (8'hae)) && {$signed(forvar3959)})))
                begin
                  for (forvar3967 = (1'h0); (forvar3967 < (1'h0)); forvar3967 = (forvar3967 + (1'h1)))
                    begin
                      reg3968 <= forvar3945[(2'h2):(1'h0)];
                      reg3969 <= $unsigned((-reg3960[(2'h3):(2'h2)]));
                    end
                end
              else
                begin
                  for (forvar3967 = (1'h0); (forvar3967 < (1'h1)); forvar3967 = (forvar3967 + (1'h1)))
                    begin
                      reg3968 <= $signed(((+forvar3945) > $unsigned({reg3969})));
                      reg3969 <= $signed(forvar3967[(1'h0):(1'h0)]);
                      reg3970 <= ((wire3937 ?
                              ((reg3965 ?
                                  forvar3949 : wire3938) & (-forvar3954)) : {reg3963[(1'h1):(1'h1)]}) ?
                          $unsigned(reg3954[(3'h5):(2'h3)]) : (-forvar3967[(1'h0):(1'h0)]));
                      reg3971 <= $signed((~&((+reg3955) <= $unsigned(reg3969))));
                    end
                  for (forvar3972 = (1'h0); (forvar3972 < (1'h0)); forvar3972 = (forvar3972 + (1'h1)))
                    begin
                      reg3973 <= (|reg3969[(3'h4):(2'h2)]);
                      reg3974 <= forvar3950;
                    end
                end
              if (forvar3967)
                begin
                  if (reg3952)
                    begin
                      reg3975 <= reg3961[(3'h7):(2'h3)];
                      reg3976 <= $unsigned(((~|reg3958[(4'h8):(4'h8)]) ?
                          (&{wire3938}) : reg3968));
                      reg3977 <= reg3953[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg3975 <= $unsigned((!reg3975));
                      reg3976 <= {reg3956[(3'h6):(2'h2)]};
                      reg3977 <= ((^~(^~reg3960)) ^ $signed(reg3971));
                      reg3978 <= (($unsigned((reg3953 ? forvar3954 : reg3956)) ?
                              ($unsigned(reg3973) < reg3964[(5'h10):(3'h7)]) : (+(^~reg3949))) ?
                          forvar3948[(3'h4):(1'h1)] : forvar3972);
                    end
                  if (wire3939)
                    begin
                      reg3979 <= ((((^reg3955) ? (~|forvar3950) : (~(8'hb3))) ?
                          $unsigned(((8'h9f) ?
                              reg3957 : wire3938)) : {(8'h9c)}) >= (reg3976 ?
                          {$signed(wire3944)} : ((wire3940 + forvar3948) << (reg3973 * reg3973))));
                      reg3980 <= reg3960[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3979 <= forvar3954[(3'h7):(3'h6)];
                    end
                end
              else
                begin
                  for (forvar3975 = (1'h0); (forvar3975 < (1'h1)); forvar3975 = (forvar3975 + (1'h1)))
                    begin
                      reg3976 <= wire3941[(1'h0):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar3967 = (1'h0); (forvar3967 < (2'h3)); forvar3967 = (forvar3967 + (1'h1)))
                begin
                  for (forvar3968 = (1'h0); (forvar3968 < (2'h2)); forvar3968 = (forvar3968 + (1'h1)))
                    begin
                      reg3969 <= (((~^reg3977) ?
                              forvar3968 : reg3958[(3'h6):(2'h2)]) ?
                          ($signed($signed(reg3949)) - reg3957[(1'h1):(1'h1)]) : (!$unsigned((forvar3954 - (8'hb2)))));
                      reg3970 <= (~^reg3966[(2'h2):(1'h1)]);
                      reg3971 <= forvar3954[(3'h7):(3'h5)];
                    end
                  for (forvar3972 = (1'h0); (forvar3972 < (2'h2)); forvar3972 = (forvar3972 + (1'h1)))
                    begin
                      reg3973 <= (&(({reg3975} ?
                          (reg3977 ?
                              forvar3945 : reg3955) : $signed(wire3937)) * forvar3949[(3'h5):(2'h2)]));
                    end
                  if ((forvar3950[(3'h7):(1'h1)] ?
                      $signed(($signed((8'ha5)) ~^ (&reg3947))) : (reg3945[(3'h4):(3'h4)] + (~&(reg3961 ~^ wire3943)))))
                    begin
                      reg3974 <= (((~&$signed(wire3943)) ?
                              ({(8'h9f)} <<< $signed(reg3979)) : $unsigned($unsigned(reg3966))) ?
                          $signed({reg3949}) : {(reg3980 ?
                                  (forvar3967 ?
                                      reg3947 : (8'ha5)) : $unsigned(reg3953))});
                    end
                  else
                    begin
                      reg3974 <= reg3945[(2'h3):(1'h0)];
                      reg3975 <= reg3947[(1'h0):(1'h0)];
                      reg3976 <= forvar3967[(2'h3):(1'h1)];
                      reg3977 <= ($signed(({wire3937} >> reg3945[(4'h8):(3'h6)])) ?
                          (~|((^~reg3963) ?
                              (+reg3979) : (8'haf))) : forvar3975);
                    end
                end
              reg3978 <= ($signed(((reg3966 ? wire3944 : reg3964) ?
                  (8'hb5) : reg3977)) << (+reg3968[(4'h9):(1'h1)]));
            end
        end
      if ($signed($unsigned({(forvar3945 * reg3975)})))
        begin
          for (forvar3981 = (1'h0); (forvar3981 < (1'h1)); forvar3981 = (forvar3981 + (1'h1)))
            begin
              for (forvar3982 = (1'h0); (forvar3982 < (2'h3)); forvar3982 = (forvar3982 + (1'h1)))
                begin
                  for (forvar3983 = (1'h0); (forvar3983 < (1'h0)); forvar3983 = (forvar3983 + (1'h1)))
                    begin
                      reg3984 <= $unsigned(((reg3963[(1'h1):(1'h0)] ?
                          reg3976 : forvar3952[(2'h2):(2'h2)]) > (|reg3973[(3'h4):(1'h1)])));
                    end
                end
              for (forvar3985 = (1'h0); (forvar3985 < (1'h1)); forvar3985 = (forvar3985 + (1'h1)))
                begin
                  for (forvar3986 = (1'h0); (forvar3986 < (1'h0)); forvar3986 = (forvar3986 + (1'h1)))
                    begin
                      reg3987 <= ($signed($signed($unsigned(forvar3968))) <= {$unsigned((-reg3953))});
                      reg3988 <= $unsigned(reg3973);
                      reg3989 <= forvar3945[(3'h6):(1'h0)];
                      reg3990 <= wire3937;
                    end
                  if ($signed(reg3946))
                    begin
                      reg3991 <= $unsigned(forvar3945);
                      reg3992 <= ((~&((reg3971 ?
                              (8'h9e) : reg3976) && $signed(reg3977))) ?
                          $unsigned(($unsigned(reg3957) ^~ (~&(8'h9f)))) : (reg3951[(3'h5):(2'h3)] ?
                              $unsigned($unsigned(forvar3972)) : reg3976[(3'h5):(2'h2)]));
                    end
                  else
                    begin
                      reg3991 <= ({forvar3985} <= reg3946[(3'h5):(1'h0)]);
                    end
                  for (forvar3993 = (1'h0); (forvar3993 < (1'h1)); forvar3993 = (forvar3993 + (1'h1)))
                    begin
                      reg3994 <= ($unsigned($signed(reg3991[(4'h8):(3'h6)])) ?
                          reg3980 : reg3977[(3'h7):(1'h0)]);
                      reg3995 <= $signed(((^forvar3986) >= (reg3950 ?
                          $unsigned(reg3984) : reg3984[(3'h4):(3'h4)])));
                      reg3996 <= $unsigned((^({(8'hb1)} << $signed((8'hac)))));
                      reg3997 <= (+{(~|{(8'h9e)})});
                    end
                  if (reg3960[(2'h3):(1'h0)])
                    begin
                      reg3998 <= (($unsigned((reg3947 && reg3964)) >>> (((8'hb0) ?
                                  (8'ha0) : reg3976) ?
                              (forvar3985 <= forvar3985) : forvar3972)) ?
                          $unsigned(reg3956) : $unsigned((|$unsigned(reg3951))));
                      reg3999 <= $unsigned(((reg3951 ?
                              (reg3964 != (8'hb5)) : (8'hac)) ?
                          $signed((~^forvar3975)) : forvar3954));
                      reg4000 <= reg3977;
                      reg4001 <= ((reg3984 ?
                          $signed({reg3973}) : forvar3945[(3'h7):(2'h2)]) - (~^($unsigned((8'had)) & (forvar3986 ?
                          reg3968 : (8'ha4)))));
                    end
                  else
                    begin
                      reg3998 <= forvar3950[(1'h1):(1'h0)];
                      reg3999 <= $unsigned(reg3948);
                      reg4000 <= $signed($signed((reg3992 ?
                          forvar3986 : $unsigned(reg3955))));
                      reg4001 <= wire3944[(2'h3):(2'h3)];
                    end
                end
              for (forvar4002 = (1'h0); (forvar4002 < (2'h3)); forvar4002 = (forvar4002 + (1'h1)))
                begin
                  for (forvar4003 = (1'h0); (forvar4003 < (1'h0)); forvar4003 = (forvar4003 + (1'h1)))
                    begin
                      reg4004 <= $unsigned(reg3992);
                    end
                  for (forvar4005 = (1'h0); (forvar4005 < (1'h1)); forvar4005 = (forvar4005 + (1'h1)))
                    begin
                      reg4006 <= (reg3946 ?
                          (!reg3951) : ((wire3938[(1'h0):(1'h0)] ?
                                  (&forvar3986) : forvar3948) ?
                              (~|$signed(reg3961)) : ((reg3971 ?
                                  reg3950 : wire3939) <<< reg3971)));
                    end
                end
              if ((forvar4005 ?
                  reg3958 : $unsigned($signed((reg3957 ? reg4004 : reg3978)))))
                begin
                  reg4007 <= reg3990[(4'hb):(3'h7)];
                end
              else
                begin
                  if ($signed(reg3995))
                    begin
                      reg4007 <= reg3963;
                      reg4008 <= $signed(forvar3993);
                      reg4009 <= {{{(!(8'h9c))}}};
                    end
                  else
                    begin
                      reg4007 <= reg4008[(3'h7):(3'h6)];
                      reg4008 <= reg3987[(3'h7):(3'h4)];
                      reg4009 <= (^~(reg3961[(4'h8):(1'h0)] ?
                          (reg3988 * (forvar4003 ?
                              reg3953 : reg3976)) : {(8'ha7)}));
                      reg4010 <= ((((~|reg3989) ?
                              reg3964 : $unsigned(forvar3986)) ?
                          reg3963 : $signed((^~reg3948))) + ($unsigned($signed((8'ha3))) * ($unsigned(reg3995) ?
                          forvar3968 : $signed(forvar3983))));
                    end
                  reg4011 <= (+(^~reg3991));
                  if ((8'hae))
                    begin
                      reg4012 <= $signed((&forvar3962[(2'h3):(1'h1)]));
                    end
                  else
                    begin
                      reg4012 <= (8'hb7);
                    end
                  for (forvar4013 = (1'h0); (forvar4013 < (2'h2)); forvar4013 = (forvar4013 + (1'h1)))
                    begin
                      reg4014 <= (reg3956[(3'h4):(3'h4)] ?
                          (($unsigned(reg4007) & reg3957) ?
                              (8'ha7) : ((reg3989 ? reg3977 : reg3954) ?
                                  reg3963 : (wire3937 <<< reg3980))) : ({$signed(forvar4002)} + $unsigned($unsigned((8'ha0)))));
                    end
                end
            end
          if (({$signed($signed(forvar3949))} ^~ ((-$signed(reg3995)) ?
              $unsigned($unsigned((8'had))) : ((!reg4007) ^~ (^~(8'h9e))))))
            begin
              for (forvar4015 = (1'h0); (forvar4015 < (1'h0)); forvar4015 = (forvar4015 + (1'h1)))
                begin
                  reg4016 <= reg3950;
                end
              for (forvar4017 = (1'h0); (forvar4017 < (2'h2)); forvar4017 = (forvar4017 + (1'h1)))
                begin
                  if ((((((8'h9f) ? reg3958 : reg3969) ?
                      $signed(reg3961) : $unsigned((8'hb5))) < $unsigned($unsigned(reg3969))) < reg3949))
                    begin
                      reg4018 <= reg3964[(4'hd):(3'h6)];
                      reg4019 <= $unsigned(($signed((forvar3954 ?
                              forvar3967 : reg3966)) ?
                          (forvar4002 >> $signed(forvar3945)) : (8'haf)));
                    end
                  else
                    begin
                      reg4018 <= (reg3970 - (8'h9e));
                    end
                end
              for (forvar4020 = (1'h0); (forvar4020 < (1'h1)); forvar4020 = (forvar4020 + (1'h1)))
                begin
                  reg4021 <= forvar3954[(2'h2):(1'h1)];
                  reg4022 <= reg3965;
                  for (forvar4023 = (1'h0); (forvar4023 < (1'h0)); forvar4023 = (forvar4023 + (1'h1)))
                    begin
                      reg4024 <= $signed({{(!reg4016)}});
                    end
                  if (reg3951[(3'h4):(1'h0)])
                    begin
                      reg4025 <= (~|$signed($signed((reg4016 <= reg3963))));
                    end
                  else
                    begin
                      reg4025 <= (reg4024[(2'h2):(2'h2)] ?
                          forvar3950[(3'h6):(1'h0)] : (-(&(forvar4013 ?
                              forvar3981 : (8'ha1)))));
                      reg4026 <= reg3994;
                    end
                end
            end
          else
            begin
              reg4015 <= reg3990;
            end
          for (forvar4027 = (1'h0); (forvar4027 < (2'h3)); forvar4027 = (forvar4027 + (1'h1)))
            begin
              if ((^~reg4026))
                begin
                  if ($signed(reg3999[(3'h5):(1'h1)]))
                    begin
                      reg4028 <= reg3996;
                    end
                  else
                    begin
                      reg4028 <= ($unsigned($unsigned($unsigned(wire3941))) ?
                          $unsigned($signed($signed(forvar3945))) : (~({forvar4017} ?
                              reg4011 : forvar3986[(2'h2):(1'h1)])));
                      reg4029 <= (8'hac);
                      reg4030 <= forvar3968;
                    end
                  for (forvar4031 = (1'h0); (forvar4031 < (2'h2)); forvar4031 = (forvar4031 + (1'h1)))
                    begin
                      reg4032 <= (({forvar3967} ?
                          (reg4029[(4'h8):(3'h4)] >>> (~|reg3976)) : ($unsigned(forvar4013) ?
                              forvar3982 : (forvar3950 || reg3989))) << $unsigned(forvar3986[(2'h3):(1'h1)]));
                      reg4033 <= reg3978[(4'ha):(1'h1)];
                    end
                  for (forvar4034 = (1'h0); (forvar4034 < (1'h1)); forvar4034 = (forvar4034 + (1'h1)))
                    begin
                      reg4035 <= $unsigned(({(~&reg4016)} ^ ((^reg3989) ~^ forvar4013[(4'ha):(4'h9)])));
                      reg4036 <= ((&$unsigned($unsigned(reg4015))) ?
                          ($signed(reg3966[(2'h2):(1'h1)]) ?
                              (-$unsigned(forvar3962)) : ($unsigned((8'h9f)) ?
                                  (8'hb4) : (~reg4006))) : wire3937);
                    end
                end
              else
                begin
                  for (forvar4028 = (1'h0); (forvar4028 < (1'h1)); forvar4028 = (forvar4028 + (1'h1)))
                    begin
                      reg4029 <= (wire3940 ~^ (reg3956[(3'h4):(3'h4)] > {$signed(reg4019)}));
                      reg4030 <= forvar3975;
                      reg4031 <= $signed($unsigned((8'hb0)));
                      reg4032 <= (forvar3981 ?
                          ((^$unsigned((8'ha4))) ?
                              (~|(reg3958 ?
                                  reg3992 : (8'ha5))) : reg4006) : (&{reg3958[(1'h1):(1'h0)]}));
                    end
                  for (forvar4033 = (1'h0); (forvar4033 < (1'h1)); forvar4033 = (forvar4033 + (1'h1)))
                    begin
                      reg4034 <= (!$unsigned($unsigned((8'ha1))));
                    end
                  for (forvar4035 = (1'h0); (forvar4035 < (2'h3)); forvar4035 = (forvar4035 + (1'h1)))
                    begin
                      reg4036 <= $signed(reg3980);
                      reg4037 <= (8'ha5);
                    end
                  for (forvar4038 = (1'h0); (forvar4038 < (2'h3)); forvar4038 = (forvar4038 + (1'h1)))
                    begin
                      reg4039 <= (+reg3976);
                    end
                end
              if ((~&$unsigned(reg3997[(1'h0):(1'h0)])))
                begin
                  for (forvar4040 = (1'h0); (forvar4040 < (1'h0)); forvar4040 = (forvar4040 + (1'h1)))
                    begin
                      reg4041 <= $unsigned($unsigned($unsigned(wire3940[(1'h0):(1'h0)])));
                      reg4042 <= $unsigned((^($signed(forvar4023) - forvar3967[(1'h1):(1'h1)])));
                    end
                  reg4043 <= forvar4003;
                  for (forvar4044 = (1'h0); (forvar4044 < (1'h0)); forvar4044 = (forvar4044 + (1'h1)))
                    begin
                      reg4045 <= $unsigned((~&(reg4031 - $unsigned((8'ha8)))));
                    end
                  if (reg4045[(1'h0):(1'h0)])
                    begin
                      reg4046 <= (!(!$unsigned((wire3943 || reg3990))));
                      reg4047 <= $signed(((^~reg4039[(2'h3):(1'h1)]) && ((&reg3945) >= (reg3969 >>> reg3994))));
                    end
                  else
                    begin
                      reg4046 <= (-(~^((forvar3967 == reg4010) <= ((8'hb5) ?
                          reg3961 : reg3960))));
                    end
                end
              else
                begin
                  if ($signed($signed(reg3960[(3'h4):(2'h3)])))
                    begin
                      reg4040 <= $signed($unsigned($unsigned($unsigned((8'hb8)))));
                      reg4041 <= ($signed(reg4001) << {(|(forvar3952 > (8'hb4)))});
                      reg4042 <= $unsigned(reg3975);
                    end
                  else
                    begin
                      reg4040 <= ((reg4019 ?
                          ((^reg3973) ?
                              forvar4034[(3'h6):(3'h5)] : (reg3995 ?
                                  (8'ha1) : reg3978)) : (reg3952 >> $unsigned(forvar3959))) >= ($signed(reg3999) ?
                          $unsigned($signed(forvar4035)) : $signed($signed(reg4039))));
                      reg4041 <= ($unsigned($signed(forvar3967)) - ((8'hb5) ?
                          (-$signed(reg3961)) : $unsigned((reg3947 ?
                              (8'h9d) : wire3943))));
                      reg4042 <= reg3947;
                    end
                  if ((^~$unsigned((reg3948 && forvar3945[(3'h7):(3'h5)]))))
                    begin
                      reg4043 <= $unsigned((forvar3949 ?
                          {$signed(reg4016)} : $signed(reg4046)));
                    end
                  else
                    begin
                      reg4043 <= ($unsigned($unsigned(reg3987[(4'ha):(2'h3)])) == reg3955);
                    end
                  if ($unsigned(((~(forvar4003 > reg4046)) ?
                      reg4019 : {(reg4006 ? forvar3983 : reg3966)})))
                    begin
                      reg4044 <= ((8'h9e) ?
                          reg4022 : $unsigned((reg3998[(4'h9):(3'h4)] ?
                              {forvar4038} : (!reg3953))));
                      reg4045 <= $unsigned((reg4019 || $unsigned($signed(reg3955))));
                    end
                  else
                    begin
                      reg4044 <= $signed(reg4028[(4'h8):(1'h0)]);
                      reg4045 <= (-(~|reg3997[(1'h1):(1'h0)]));
                    end
                  if ({reg3995[(2'h2):(2'h2)]})
                    begin
                      reg4046 <= $unsigned(((~&$unsigned((8'ha4))) ?
                          $signed($signed((8'hb7))) : (reg4032[(3'h4):(2'h3)] ?
                              reg4040 : $signed(reg4034))));
                      reg4047 <= {reg4041[(4'hc):(2'h2)]};
                      reg4048 <= (reg3979[(2'h3):(1'h0)] ?
                          $unsigned($signed({(8'hba)})) : (((reg4018 >= wire3943) | $unsigned(reg4037)) ?
                              (reg4041 ?
                                  $unsigned(forvar4013) : (reg4016 ?
                                      reg4032 : reg4042)) : $signed($signed((8'hba)))));
                      reg4049 <= (&($signed($signed((8'h9d))) ?
                          ((8'hb3) ?
                              reg4011[(2'h2):(2'h2)] : (|(8'hb8))) : (((8'hb5) ~^ forvar3952) || {forvar3972})));
                    end
                  else
                    begin
                      reg4046 <= forvar4013;
                    end
                end
              for (forvar4050 = (1'h0); (forvar4050 < (1'h0)); forvar4050 = (forvar4050 + (1'h1)))
                begin
                  for (forvar4051 = (1'h0); (forvar4051 < (2'h3)); forvar4051 = (forvar4051 + (1'h1)))
                    begin
                      reg4052 <= ((^(+$unsigned(reg3945))) ?
                          $unsigned((reg4042 ^ (8'hb4))) : $unsigned((+(reg4001 << reg3989))));
                      reg4053 <= (!(^reg4014));
                      reg4054 <= {reg4006[(1'h1):(1'h0)]};
                      reg4055 <= {$signed({wire3937[(1'h1):(1'h1)]})};
                    end
                  if ((reg3970[(4'h8):(3'h5)] ?
                      (8'h9c) : $signed((((8'hba) ? reg4041 : reg3952) ?
                          (8'h9d) : {(8'had)}))))
                    begin
                      reg4056 <= (!((~&{forvar3948}) ?
                          (|(8'hb2)) : (reg3953[(1'h1):(1'h1)] ?
                              $signed(wire3941) : wire3943[(3'h4):(3'h4)])));
                      reg4057 <= ($signed($signed((reg4049 > reg4012))) * $unsigned((8'h9f)));
                    end
                  else
                    begin
                      reg4056 <= (reg4019[(2'h3):(2'h3)] ?
                          reg4022[(3'h7):(1'h1)] : ($unsigned((~^(8'hac))) ?
                              (-$signed((8'ha9))) : $signed((!reg3945))));
                    end
                  if ((((~^$unsigned(reg4026)) >>> reg4014) ?
                      $signed($unsigned((8'ha2))) : $unsigned($signed((8'hb3)))))
                    begin
                      reg4058 <= $unsigned($signed($signed(reg4047)));
                      reg4059 <= reg4034;
                    end
                  else
                    begin
                      reg4058 <= (-$unsigned((reg4026 >> forvar3962)));
                      reg4059 <= (((reg4045[(3'h4):(2'h3)] ?
                          (reg4058 <= reg4018) : $unsigned(reg4024)) || (reg3948[(5'h10):(1'h0)] < reg3957[(1'h0):(1'h0)])) || (((reg4049 ?
                              forvar3954 : (8'hb7)) ?
                          $unsigned((8'haa)) : forvar3950) <= (|$signed(forvar3945))));
                      reg4060 <= forvar3968[(4'h8):(1'h1)];
                      reg4061 <= ((~(|reg3995)) != (~|((!(8'hb4)) ?
                          {forvar3959} : (reg3946 || reg4037))));
                    end
                  if ({reg3956[(1'h1):(1'h1)]})
                    begin
                      reg4062 <= reg4009;
                      reg4063 <= $unsigned(($signed(reg3971) ?
                          ($signed(forvar4031) ?
                              $signed(reg3960) : ((8'ha3) > reg4061)) : ({reg3978} > (reg3951 >= reg4043))));
                      reg4064 <= forvar4020;
                      reg4065 <= ((^~reg4030[(1'h1):(1'h1)]) ?
                          $signed($unsigned((|reg3987))) : reg3975);
                    end
                  else
                    begin
                      reg4062 <= ({$signed(reg4054)} != (^~wire3940));
                      reg4063 <= (~$unsigned((^(reg3992 ?
                          forvar3985 : reg4026))));
                      reg4064 <= $signed($unsigned(((forvar3983 ?
                              reg4025 : reg3991) ?
                          $unsigned(reg3973) : reg4065)));
                    end
                end
              if ($unsigned($unsigned($signed((|reg4053)))))
                begin
                  reg4066 <= {(^~{reg3965[(3'h6):(1'h0)]})};
                  if ($signed(reg4037[(4'hb):(1'h1)]))
                    begin
                      reg4067 <= $signed((wire3940[(1'h0):(1'h0)] ?
                          forvar4044[(4'hf):(1'h0)] : (((8'haf) << reg4009) << ((8'hb2) ?
                              reg4037 : reg3953))));
                      reg4068 <= (((reg3974[(2'h3):(1'h0)] ?
                              $unsigned(reg4044) : reg3946[(2'h3):(1'h1)]) & reg4040[(4'h8):(2'h3)]) ?
                          (8'ha7) : (-(reg4009 != forvar3985)));
                      reg4069 <= ($signed(reg4018[(4'h8):(2'h2)]) <<< $unsigned({(reg3999 ?
                              wire3937 : forvar4033)}));
                    end
                  else
                    begin
                      reg4067 <= $signed((($unsigned(reg4028) > (+reg3974)) ?
                          forvar4035 : $unsigned($signed(reg4031))));
                      reg4068 <= (reg4022[(3'h5):(1'h0)] - ({reg3968} ?
                          $signed((forvar3962 ?
                              forvar3962 : forvar3993)) : reg4055[(2'h2):(1'h1)]));
                      reg4069 <= ({$unsigned((-wire3938))} | (((reg3969 >>> forvar4020) ?
                          $unsigned(reg4046) : {(8'ha9)}) >>> reg3988));
                      reg4070 <= $unsigned($signed((&reg3950[(2'h3):(1'h0)])));
                    end
                end
              else
                begin
                  if (($signed((8'hac)) - reg4036[(1'h0):(1'h0)]))
                    begin
                      reg4066 <= reg4053;
                      reg4067 <= reg4061;
                    end
                  else
                    begin
                      reg4066 <= $unsigned(reg3976);
                    end
                  reg4068 <= ({reg4025[(3'h6):(2'h2)]} < (~|forvar4013));
                  reg4069 <= ((~(~|reg3990)) ?
                      $unsigned(((-(8'hb9)) != $signed(reg3952))) : $unsigned((-$unsigned(reg3988))));
                  if ($unsigned((reg3948 ?
                      reg4016[(3'h6):(2'h2)] : (^$unsigned(wire3940)))))
                    begin
                      reg4070 <= ({reg4025[(4'hf):(3'h4)]} >= (-{wire3942[(1'h1):(1'h1)]}));
                    end
                  else
                    begin
                      reg4070 <= $signed(reg4030[(1'h0):(1'h0)]);
                    end
                end
            end
          if ($unsigned($unsigned((+forvar4015))))
            begin
              reg4071 <= $signed((((~|(8'hb9)) & (^reg4008)) ?
                  reg4066 : ({reg4035} ?
                      $signed(reg3951) : ((8'hb8) || reg3998))));
              for (forvar4072 = (1'h0); (forvar4072 < (1'h0)); forvar4072 = (forvar4072 + (1'h1)))
                begin
                  if ($unsigned($unsigned((forvar3959[(2'h2):(1'h1)] * (reg3951 ?
                      reg4049 : forvar3983)))))
                    begin
                      reg4073 <= $signed(((8'hb8) ?
                          $signed(reg4063[(4'h8):(2'h2)]) : (~$signed(reg4053))));
                    end
                  else
                    begin
                      reg4073 <= $signed({forvar4028[(2'h2):(1'h0)]});
                      reg4074 <= forvar4051[(2'h2):(1'h0)];
                      reg4075 <= ($signed(((!reg3955) ?
                          forvar3975 : reg3995[(1'h1):(1'h1)])) == {({reg3948} - $signed(reg4029))});
                    end
                  for (forvar4076 = (1'h0); (forvar4076 < (2'h3)); forvar4076 = (forvar4076 + (1'h1)))
                    begin
                      reg4077 <= forvar3972;
                      reg4078 <= $signed(reg4039);
                    end
                  if ((~$signed(($unsigned(reg4018) ?
                      $signed(reg3949) : reg3945[(3'h7):(3'h5)]))))
                    begin
                      reg4079 <= reg3975[(4'hb):(3'h7)];
                      reg4080 <= $unsigned($signed((~|(&forvar3959))));
                    end
                  else
                    begin
                      reg4079 <= ((forvar3968[(4'h9):(4'h8)] ?
                              $signed(forvar3985[(4'h8):(3'h5)]) : $signed(reg3945[(4'h9):(2'h3)])) ?
                          (~^(^{reg4054})) : (^~(-$unsigned(reg3987))));
                      reg4080 <= {((~|$signed(forvar4044)) ?
                              ((reg3974 * reg4008) ?
                                  {forvar3952} : reg4048) : ($signed(reg4026) ~^ reg3958[(3'h5):(2'h3)]))};
                      reg4081 <= (((8'ha0) ?
                              ($unsigned(reg3961) ?
                                  {reg3984} : {reg3950}) : ((-reg4053) ?
                                  forvar3949[(4'ha):(2'h3)] : $signed(forvar3981))) ?
                          forvar3952 : ($signed({forvar4028}) ?
                              {(reg4058 ?
                                      reg3975 : reg4080)} : (^~$unsigned(forvar4038))));
                    end
                end
            end
          else
            begin
              for (forvar4071 = (1'h0); (forvar4071 < (1'h1)); forvar4071 = (forvar4071 + (1'h1)))
                begin
                  for (forvar4072 = (1'h0); (forvar4072 < (1'h0)); forvar4072 = (forvar4072 + (1'h1)))
                    begin
                      reg4073 <= (|$signed($unsigned((|reg4015))));
                      reg4074 <= $signed({(|(forvar4038 ? (8'hb5) : reg4041))});
                      reg4075 <= (|$unsigned($unsigned($signed(reg3980))));
                      reg4076 <= (reg3987[(1'h1):(1'h0)] ?
                          $unsigned(($signed(reg4022) ~^ forvar4033[(4'hf):(4'hd)])) : (+($signed((8'ha9)) > $unsigned(reg4060))));
                    end
                  reg4077 <= {reg4016[(3'h7):(1'h1)]};
                end
              for (forvar4078 = (1'h0); (forvar4078 < (1'h0)); forvar4078 = (forvar4078 + (1'h1)))
                begin
                  if (((^((reg4055 - forvar3968) ?
                          reg4064[(3'h7):(1'h0)] : reg3969[(2'h2):(1'h0)])) ?
                      reg4035 : (!(((8'h9d) ? reg3978 : forvar4034) ?
                          forvar4003[(4'h8):(2'h3)] : (reg3976 ?
                              reg3953 : forvar4013)))))
                    begin
                      reg4079 <= reg3995[(2'h2):(1'h0)];
                      reg4080 <= reg3958[(4'h8):(3'h6)];
                      reg4081 <= (&(wire3942[(3'h4):(1'h1)] != {(forvar3952 ^~ reg4078)}));
                    end
                  else
                    begin
                      reg4079 <= (|$signed(reg4058[(4'h9):(4'h9)]));
                      reg4080 <= (|((reg4024[(3'h5):(1'h0)] > reg3991) & (reg4035[(3'h6):(2'h3)] ?
                          forvar3952[(3'h4):(1'h1)] : $unsigned((8'haf)))));
                      reg4081 <= reg4058[(3'h4):(2'h2)];
                      reg4082 <= ({$unsigned($unsigned(reg4018))} ?
                          wire3943[(3'h5):(2'h2)] : $unsigned(reg3984));
                    end
                  if (($signed(($unsigned(reg4029) && $unsigned(reg4001))) > $unsigned(reg4041[(2'h2):(1'h0)])))
                    begin
                      reg4083 <= ($signed(reg3996) ~^ $signed(reg3992));
                      reg4084 <= (($signed((!forvar4017)) >> reg4010) << (!$unsigned((forvar4044 - (8'ha3)))));
                      reg4085 <= (reg4056[(1'h0):(1'h0)] ?
                          forvar4031 : (($unsigned(reg4016) ?
                              forvar3967 : $unsigned(reg4041)) >> (+reg3946[(3'h4):(1'h0)])));
                    end
                  else
                    begin
                      reg4083 <= reg3973;
                      reg4084 <= forvar4023;
                      reg4085 <= ({reg4014[(4'hc):(1'h1)]} <<< reg3956);
                    end
                  if ({$signed(forvar4071[(3'h6):(3'h6)])})
                    begin
                      reg4086 <= $signed(reg4042);
                      reg4087 <= ($signed((reg4007[(4'h9):(2'h2)] ^~ reg4011)) ^~ (((|forvar3993) <= {reg4067}) < $unsigned($signed((8'haa)))));
                    end
                  else
                    begin
                      reg4086 <= reg4046;
                      reg4087 <= reg3968[(1'h0):(1'h0)];
                      reg4088 <= $signed(forvar4023[(4'hd):(1'h1)]);
                    end
                  if (($signed((~^(+reg4004))) ?
                      $unsigned(($unsigned(forvar4034) ?
                          reg3991 : (reg4036 ?
                              reg3992 : reg3956))) : ((~^reg3999) ?
                          $unsigned(((8'ha2) ^~ reg4000)) : (reg4064[(2'h2):(1'h1)] ?
                              (forvar4031 ?
                                  reg3957 : reg4021) : reg4061[(1'h1):(1'h1)]))))
                    begin
                      reg4089 <= reg3976;
                      reg4090 <= ((~|$unsigned(reg4084)) ?
                          ((reg3978[(3'h7):(3'h7)] >= $unsigned((8'ha6))) >> ((forvar3967 ?
                              forvar4015 : reg4033) + $unsigned(reg3976))) : ($signed(wire3940[(1'h0):(1'h0)]) ~^ wire3944));
                    end
                  else
                    begin
                      reg4089 <= $unsigned(reg4001);
                    end
                end
              if ($signed({reg4032}))
                begin
                  for (forvar4091 = (1'h0); (forvar4091 < (2'h2)); forvar4091 = (forvar4091 + (1'h1)))
                    begin
                      reg4092 <= ($signed({reg4049[(3'h4):(1'h0)]}) > $signed($unsigned((forvar3967 ?
                          forvar4038 : reg4083))));
                      reg4093 <= {reg3966[(1'h0):(1'h0)]};
                      reg4094 <= {(forvar3949[(3'h6):(3'h5)] ?
                              reg4033 : ((!reg4043) && {reg3973}))};
                      reg4095 <= ({$unsigned($unsigned(reg4054))} > $signed((8'ha0)));
                    end
                end
              else
                begin
                  if (((~|reg4078[(2'h3):(2'h2)]) ?
                      ((forvar4033[(3'h4):(3'h4)] ^ (forvar3967 >= forvar3972)) * forvar3952[(4'h9):(1'h0)]) : {reg4082}))
                    begin
                      reg4091 <= (^(|($unsigned(reg4062) ?
                          reg3995[(2'h2):(1'h0)] : reg4032[(3'h5):(3'h5)])));
                    end
                  else
                    begin
                      reg4091 <= (&reg4040);
                      reg4092 <= reg3958[(2'h2):(2'h2)];
                    end
                  if ((~$signed((~^(~|(8'hb7))))))
                    begin
                      reg4093 <= reg4016[(1'h0):(1'h0)];
                      reg4094 <= $unsigned($signed($signed({(8'ha0)})));
                    end
                  else
                    begin
                      reg4093 <= $unsigned((8'h9c));
                      reg4094 <= (reg4080[(3'h4):(2'h3)] ?
                          (~&$signed(forvar3952)) : $signed(reg3948));
                      reg4095 <= (+($unsigned(forvar4044) ?
                          {reg3964} : ({reg4019} ?
                              (reg4045 ? wire3939 : reg4046) : (8'hba))));
                      reg4096 <= reg3970;
                    end
                end
            end
        end
      else
        begin
          if (reg3992)
            begin
              reg3981 <= ($unsigned((8'hb6)) ?
                  (((8'hb9) ?
                      $signed(forvar3975) : (reg4016 >> forvar4033)) >> ((forvar4031 ?
                      reg3991 : reg4033) != reg4039)) : ({reg3949} ^~ forvar4034));
            end
          else
            begin
              if ($unsigned((8'hb1)))
                begin
                  for (forvar3981 = (1'h0); (forvar3981 < (1'h0)); forvar3981 = (forvar3981 + (1'h1)))
                    begin
                      reg3982 <= ((8'h9d) ?
                          reg3971[(4'h9):(4'h8)] : forvar4035[(3'h6):(2'h2)]);
                      reg3983 <= $unsigned(reg4073[(3'h5):(1'h1)]);
                      reg3984 <= {(+reg4049[(3'h5):(1'h1)])};
                    end
                  for (forvar3985 = (1'h0); (forvar3985 < (1'h1)); forvar3985 = (forvar3985 + (1'h1)))
                    begin
                      reg3986 <= ($signed(({reg4012} >= (&reg4095))) ?
                          (!forvar3968) : ($signed((reg4065 <= forvar3962)) ?
                              $unsigned($unsigned((8'hb6))) : $unsigned($unsigned(forvar4076))));
                      reg3987 <= forvar3945[(1'h1):(1'h0)];
                      reg3988 <= reg4046[(2'h3):(2'h2)];
                    end
                end
              else
                begin
                  reg3981 <= (+reg4064[(3'h5):(2'h2)]);
                  if (reg4054[(1'h1):(1'h1)])
                    begin
                      reg3982 <= ((~^$unsigned((reg4059 <<< reg4039))) ?
                          reg4059[(1'h1):(1'h1)] : $signed(((&reg3994) ^ (reg3956 ?
                              reg3977 : forvar4071))));
                      reg3983 <= reg4030;
                    end
                  else
                    begin
                      reg3982 <= wire3937[(1'h1):(1'h1)];
                      reg3983 <= (~&(~|reg4075[(3'h7):(1'h0)]));
                      reg3984 <= reg3998;
                      reg3985 <= $unsigned((reg4064[(2'h3):(2'h3)] ?
                          forvar3975 : $unsigned((reg4069 || reg3999))));
                    end
                  if (reg4095[(3'h6):(3'h4)])
                    begin
                      reg3986 <= (|reg4063[(4'hc):(2'h3)]);
                      reg3987 <= ($unsigned(($unsigned(forvar4020) ?
                              $signed(reg4086) : (reg4008 <= reg3948))) ?
                          wire3943 : ((reg4006[(1'h0):(1'h0)] >> $unsigned(reg4096)) || reg3961[(4'h8):(2'h2)]));
                      reg3988 <= reg4091[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg3986 <= $unsigned(forvar3962);
                      reg3987 <= (&(+($unsigned(reg4009) * (reg4019 + reg4059))));
                      reg3988 <= (!reg4016);
                      reg3989 <= $unsigned($signed((~&(^reg3984))));
                    end
                  if (reg4070)
                    begin
                      reg3990 <= $signed((reg4004[(1'h1):(1'h0)] ?
                          reg4065[(3'h7):(3'h6)] : (8'ha2)));
                      reg3991 <= (8'hb0);
                      reg3992 <= (!reg3974[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg3990 <= forvar4035[(4'ha):(4'h8)];
                      reg3991 <= (-{({forvar4035} ?
                              {reg3982} : forvar4028[(1'h0):(1'h0)])});
                    end
                end
              if (($unsigned($signed((reg4080 ^ reg4046))) ?
                  {(8'ha0)} : $unsigned((+(|reg4073)))))
                begin
                  for (forvar3993 = (1'h0); (forvar3993 < (1'h0)); forvar3993 = (forvar3993 + (1'h1)))
                    begin
                      reg3994 <= $signed(((|$signed(reg3983)) ^~ ((forvar3982 ?
                          (8'ha2) : forvar4038) >= $unsigned(wire3942))));
                      reg3995 <= ($signed((^~(~reg4032))) && ({$signed(forvar4038)} ?
                          reg4078[(1'h1):(1'h1)] : (~&$unsigned(reg3987))));
                      reg3996 <= $signed(reg4054);
                    end
                  if ($unsigned($signed((+$signed((8'hb3))))))
                    begin
                      reg3997 <= $unsigned({reg3950});
                      reg3998 <= $signed({{$signed((8'h9d))}});
                      reg3999 <= $unsigned(wire3942[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg3997 <= $signed($signed(forvar3952));
                      reg3998 <= reg3982;
                    end
                  if (reg4049)
                    begin
                      reg4000 <= (8'hb1);
                      reg4001 <= $signed($unsigned($unsigned($signed(reg4069))));
                    end
                  else
                    begin
                      reg4000 <= reg4076[(4'h8):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar3993 = (1'h0); (forvar3993 < (1'h1)); forvar3993 = (forvar3993 + (1'h1)))
                    begin
                      reg3994 <= forvar3985[(3'h4):(1'h1)];
                      reg3995 <= ($signed(reg4064) ?
                          $unsigned((reg4066 ~^ forvar3982)) : $unsigned(reg4043[(4'ha):(3'h6)]));
                    end
                  if ((reg4095[(3'h4):(3'h4)] && reg4059))
                    begin
                      reg3996 <= ((8'h9d) ?
                          $signed(((^reg4039) ?
                              (-wire3944) : ((8'ha4) ^~ reg3966))) : (reg4049[(3'h5):(3'h5)] | forvar4038));
                      reg3997 <= reg3983[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg3996 <= (((8'ha0) ^~ ($signed(reg4064) ?
                              {reg4036} : $unsigned(reg4022))) ?
                          ((!(&(8'hab))) ?
                              ((reg4015 ? (8'haf) : reg3971) ?
                                  $unsigned(reg4075) : reg4063[(4'ha):(3'h5)]) : ((forvar3968 ~^ reg3965) ?
                                  (8'hb0) : (reg4071 ?
                                      forvar4035 : (8'hb0)))) : forvar4071[(3'h7):(3'h6)]);
                      reg3997 <= $unsigned(($signed((reg4092 ^ (8'had))) >> $signed(reg4070)));
                      reg3998 <= {reg4006[(2'h2):(1'h1)]};
                      reg3999 <= $signed(({(reg4084 ?
                              reg4045 : reg4044)} >= $unsigned({reg4033})));
                    end
                  reg4000 <= (!((forvar3950 ?
                          (|forvar3981) : $signed(reg4046)) ?
                      (reg4087 ?
                          {reg4085} : reg4057[(3'h6):(1'h1)]) : $unsigned(reg4086[(4'ha):(4'h9)])));
                  if (reg3999[(4'hc):(3'h5)])
                    begin
                      reg4001 <= reg3978[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg4001 <= $unsigned(reg3960);
                      reg4002 <= ((&($unsigned(reg3980) + (reg4042 ?
                              forvar4005 : (8'hb3)))) ?
                          $unsigned($signed((reg4039 << forvar4033))) : (^((reg4041 ?
                              reg3999 : reg4079) & (reg4012 + reg4081))));
                      reg4003 <= $signed((8'hb9));
                    end
                end
              for (forvar4004 = (1'h0); (forvar4004 < (1'h0)); forvar4004 = (forvar4004 + (1'h1)))
                begin
                  for (forvar4005 = (1'h0); (forvar4005 < (2'h3)); forvar4005 = (forvar4005 + (1'h1)))
                    begin
                      reg4006 <= $signed({(8'had)});
                      reg4007 <= ((($signed(reg4092) ?
                              reg4007[(2'h3):(2'h3)] : (reg3976 && reg3980)) ?
                          reg4025 : (8'ha0)) ^~ $signed($unsigned(reg3955)));
                      reg4008 <= (^~(~&({(8'ha0)} - reg4014[(4'hb):(4'ha)])));
                      reg4009 <= (forvar3945 ?
                          $signed($signed($signed(reg4026))) : {($signed((8'ha4)) ?
                                  $unsigned(reg4049) : $signed(reg4044))});
                    end
                  if ((~^forvar3975[(1'h0):(1'h0)]))
                    begin
                      reg4010 <= $unsigned((8'had));
                      reg4011 <= wire3940;
                      reg4012 <= ((^$signed({(8'h9d)})) ?
                          {(-(reg3999 >> reg4033))} : {(reg3975[(4'h8):(1'h1)] ?
                                  $signed(reg3975) : $signed(reg3987))});
                    end
                  else
                    begin
                      reg4010 <= reg4008[(1'h0):(1'h0)];
                      reg4011 <= ((($signed(reg4073) >>> reg3989[(4'hb):(1'h1)]) ?
                          $unsigned($unsigned(forvar4013)) : $unsigned(forvar4051[(2'h3):(2'h3)])) <<< (reg3999 < $signed($unsigned(reg3976))));
                      reg4012 <= (|forvar4017[(1'h1):(1'h1)]);
                    end
                end
              for (forvar4013 = (1'h0); (forvar4013 < (2'h3)); forvar4013 = (forvar4013 + (1'h1)))
                begin
                  if ($signed((+(&{reg3984}))))
                    begin
                      reg4014 <= (wire3939[(1'h0):(1'h0)] ?
                          ((~$unsigned(reg3948)) ~^ ($signed(wire3939) & forvar4013[(4'ha):(3'h5)])) : ($unsigned(reg4033[(1'h1):(1'h1)]) ?
                              $unsigned({reg3958}) : $unsigned(forvar3948)));
                    end
                  else
                    begin
                      reg4014 <= {forvar4035[(4'hd):(4'hc)]};
                    end
                end
            end
          for (forvar4015 = (1'h0); (forvar4015 < (2'h2)); forvar4015 = (forvar4015 + (1'h1)))
            begin
              if ($signed(($unsigned((reg3955 <= reg3945)) >>> (wire3944 ?
                  $unsigned((8'ha1)) : (|(8'ha4))))))
                begin
                  reg4016 <= ($signed($unsigned($unsigned(reg4052))) & (~reg3996[(1'h1):(1'h1)]));
                  for (forvar4017 = (1'h0); (forvar4017 < (1'h0)); forvar4017 = (forvar4017 + (1'h1)))
                    begin
                      reg4018 <= (^{$unsigned($signed((8'h9e)))});
                    end
                  reg4019 <= ($signed(reg4076) ?
                      ((((8'ha9) ? forvar4003 : forvar4078) ?
                              $unsigned(reg4024) : $signed(forvar3959)) ?
                          (reg3999[(4'hc):(4'ha)] ?
                              (reg3958 | forvar3981) : $signed(reg3965)) : reg3998) : $signed($unsigned($unsigned((8'hb0)))));
                  for (forvar4020 = (1'h0); (forvar4020 < (1'h0)); forvar4020 = (forvar4020 + (1'h1)))
                    begin
                      reg4021 <= $unsigned((forvar3986[(1'h0):(1'h0)] < (~|(^reg4036))));
                      reg4022 <= $signed($signed($signed($signed(reg4029))));
                      reg4023 <= ((((-reg3989) != forvar3967[(1'h1):(1'h1)]) ^ reg4014) ?
                          $unsigned(reg3969[(1'h0):(1'h0)]) : forvar4017[(2'h2):(1'h0)]);
                    end
                end
              else
                begin
                  reg4016 <= {$signed(forvar4044[(2'h3):(1'h1)])};
                  for (forvar4017 = (1'h0); (forvar4017 < (1'h0)); forvar4017 = (forvar4017 + (1'h1)))
                    begin
                      reg4018 <= $signed({$unsigned({reg4068})});
                    end
                  reg4019 <= $signed(({forvar3985[(3'h7):(2'h2)]} ~^ (^~$signed((8'ha4)))));
                end
              if (($signed(({reg4079} >>> (reg3955 & reg3971))) ?
                  $unsigned($unsigned({reg3947})) : reg4032[(3'h7):(3'h4)]))
                begin
                  for (forvar4024 = (1'h0); (forvar4024 < (1'h1)); forvar4024 = (forvar4024 + (1'h1)))
                    begin
                      reg4025 <= $unsigned(reg4063);
                      reg4026 <= reg4042;
                      reg4027 <= reg4035;
                      reg4028 <= (^reg3973[(4'h9):(3'h4)]);
                    end
                  for (forvar4029 = (1'h0); (forvar4029 < (2'h3)); forvar4029 = (forvar4029 + (1'h1)))
                    begin
                      reg4030 <= forvar3985[(1'h0):(1'h0)];
                      reg4031 <= $unsigned({{reg3996[(3'h4):(2'h3)]}});
                      reg4032 <= (^($unsigned(reg3950[(1'h1):(1'h1)]) ?
                          ($signed((8'h9e)) ?
                              $unsigned(reg3986) : (reg4094 ~^ (8'hb6))) : reg4078));
                    end
                end
              else
                begin
                  if ((-$signed($signed((&(8'hb4))))))
                    begin
                      reg4024 <= (($unsigned((^~reg4014)) + forvar3967[(3'h4):(2'h2)]) > (^~{wire3939}));
                      reg4025 <= (8'hb6);
                      reg4026 <= ((~^(~&reg4064)) ?
                          ({reg4084} ?
                              ((reg3980 ?
                                  reg3989 : reg4032) ^~ reg3991) : $signed((forvar3993 + reg4056))) : forvar4034);
                      reg4027 <= (({{(8'hb1)}} ?
                          (|(reg4067 >>> (8'haf))) : (-forvar3993[(1'h0):(1'h0)])) >= (reg3974[(2'h3):(1'h0)] <<< (+(reg4052 ?
                          reg3950 : reg4033))));
                    end
                  else
                    begin
                      reg4024 <= ($unsigned((8'hb2)) << (-$unsigned(((8'h9e) ?
                          reg4054 : reg4086))));
                      reg4025 <= (forvar4005 ?
                          $signed($signed((forvar4044 ?
                              forvar3982 : forvar4050))) : reg3950[(2'h3):(1'h0)]);
                      reg4026 <= reg3981[(1'h0):(1'h0)];
                    end
                  if (({(+$signed(reg3975))} != reg3996[(3'h4):(2'h2)]))
                    begin
                      reg4028 <= (&(((reg3991 ? reg3994 : (8'hb4)) ?
                          (reg4012 ?
                              forvar4034 : forvar4017) : {forvar3972}) > ($unsigned(reg4063) <<< reg4074[(4'hc):(2'h2)])));
                      reg4029 <= reg4012[(2'h2):(1'h0)];
                      reg4030 <= $unsigned(forvar3959[(3'h5):(3'h4)]);
                      reg4031 <= $unsigned(((-(reg3946 | reg3960)) ~^ ((forvar4076 + forvar3983) * $signed(reg4019))));
                    end
                  else
                    begin
                      reg4028 <= reg4015;
                    end
                  if ($signed(reg4034))
                    begin
                      reg4032 <= (8'ha5);
                    end
                  else
                    begin
                      reg4032 <= (^~(reg4047[(3'h4):(1'h0)] - $unsigned(reg4073)));
                      reg4033 <= (reg4024[(3'h5):(1'h1)] ?
                          reg4071[(2'h2):(1'h1)] : (reg3950 ?
                              (reg4026[(1'h1):(1'h1)] ?
                                  (reg3965 ?
                                      reg4062 : reg4047) : $unsigned(forvar3945)) : (^((8'hb7) - forvar4020))));
                      reg4034 <= $unsigned(($signed($signed(reg3980)) == reg3983));
                      reg4035 <= {$unsigned($signed($signed(reg4058)))};
                    end
                end
              for (forvar4036 = (1'h0); (forvar4036 < (1'h1)); forvar4036 = (forvar4036 + (1'h1)))
                begin
                  for (forvar4037 = (1'h0); (forvar4037 < (1'h0)); forvar4037 = (forvar4037 + (1'h1)))
                    begin
                      reg4038 <= reg4026[(4'h8):(2'h3)];
                    end
                  if ((-({(reg4088 ?
                          reg4041 : reg4054)} != {(forvar4071 ^ reg3996)})))
                    begin
                      reg4039 <= $unsigned($unsigned(forvar4037));
                    end
                  else
                    begin
                      reg4039 <= (~^$signed($signed(reg4011[(2'h3):(2'h2)])));
                      reg4040 <= reg3970;
                    end
                  if (({((-reg4076) ?
                          reg3958[(4'h8):(3'h4)] : (reg4031 ?
                              (8'hb0) : forvar3959))} >= (($signed(reg4074) ?
                      reg3985[(4'ha):(3'h5)] : (reg4079 ?
                          reg4029 : reg4010)) && (~(8'hb2)))))
                    begin
                      reg4041 <= (!$signed($unsigned({(8'ha8)})));
                      reg4042 <= reg4030;
                      reg4043 <= $signed((8'h9e));
                      reg4044 <= (+(((^reg4065) ?
                          reg4067[(3'h7):(2'h3)] : forvar4044[(1'h0):(1'h0)]) >>> ({reg3971} || $signed(reg4080))));
                    end
                  else
                    begin
                      reg4041 <= $signed((|$signed(reg3965[(2'h2):(1'h0)])));
                      reg4042 <= (~&(reg3988[(3'h7):(3'h6)] ^~ ((forvar4078 ?
                          wire3944 : (8'haf)) & $signed(forvar4013))));
                    end
                  reg4045 <= reg4011;
                end
              for (forvar4046 = (1'h0); (forvar4046 < (1'h1)); forvar4046 = (forvar4046 + (1'h1)))
                begin
                  for (forvar4047 = (1'h0); (forvar4047 < (2'h2)); forvar4047 = (forvar4047 + (1'h1)))
                    begin
                      reg4048 <= {$unsigned(reg4094[(1'h1):(1'h0)])};
                      reg4049 <= reg4012[(2'h3):(1'h0)];
                      reg4050 <= $signed($unsigned(reg3965));
                    end
                  if ($unsigned((reg4079[(1'h1):(1'h0)] + {(+reg4048)})))
                    begin
                      reg4051 <= $unsigned(($unsigned($unsigned((8'ha9))) ?
                          $signed($unsigned(reg4050)) : (((8'hb7) ?
                                  reg3978 : reg4067) ?
                              {(8'ha7)} : (+(8'h9f)))));
                      reg4052 <= $unsigned((!((-reg3984) ?
                          forvar3968[(1'h1):(1'h1)] : $signed((8'ha6)))));
                      reg4053 <= reg4076;
                    end
                  else
                    begin
                      reg4051 <= (~&reg3958);
                    end
                  for (forvar4054 = (1'h0); (forvar4054 < (2'h2)); forvar4054 = (forvar4054 + (1'h1)))
                    begin
                      reg4055 <= ({$signed(((8'haa) ^ wire3939))} ?
                          reg4039[(3'h6):(3'h4)] : {forvar4046});
                      reg4056 <= (wire3939[(3'h6):(2'h3)] >>> (reg4004[(1'h0):(1'h0)] >= ((reg4018 << forvar3950) ?
                          (reg3992 ? forvar3985 : reg3961) : forvar4047)));
                      reg4057 <= $unsigned($unsigned((^~reg4015[(3'h4):(2'h3)])));
                    end
                end
            end
          if ((reg4090[(2'h2):(1'h0)] ?
              reg4021 : ((!(~&reg4080)) && {$signed(reg3979)})))
            begin
              reg4058 <= (~|forvar4054[(3'h4):(1'h1)]);
              for (forvar4059 = (1'h0); (forvar4059 < (1'h0)); forvar4059 = (forvar4059 + (1'h1)))
                begin
                  for (forvar4060 = (1'h0); (forvar4060 < (2'h3)); forvar4060 = (forvar4060 + (1'h1)))
                    begin
                      reg4061 <= $unsigned((reg3978[(3'h7):(1'h1)] ?
                          (~^(reg4035 ~^ reg4068)) : ((forvar4051 ?
                                  forvar4034 : wire3938) ?
                              reg3965[(4'hc):(3'h5)] : $signed(reg3948))));
                      reg4062 <= wire3943[(2'h3):(2'h2)];
                      reg4063 <= {forvar3981[(1'h1):(1'h0)]};
                      reg4064 <= reg3949;
                    end
                  if ($signed((&$unsigned($signed(reg4028)))))
                    begin
                      reg4065 <= reg3946[(2'h3):(2'h2)];
                      reg4066 <= (reg4082[(4'he):(4'ha)] ?
                          forvar4054[(3'h5):(1'h1)] : (reg3983[(3'h7):(3'h6)] ?
                              forvar4059[(4'hd):(2'h2)] : $unsigned({reg3960})));
                      reg4067 <= $unsigned((reg4094 - $unsigned((+reg3952))));
                    end
                  else
                    begin
                      reg4065 <= reg3978[(2'h2):(1'h1)];
                    end
                end
              reg4068 <= $signed({(((8'ha8) ? (8'h9d) : reg4081) << reg3989)});
              for (forvar4069 = (1'h0); (forvar4069 < (1'h0)); forvar4069 = (forvar4069 + (1'h1)))
                begin
                  reg4070 <= $signed(reg4087);
                  reg4071 <= $unsigned(reg4011);
                  for (forvar4072 = (1'h0); (forvar4072 < (1'h0)); forvar4072 = (forvar4072 + (1'h1)))
                    begin
                      reg4073 <= ($signed({(reg4014 < forvar3945)}) ?
                          (-forvar4003) : wire3944);
                      reg4074 <= (8'hb0);
                    end
                  for (forvar4075 = (1'h0); (forvar4075 < (2'h3)); forvar4075 = (forvar4075 + (1'h1)))
                    begin
                      reg4076 <= reg4093[(2'h2):(1'h1)];
                      reg4077 <= ($signed({reg3976}) ?
                          ((reg4066 && (reg4009 ? reg3961 : reg3964)) ?
                              ((reg4086 ? reg4031 : forvar4078) ?
                                  {forvar3968} : $signed(reg4068)) : {(reg4048 ?
                                      forvar3968 : reg3945)}) : reg4050[(1'h0):(1'h0)]);
                      reg4078 <= reg4012[(4'h8):(3'h6)];
                    end
                end
            end
          else
            begin
              for (forvar4058 = (1'h0); (forvar4058 < (2'h3)); forvar4058 = (forvar4058 + (1'h1)))
                begin
                  for (forvar4059 = (1'h0); (forvar4059 < (1'h1)); forvar4059 = (forvar4059 + (1'h1)))
                    begin
                      reg4060 <= (8'hae);
                      reg4061 <= (((^~(~|forvar4046)) ^ forvar3950) >> (!{reg3971[(3'h7):(3'h6)]}));
                      reg4062 <= forvar4023;
                      reg4063 <= forvar4027[(4'he):(1'h1)];
                    end
                  if ($unsigned((~^(8'h9d))))
                    begin
                      reg4064 <= ((~^reg3987) == ((|(+(8'hb5))) * (reg4034 >> forvar4036[(4'ha):(3'h7)])));
                      reg4065 <= (8'h9f);
                    end
                  else
                    begin
                      reg4064 <= $signed(reg4023[(1'h0):(1'h0)]);
                      reg4065 <= {($unsigned((~reg4064)) ?
                              $signed(forvar3959) : reg3947)};
                    end
                  if (reg4037)
                    begin
                      reg4066 <= $unsigned((reg4088 ?
                          $signed((reg4012 > forvar4069)) : forvar3962[(2'h3):(2'h3)]));
                      reg4067 <= $signed($unsigned(forvar4020[(2'h3):(1'h1)]));
                      reg4068 <= reg4052[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg4066 <= reg3965[(4'hc):(4'ha)];
                      reg4067 <= ((+$unsigned((reg4043 ?
                              forvar3945 : forvar3993))) ?
                          (8'ha0) : (+forvar4037[(4'h9):(3'h4)]));
                      reg4068 <= ({(|$unsigned(reg4093))} ?
                          reg3990 : $signed(wire3939[(1'h1):(1'h1)]));
                    end
                  reg4069 <= (~&(reg4064 != {(wire3937 ?
                          forvar4005 : reg4071)}));
                end
            end
        end
      if (($unsigned($unsigned((&reg3983))) <= $signed(forvar4071[(2'h2):(2'h2)])))
        begin
          for (forvar4097 = (1'h0); (forvar4097 < (1'h0)); forvar4097 = (forvar4097 + (1'h1)))
            begin
              for (forvar4098 = (1'h0); (forvar4098 < (2'h3)); forvar4098 = (forvar4098 + (1'h1)))
                begin
                  reg4099 <= (reg3977[(1'h0):(1'h0)] ? {reg3964} : forvar3945);
                  for (forvar4100 = (1'h0); (forvar4100 < (2'h2)); forvar4100 = (forvar4100 + (1'h1)))
                    begin
                      reg4101 <= reg4068[(2'h3):(1'h0)];
                      reg4102 <= reg4060[(2'h2):(2'h2)];
                    end
                end
              for (forvar4103 = (1'h0); (forvar4103 < (2'h3)); forvar4103 = (forvar4103 + (1'h1)))
                begin
                  for (forvar4104 = (1'h0); (forvar4104 < (1'h0)); forvar4104 = (forvar4104 + (1'h1)))
                    begin
                      reg4105 <= $signed(reg4063);
                      reg4106 <= (forvar4071 ?
                          $signed($unsigned($signed(reg4042))) : (reg4080 - (forvar4040 <<< forvar3959[(1'h0):(1'h0)])));
                    end
                end
            end
          reg4107 <= reg4063;
          for (forvar4108 = (1'h0); (forvar4108 < (2'h3)); forvar4108 = (forvar4108 + (1'h1)))
            begin
              if ({$signed($unsigned(forvar4072))})
                begin
                  for (forvar4109 = (1'h0); (forvar4109 < (1'h1)); forvar4109 = (forvar4109 + (1'h1)))
                    begin
                      reg4110 <= $signed({((reg4083 ?
                              reg3946 : (8'haa)) <<< $unsigned(forvar4036))});
                      reg4111 <= forvar4046;
                    end
                  if ((~($signed((reg4088 == reg3955)) <<< (+(+reg3971)))))
                    begin
                      reg4112 <= (8'hab);
                      reg4113 <= forvar3945;
                    end
                  else
                    begin
                      reg4112 <= reg3987[(4'hc):(2'h2)];
                      reg4113 <= forvar3993;
                      reg4114 <= reg4070;
                      reg4115 <= ($signed(((forvar4071 > forvar4078) ?
                              (|(8'hb5)) : (8'hb5))) ?
                          ((reg3985 << forvar4017) ?
                              $signed(reg3958[(3'h4):(2'h3)]) : reg3950[(1'h0):(1'h0)]) : (reg4073[(2'h2):(1'h0)] < {$unsigned(reg3948)}));
                    end
                end
              else
                begin
                  if (reg3984)
                    begin
                      reg4109 <= (^$signed(((~^(8'ha0)) ?
                          reg3974 : forvar4027)));
                      reg4110 <= forvar4034[(3'h7):(3'h6)];
                      reg4111 <= forvar3986;
                      reg4112 <= {{($signed(reg4091) ?
                                  $unsigned(reg3973) : (8'hb2))}};
                    end
                  else
                    begin
                      reg4109 <= reg4091[(1'h0):(1'h0)];
                      reg4110 <= (((~|reg4058[(2'h3):(1'h1)]) ?
                              ((reg4066 ? reg4112 : reg4068) ?
                                  ((8'ha9) != (8'ha1)) : (~reg4027)) : ($signed(wire3943) & reg4030)) ?
                          reg4025 : (~&reg4067[(3'h4):(1'h1)]));
                      reg4111 <= (!(+wire3942[(1'h0):(1'h0)]));
                      reg4112 <= reg4054;
                    end
                end
              if ($unsigned(($signed(forvar3949[(3'h5):(3'h4)]) >>> (+$signed(reg3963)))))
                begin
                  reg4116 <= (!(forvar4037[(4'ha):(3'h5)] || $unsigned($unsigned(reg4030))));
                end
              else
                begin
                  reg4116 <= ($signed({$unsigned(reg3958)}) ?
                      $unsigned(reg3963[(1'h1):(1'h1)]) : forvar3985[(3'h6):(2'h2)]);
                  if ((~^{reg4069[(2'h2):(1'h0)]}))
                    begin
                      reg4117 <= $unsigned(forvar4038);
                      reg4118 <= reg4107[(1'h1):(1'h0)];
                      reg4119 <= reg4090[(1'h0):(1'h0)];
                      reg4120 <= reg3951;
                    end
                  else
                    begin
                      reg4117 <= ((8'h9e) ?
                          (8'hae) : (reg4110 ?
                              ($unsigned(reg3953) ?
                                  (~reg3998) : {reg4093}) : $unsigned((reg3976 ?
                                  reg3966 : reg4009))));
                    end
                  for (forvar4121 = (1'h0); (forvar4121 < (2'h3)); forvar4121 = (forvar4121 + (1'h1)))
                    begin
                      reg4122 <= ($unsigned(((&forvar4104) ?
                          reg3981[(1'h0):(1'h0)] : (8'ha3))) + $unsigned((~reg3953)));
                      reg4123 <= (+reg3992[(1'h0):(1'h0)]);
                    end
                  reg4124 <= (forvar4091[(3'h6):(2'h2)] < $signed($signed((^reg4074))));
                end
            end
        end
      else
        begin
          reg4097 <= reg4105[(3'h5):(2'h2)];
          for (forvar4098 = (1'h0); (forvar4098 < (2'h2)); forvar4098 = (forvar4098 + (1'h1)))
            begin
              reg4099 <= $signed($unsigned(({forvar4091} ?
                  reg4081[(1'h0):(1'h0)] : reg3979[(4'hb):(2'h3)])));
              if ($signed(({(forvar4100 ? reg3973 : forvar4029)} ?
                  (reg3955[(3'h7):(1'h0)] ?
                      $signed(reg3983) : (reg4026 - (8'ha6))) : (|reg4068[(2'h2):(1'h1)]))))
                begin
                  for (forvar4100 = (1'h0); (forvar4100 < (2'h2)); forvar4100 = (forvar4100 + (1'h1)))
                    begin
                      reg4101 <= (~$unsigned((!$signed(reg4039))));
                    end
                  for (forvar4102 = (1'h0); (forvar4102 < (1'h0)); forvar4102 = (forvar4102 + (1'h1)))
                    begin
                      reg4103 <= $signed(forvar4109);
                      reg4104 <= forvar4024;
                      reg4105 <= (~(8'ha3));
                      reg4106 <= $unsigned((($signed(forvar4103) ?
                          reg4068 : (8'hac)) << $signed($signed(reg4025))));
                    end
                  for (forvar4107 = (1'h0); (forvar4107 < (2'h3)); forvar4107 = (forvar4107 + (1'h1)))
                    begin
                      reg4108 <= (((reg3983[(4'h9):(4'h9)] ?
                          ((8'h9c) ? reg4062 : (8'ha5)) : (forvar4060 ?
                              (8'hb0) : forvar4005)) <<< (reg3945[(3'h7):(1'h0)] ?
                          $unsigned(reg4073) : (reg4026 & reg4088))) >>> reg4120[(3'h4):(3'h4)]);
                      reg4109 <= $signed((8'had));
                      reg4110 <= (~$unsigned(reg4068[(1'h1):(1'h0)]));
                      reg4111 <= reg4022;
                    end
                  if ($unsigned($unsigned(((8'hb8) > (^~reg4099)))))
                    begin
                      reg4112 <= $unsigned((((reg4031 && reg4010) ?
                          reg4046[(1'h0):(1'h0)] : reg4081) && reg3948));
                    end
                  else
                    begin
                      reg4112 <= (|((~&(|reg4021)) ^ reg4016[(2'h2):(1'h0)]));
                      reg4113 <= {$signed(wire3937)};
                    end
                end
              else
                begin
                  if (($signed({$unsigned(forvar4091)}) ?
                      (reg4093[(4'h9):(3'h6)] ?
                          ((~&reg4102) ?
                              {reg4068} : reg4015) : reg4056) : (+reg4030[(1'h0):(1'h0)])))
                    begin
                      reg4100 <= ($unsigned(reg4056[(2'h3):(2'h2)]) ?
                          reg3998[(2'h2):(1'h0)] : {(!forvar3967[(1'h1):(1'h0)])});
                    end
                  else
                    begin
                      reg4100 <= $unsigned(reg4018[(3'h7):(1'h0)]);
                      reg4101 <= $signed($signed(((reg3948 == reg4042) ?
                          (~^reg3966) : (reg3956 + reg4109))));
                    end
                end
            end
        end
      reg4125 <= forvar4100;
    end
  always
    @(posedge clk) begin
      if ((($signed(reg4105[(2'h3):(2'h2)]) ^~ ((&reg4088) ?
          reg4120[(4'ha):(4'h8)] : reg3971)) >= $signed($unsigned($unsigned((8'had))))))
        begin
          if ((8'ha1))
            begin
              for (forvar4126 = (1'h0); (forvar4126 < (2'h2)); forvar4126 = (forvar4126 + (1'h1)))
                begin
                  reg4127 <= (~$signed(reg4009));
                  for (forvar4128 = (1'h0); (forvar4128 < (1'h1)); forvar4128 = (forvar4128 + (1'h1)))
                    begin
                      reg4129 <= ($signed(((&reg4116) ?
                              $signed((8'hb1)) : (^~reg4106))) ?
                          $unsigned(reg4087) : {reg3960[(1'h1):(1'h0)]});
                      reg4130 <= $unsigned(((~^reg4064[(3'h7):(3'h5)]) ^ {(reg3957 ?
                              reg3978 : (8'hb0))}));
                      reg4131 <= ($signed((!reg4084)) ?
                          ($unsigned((reg4032 + reg3965)) ?
                              reg3999 : ($unsigned((8'hae)) != reg4057[(1'h1):(1'h1)])) : (reg4018[(3'h5):(3'h5)] ?
                              (((8'hb0) ? reg4023 : reg4019) ?
                                  (reg4059 >= reg4101) : (reg4002 + (8'hb0))) : ($signed((8'hb7)) ?
                                  (reg4025 ?
                                      reg4105 : reg4109) : reg3975[(1'h1):(1'h0)])));
                      reg4132 <= reg3977[(2'h2):(1'h1)];
                    end
                  for (forvar4133 = (1'h0); (forvar4133 < (2'h2)); forvar4133 = (forvar4133 + (1'h1)))
                    begin
                      reg4134 <= reg4090[(4'h9):(4'h8)];
                      reg4135 <= $signed(reg3991[(4'h8):(1'h0)]);
                      reg4136 <= ((reg3985 ?
                          reg4112[(4'h9):(4'h9)] : reg4062) ~^ ($unsigned(reg4019) >= ((~wire3943) ?
                          reg4063[(2'h3):(2'h2)] : (wire3939 ?
                              wire3944 : reg4119))));
                      reg4137 <= reg4090[(3'h6):(2'h3)];
                    end
                  for (forvar4138 = (1'h0); (forvar4138 < (2'h3)); forvar4138 = (forvar4138 + (1'h1)))
                    begin
                      reg4139 <= $signed((-{(|reg4027)}));
                    end
                end
            end
          else
            begin
              for (forvar4126 = (1'h0); (forvar4126 < (1'h0)); forvar4126 = (forvar4126 + (1'h1)))
                begin
                  for (forvar4127 = (1'h0); (forvar4127 < (1'h0)); forvar4127 = (forvar4127 + (1'h1)))
                    begin
                      reg4128 <= $signed($signed($signed({(8'ha6)})));
                    end
                  for (forvar4129 = (1'h0); (forvar4129 < (2'h2)); forvar4129 = (forvar4129 + (1'h1)))
                    begin
                      reg4130 <= $signed($signed((8'ha0)));
                      reg4131 <= $signed($signed((8'hab)));
                      reg4132 <= $signed({reg4083});
                      reg4133 <= ((~|reg4050[(2'h2):(2'h2)]) ?
                          reg4044 : ({$signed(reg4037)} ~^ $unsigned($signed(reg4093))));
                    end
                end
              for (forvar4134 = (1'h0); (forvar4134 < (2'h3)); forvar4134 = (forvar4134 + (1'h1)))
                begin
                  for (forvar4135 = (1'h0); (forvar4135 < (2'h2)); forvar4135 = (forvar4135 + (1'h1)))
                    begin
                      reg4136 <= {reg4090[(2'h3):(2'h3)]};
                      reg4137 <= ((+$unsigned(reg3965)) & reg4036);
                    end
                end
            end
          for (forvar4140 = (1'h0); (forvar4140 < (2'h2)); forvar4140 = (forvar4140 + (1'h1)))
            begin
              reg4141 <= (^~(~(reg4011[(3'h4):(3'h4)] ? reg4133 : (&reg3951))));
            end
          if ($unsigned(({reg3953[(1'h1):(1'h1)]} ?
              reg4012[(2'h2):(1'h1)] : (reg3952[(1'h1):(1'h0)] > (~|(8'ha4))))))
            begin
              if (reg3998)
                begin
                  for (forvar4142 = (1'h0); (forvar4142 < (1'h1)); forvar4142 = (forvar4142 + (1'h1)))
                    begin
                      reg4143 <= reg4058;
                    end
                  for (forvar4144 = (1'h0); (forvar4144 < (2'h2)); forvar4144 = (forvar4144 + (1'h1)))
                    begin
                      reg4145 <= {reg4042[(1'h0):(1'h0)]};
                      reg4146 <= reg3983[(3'h6):(3'h6)];
                    end
                end
              else
                begin
                  for (forvar4142 = (1'h0); (forvar4142 < (1'h0)); forvar4142 = (forvar4142 + (1'h1)))
                    begin
                      reg4143 <= (~|(-(~reg4123)));
                      reg4144 <= reg4117;
                      reg4145 <= $unsigned($unsigned({(^~(8'hb0))}));
                      reg4146 <= {$signed($unsigned(reg4129))};
                    end
                  reg4147 <= $signed((!(~{reg4134})));
                  for (forvar4148 = (1'h0); (forvar4148 < (1'h0)); forvar4148 = (forvar4148 + (1'h1)))
                    begin
                      reg4149 <= (^reg3961[(3'h4):(3'h4)]);
                      reg4150 <= (~^reg4132);
                      reg4151 <= ($unsigned({reg4079}) ?
                          $signed((reg3977 | (reg4033 + (8'hb3)))) : $unsigned((8'ha1)));
                      reg4152 <= ({(+{(8'h9f)})} ?
                          (!(8'h9f)) : ($signed(reg4086) == ($unsigned(reg4128) <<< ((8'hb8) >>> reg3982))));
                    end
                  for (forvar4153 = (1'h0); (forvar4153 < (2'h3)); forvar4153 = (forvar4153 + (1'h1)))
                    begin
                      reg4154 <= {reg3960};
                      reg4155 <= (reg4152 <<< $signed($unsigned((reg3964 ~^ (8'ha8)))));
                      reg4156 <= reg4044;
                    end
                end
              if (($unsigned({((8'hb4) ?
                      reg4032 : reg4011)}) | $unsigned($unsigned((reg4129 <= reg4088)))))
                begin
                  reg4157 <= {$unsigned((^(reg4035 ? (8'hb0) : reg4049)))};
                  for (forvar4158 = (1'h0); (forvar4158 < (2'h2)); forvar4158 = (forvar4158 + (1'h1)))
                    begin
                      reg4159 <= (reg4041[(2'h3):(2'h3)] ?
                          $signed((8'h9f)) : reg4095[(2'h3):(2'h2)]);
                      reg4160 <= {(reg4112[(3'h6):(3'h6)] ~^ ($signed(reg4036) ?
                              (reg4119 ? reg4044 : reg3997) : (reg4026 ?
                                  reg3980 : reg4095)))};
                      reg4161 <= ((^~(-{reg3999})) * (|(~&$signed(reg4038))));
                    end
                  reg4162 <= {(forvar4144[(4'h8):(2'h2)] > (|reg3975[(1'h0):(1'h0)]))};
                  reg4163 <= ((reg4139 ?
                          $signed((-reg4022)) : $signed((&reg3963))) ?
                      reg4038[(3'h4):(1'h1)] : (~^($signed(reg4156) ?
                          {reg4120} : {reg3966})));
                end
              else
                begin
                  for (forvar4157 = (1'h0); (forvar4157 < (2'h3)); forvar4157 = (forvar4157 + (1'h1)))
                    begin
                      reg4158 <= $signed((^reg4029[(4'h8):(2'h2)]));
                      reg4159 <= (forvar4158 ?
                          ((+$signed(reg4011)) & (reg3958 ^~ $unsigned(reg4103))) : ((|(~(8'ha3))) ?
                              forvar4128 : (reg3974 <= $unsigned(reg3979))));
                    end
                  if (($unsigned((reg4133[(3'h5):(3'h4)] * $signed((8'hae)))) <<< reg4132))
                    begin
                      reg4160 <= (wire3941[(1'h1):(1'h0)] ?
                          $signed(($unsigned(reg4113) ?
                              {reg4041} : forvar4127)) : forvar4140[(1'h1):(1'h0)]);
                      reg4161 <= reg4031[(2'h3):(1'h1)];
                      reg4162 <= $unsigned({(8'hab)});
                      reg4163 <= (reg3982 >= reg4094[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg4160 <= reg4158;
                      reg4161 <= (8'haf);
                    end
                  if (((+$signed($signed(forvar4128))) > {(reg3968[(3'h4):(3'h4)] < (^reg4007))}))
                    begin
                      reg4164 <= $unsigned((8'ha3));
                      reg4165 <= ({reg4060} > $unsigned($signed(reg3979)));
                      reg4166 <= ($unsigned({(|reg4036)}) && $signed(($signed(reg4003) ?
                          {forvar4128} : $signed(reg4038))));
                      reg4167 <= {({reg3968[(1'h0):(1'h0)]} ?
                              (8'h9c) : (8'had))};
                    end
                  else
                    begin
                      reg4164 <= $unsigned($unsigned(($unsigned(reg3958) <<< (|reg4160))));
                    end
                  for (forvar4168 = (1'h0); (forvar4168 < (2'h2)); forvar4168 = (forvar4168 + (1'h1)))
                    begin
                      reg4169 <= $signed((^~$unsigned($signed(reg4151))));
                    end
                end
              for (forvar4170 = (1'h0); (forvar4170 < (2'h2)); forvar4170 = (forvar4170 + (1'h1)))
                begin
                  for (forvar4171 = (1'h0); (forvar4171 < (1'h1)); forvar4171 = (forvar4171 + (1'h1)))
                    begin
                      reg4172 <= ((reg4135[(1'h1):(1'h1)] ?
                              ($unsigned(reg4146) <= reg4169) : reg4026[(4'hc):(1'h0)]) ?
                          {((reg4084 < (8'ha7)) ?
                                  (&forvar4158) : {reg4019})} : $signed($unsigned({reg4160})));
                    end
                  for (forvar4173 = (1'h0); (forvar4173 < (1'h1)); forvar4173 = (forvar4173 + (1'h1)))
                    begin
                      reg4174 <= reg4059[(2'h2):(1'h1)];
                      reg4175 <= (-({{reg3999}} ? reg3950 : (!reg3960)));
                      reg4176 <= reg4027[(2'h2):(1'h0)];
                    end
                  if ($unsigned(reg4090))
                    begin
                      reg4177 <= reg4156;
                      reg4178 <= $unsigned($signed((wire3937[(2'h2):(1'h1)] <<< reg4039)));
                    end
                  else
                    begin
                      reg4177 <= $unsigned(reg4089);
                      reg4178 <= $unsigned($unsigned(reg4165));
                    end
                end
              for (forvar4179 = (1'h0); (forvar4179 < (2'h2)); forvar4179 = (forvar4179 + (1'h1)))
                begin
                  if ((&(reg3992 ?
                      {$unsigned(reg4046)} : $signed($unsigned((8'hab))))))
                    begin
                      reg4180 <= reg4002[(4'he):(4'hc)];
                      reg4181 <= ((~|{$unsigned((8'ha2))}) ?
                          $signed(((-reg4134) && (&(8'hb6)))) : reg4060[(3'h6):(2'h2)]);
                      reg4182 <= reg4160;
                    end
                  else
                    begin
                      reg4180 <= ({reg4028[(2'h3):(2'h2)]} != (!(8'had)));
                      reg4181 <= reg4107;
                      reg4182 <= reg4008;
                      reg4183 <= $unsigned(wire3944[(1'h1):(1'h1)]);
                    end
                  if ($signed((&$unsigned((reg4131 ? (8'hb3) : reg4175)))))
                    begin
                      reg4184 <= reg3968[(2'h2):(1'h1)];
                      reg4185 <= reg4009;
                    end
                  else
                    begin
                      reg4184 <= (8'haa);
                      reg4185 <= (!reg4129[(2'h2):(2'h2)]);
                    end
                  for (forvar4186 = (1'h0); (forvar4186 < (1'h0)); forvar4186 = (forvar4186 + (1'h1)))
                    begin
                      reg4187 <= $signed((^reg3997));
                    end
                  if ($signed(reg4066[(3'h5):(1'h0)]))
                    begin
                      reg4188 <= (~|$unsigned({reg3987}));
                      reg4189 <= $signed((reg4177[(4'h8):(1'h1)] >>> ({(8'ha6)} & $unsigned(reg4163))));
                      reg4190 <= ($unsigned(($signed(reg4078) | (reg3960 != reg3974))) ?
                          $unsigned($signed((reg4105 ^~ reg4078))) : reg4009[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg4188 <= reg4077[(2'h3):(2'h2)];
                      reg4189 <= (((-reg4089[(3'h4):(1'h0)]) ?
                              {reg4136[(1'h0):(1'h0)]} : $signed(reg4076)) ?
                          (&(!$unsigned(wire3941))) : forvar4133[(4'h8):(2'h3)]);
                      reg4190 <= (+((^reg4131[(1'h0):(1'h0)]) ?
                          reg4131 : ($unsigned(reg3947) ?
                              {wire3941} : $signed(reg4045))));
                      reg4191 <= $unsigned((^forvar4170[(2'h3):(2'h2)]));
                    end
                end
            end
          else
            begin
              for (forvar4142 = (1'h0); (forvar4142 < (1'h0)); forvar4142 = (forvar4142 + (1'h1)))
                begin
                  if (wire3937)
                    begin
                      reg4143 <= $unsigned((($unsigned(reg3965) ?
                              (reg4041 != reg4069) : forvar4126) ?
                          ($signed((8'ha5)) - ((8'ha5) << reg4086)) : reg4069[(2'h3):(2'h3)]));
                      reg4144 <= $signed((~^{forvar4173[(2'h3):(1'h1)]}));
                    end
                  else
                    begin
                      reg4143 <= reg3950[(1'h0):(1'h0)];
                      reg4144 <= $signed(reg4067[(2'h2):(1'h0)]);
                      reg4145 <= (((^$unsigned(reg4018)) ?
                              $signed((forvar4144 ?
                                  (8'ha8) : reg4128)) : (+reg4069)) ?
                          (-reg4061) : reg4074);
                      reg4146 <= ({$signed($signed(reg3946))} ?
                          $unsigned(((+reg3995) << (-(8'hb5)))) : forvar4134);
                    end
                end
              if (($signed(($signed(reg3958) | (reg4167 | (8'hb4)))) ?
                  reg4037 : reg4133[(2'h2):(1'h0)]))
                begin
                  if (reg3997[(1'h1):(1'h0)])
                    begin
                      reg4147 <= ((($unsigned(reg4147) ?
                          (reg4110 < (8'hab)) : (reg4190 + reg3999)) != reg3964) + $unsigned(($signed(reg4132) ?
                          (8'haa) : reg4000)));
                      reg4148 <= $signed($unsigned((~^{reg4111})));
                    end
                  else
                    begin
                      reg4147 <= $unsigned(reg4190);
                      reg4148 <= $signed(($signed($signed(reg4151)) >>> {reg4129[(1'h1):(1'h0)]}));
                      reg4149 <= reg4084[(1'h1):(1'h1)];
                    end
                  if ($unsigned((reg3990[(2'h2):(2'h2)] ?
                      (~$unsigned(reg4095)) : ($signed((8'hb7)) ?
                          forvar4128[(2'h2):(1'h1)] : (reg4055 - (8'hac))))))
                    begin
                      reg4150 <= {((reg4111[(2'h3):(1'h0)] << $unsigned(reg4039)) ?
                              reg4176[(4'h8):(1'h0)] : {reg4087[(2'h3):(2'h2)]})};
                      reg4151 <= reg4092[(4'h9):(3'h4)];
                      reg4152 <= $unsigned($unsigned($unsigned((reg4006 >> reg4172))));
                      reg4153 <= reg4053;
                    end
                  else
                    begin
                      reg4150 <= forvar4135;
                      reg4151 <= reg4102;
                    end
                  if (reg4071)
                    begin
                      reg4154 <= reg4097;
                      reg4155 <= (^reg3955);
                      reg4156 <= (({(wire3938 ^~ reg4128)} ?
                          (8'ha3) : $signed((reg4182 << reg3996))) >>> reg4087[(3'h5):(1'h1)]);
                    end
                  else
                    begin
                      reg4154 <= (~&($signed((reg3977 | reg3964)) ?
                          ((+reg4064) != reg4165[(4'h8):(2'h3)]) : reg4164[(1'h1):(1'h1)]));
                    end
                end
              else
                begin
                  if (reg4045[(3'h4):(1'h0)])
                    begin
                      reg4147 <= $unsigned(($unsigned(reg4093[(1'h1):(1'h0)]) + ((|wire3938) ^ reg4145[(2'h3):(2'h3)])));
                      reg4148 <= (8'hac);
                      reg4149 <= reg4125;
                    end
                  else
                    begin
                      reg4147 <= (8'hba);
                      reg4148 <= (reg4158 ?
                          ((((8'ha6) | reg4191) - ((8'ha2) ?
                                  reg3994 : reg4033)) ?
                              ($signed((8'ha0)) <= (^forvar4126)) : $signed((~|reg4070))) : reg4117);
                      reg4149 <= (8'hae);
                      reg4150 <= (~$unsigned((8'h9c)));
                    end
                  reg4151 <= (wire3937[(1'h0):(1'h0)] > $signed((!forvar4186[(2'h2):(2'h2)])));
                  for (forvar4152 = (1'h0); (forvar4152 < (1'h1)); forvar4152 = (forvar4152 + (1'h1)))
                    begin
                      reg4153 <= forvar4179;
                      reg4154 <= (~$unsigned(wire3944[(1'h1):(1'h1)]));
                      reg4155 <= $unsigned($signed((~^(reg3956 ?
                          reg4176 : reg4054))));
                    end
                  if ($unsigned(reg4119[(2'h2):(1'h0)]))
                    begin
                      reg4156 <= reg4058[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg4156 <= reg4105;
                      reg4157 <= $signed(reg4155);
                    end
                end
              for (forvar4158 = (1'h0); (forvar4158 < (2'h3)); forvar4158 = (forvar4158 + (1'h1)))
                begin
                  reg4159 <= ($signed(reg4174) ?
                      (($unsigned(reg3968) ?
                          $signed(reg4053) : $unsigned(reg3974)) << ($unsigned(reg4143) ?
                          reg4068[(3'h4):(2'h2)] : ((8'ha6) ?
                              reg4174 : reg4056))) : reg4097[(3'h4):(3'h4)]);
                  for (forvar4160 = (1'h0); (forvar4160 < (1'h1)); forvar4160 = (forvar4160 + (1'h1)))
                    begin
                      reg4161 <= ((^reg4014[(3'h7):(2'h3)]) <<< {(+{reg4089})});
                    end
                end
            end
          for (forvar4192 = (1'h0); (forvar4192 < (1'h0)); forvar4192 = (forvar4192 + (1'h1)))
            begin
              if (forvar4133[(1'h1):(1'h0)])
                begin
                  reg4193 <= (^~reg4080[(3'h7):(2'h3)]);
                  for (forvar4194 = (1'h0); (forvar4194 < (1'h0)); forvar4194 = (forvar4194 + (1'h1)))
                    begin
                      reg4195 <= $unsigned($unsigned($unsigned((+reg4042))));
                      reg4196 <= $signed((8'hb4));
                    end
                end
              else
                begin
                  if ({reg4010})
                    begin
                      reg4193 <= reg4077;
                      reg4194 <= (wire3941 ?
                          $unsigned(reg3980) : $signed(reg4046));
                    end
                  else
                    begin
                      reg4193 <= reg3947[(2'h2):(1'h1)];
                      reg4194 <= ((reg4154 ?
                              $signed($signed(reg4178)) : ({reg3956} ~^ $unsigned(reg4048))) ?
                          (reg4057[(3'h4):(1'h0)] ^~ (reg4152[(3'h6):(1'h1)] ?
                              (reg4110 ?
                                  reg4129 : reg4075) : reg4115[(1'h1):(1'h0)])) : $signed({reg3957[(2'h2):(1'h0)]}));
                    end
                end
              for (forvar4197 = (1'h0); (forvar4197 < (2'h2)); forvar4197 = (forvar4197 + (1'h1)))
                begin
                  if ($signed(reg4095[(1'h0):(1'h0)]))
                    begin
                      reg4198 <= ($unsigned((~&{(8'ha0)})) ?
                          (^~(~^(reg4099 ? reg4161 : reg4116))) : reg3998);
                      reg4199 <= (8'hb7);
                    end
                  else
                    begin
                      reg4198 <= reg4148;
                      reg4199 <= (reg4048 <<< $signed((+(reg4027 & reg4075))));
                      reg4200 <= $unsigned((reg4177[(4'ha):(3'h5)] == ($unsigned(reg4011) >= $signed(reg4116))));
                    end
                end
              if (reg4194)
                begin
                  for (forvar4201 = (1'h0); (forvar4201 < (1'h1)); forvar4201 = (forvar4201 + (1'h1)))
                    begin
                      reg4202 <= (&reg4124[(1'h0):(1'h0)]);
                      reg4203 <= $signed(((reg4007 >= reg4090) ?
                          $unsigned($signed(reg3954)) : (-(reg4047 ?
                              reg4145 : (8'ha3)))));
                      reg4204 <= $signed((~|(!$unsigned((8'h9e)))));
                    end
                  for (forvar4205 = (1'h0); (forvar4205 < (2'h2)); forvar4205 = (forvar4205 + (1'h1)))
                    begin
                      reg4206 <= $unsigned($unsigned((~|{forvar4158})));
                    end
                end
              else
                begin
                  for (forvar4201 = (1'h0); (forvar4201 < (1'h0)); forvar4201 = (forvar4201 + (1'h1)))
                    begin
                      reg4202 <= (|($signed(reg3973[(4'h8):(4'h8)]) > reg4129[(4'he):(4'ha)]));
                      reg4203 <= (&$unsigned(((wire3940 || reg4019) ?
                          (forvar4186 <= reg4184) : $signed((8'h9e)))));
                    end
                  for (forvar4204 = (1'h0); (forvar4204 < (2'h2)); forvar4204 = (forvar4204 + (1'h1)))
                    begin
                      reg4205 <= $signed((~&$signed(forvar4128)));
                      reg4206 <= forvar4158[(2'h2):(1'h0)];
                      reg4207 <= forvar4179[(4'h9):(1'h1)];
                      reg4208 <= reg4104;
                    end
                  for (forvar4209 = (1'h0); (forvar4209 < (2'h2)); forvar4209 = (forvar4209 + (1'h1)))
                    begin
                      reg4210 <= $signed($unsigned(({reg3982} <<< $unsigned(reg4113))));
                    end
                  reg4211 <= {{reg4049}};
                end
            end
        end
      else
        begin
          reg4126 <= (-((|reg4084) ? reg4125 : ($unsigned(reg3960) - reg4049)));
        end
    end
  assign wire4212 = $unsigned(reg4091);
  assign wire4213 = ((wire3937 == (~^(reg4008 | reg4077))) >>> reg3951);
  module4214 #() modinst4534 (.clk(clk), .wire4216(reg4039), .y(wire4533), .wire4215(reg4176), .wire4218(reg3961), .wire4217(reg4148));
  assign wire4535 = (reg4200[(2'h3):(1'h0)] && reg4106);
  assign wire4536 = (reg3998 < (-$unsigned((reg4049 ? reg3961 : reg4045))));
  assign wire4537 = ($signed(reg3950[(1'h0):(1'h0)]) ?
                        reg4086 : {({reg4102} ~^ $signed((8'ha4)))});
  assign wire4538 = (&{$signed((-reg4165))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4214  (y, clk, wire4218, wire4217, wire4216, wire4215);
  output wire [(32'hd46):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire4218;
  input wire [(3'h6):(1'h0)] wire4217;
  input wire signed [(3'h6):(1'h0)] wire4216;
  input wire signed [(4'hf):(1'h0)] wire4215;
  wire [(3'h7):(1'h0)] wire4532;
  wire [(3'h5):(1'h0)] wire4430;
  wire [(4'ha):(1'h0)] wire4270;
  reg [(3'h7):(1'h0)] reg4531 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4530 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4528 = (1'h0);
  reg [(4'hd):(1'h0)] reg4527 = (1'h0);
  reg [(4'hd):(1'h0)] reg4526 = (1'h0);
  reg [(3'h5):(1'h0)] reg4525 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4524 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4523 = (1'h0);
  reg [(3'h5):(1'h0)] reg4522 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4521 = (1'h0);
  reg [(4'h9):(1'h0)] reg4514 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4519 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4518 = (1'h0);
  reg [(4'hb):(1'h0)] reg4517 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4516 = (1'h0);
  reg [(2'h2):(1'h0)] reg4515 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4513 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4512 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4511 = (1'h0);
  reg [(3'h5):(1'h0)] reg4507 = (1'h0);
  reg [(4'ha):(1'h0)] reg4504 = (1'h0);
  reg [(3'h7):(1'h0)] reg4501 = (1'h0);
  reg [(4'hb):(1'h0)] reg4500 = (1'h0);
  reg [(5'h10):(1'h0)] reg4510 = (1'h0);
  reg [(4'h8):(1'h0)] reg4509 = (1'h0);
  reg [(4'hc):(1'h0)] reg4508 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4506 = (1'h0);
  reg [(4'he):(1'h0)] reg4505 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4503 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4502 = (1'h0);
  reg [(3'h4):(1'h0)] reg4499 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4498 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4497 = (1'h0);
  reg [(4'h9):(1'h0)] reg4496 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4494 = (1'h0);
  reg [(5'h10):(1'h0)] reg4493 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4492 = (1'h0);
  reg [(3'h5):(1'h0)] reg4491 = (1'h0);
  reg [(4'hd):(1'h0)] reg4490 = (1'h0);
  reg [(4'hb):(1'h0)] reg4489 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4488 = (1'h0);
  reg [(5'h10):(1'h0)] reg4487 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4485 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4484 = (1'h0);
  reg [(4'h9):(1'h0)] reg4483 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4479 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4478 = (1'h0);
  reg [(4'ha):(1'h0)] reg4477 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4476 = (1'h0);
  reg [(4'ha):(1'h0)] reg4475 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4474 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4473 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4462 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4471 = (1'h0);
  reg [(4'hd):(1'h0)] reg4470 = (1'h0);
  reg [(3'h5):(1'h0)] reg4469 = (1'h0);
  reg [(2'h3):(1'h0)] reg4468 = (1'h0);
  reg [(5'h10):(1'h0)] reg4467 = (1'h0);
  reg [(4'h8):(1'h0)] reg4465 = (1'h0);
  reg [(3'h4):(1'h0)] reg4464 = (1'h0);
  reg [(3'h7):(1'h0)] reg4463 = (1'h0);
  reg [(3'h4):(1'h0)] reg4461 = (1'h0);
  reg [(5'h10):(1'h0)] reg4460 = (1'h0);
  reg [(4'hf):(1'h0)] reg4445 = (1'h0);
  reg [(4'hb):(1'h0)] reg4455 = (1'h0);
  reg [(4'hf):(1'h0)] reg4454 = (1'h0);
  reg [(4'h9):(1'h0)] reg4453 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4451 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4450 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4449 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4448 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4447 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4446 = (1'h0);
  reg [(5'h10):(1'h0)] reg4435 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4444 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4443 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4433 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4442 = (1'h0);
  reg [(4'ha):(1'h0)] reg4441 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4440 = (1'h0);
  reg [(4'ha):(1'h0)] reg4439 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4438 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4437 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4436 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4434 = (1'h0);
  reg [(2'h3):(1'h0)] reg4429 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4428 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4427 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4423 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4426 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4425 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4424 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4422 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4421 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4420 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4419 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4418 = (1'h0);
  reg [(4'ha):(1'h0)] reg4417 = (1'h0);
  reg [(4'hf):(1'h0)] reg4416 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4415 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4414 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4413 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4412 = (1'h0);
  reg [(4'hc):(1'h0)] reg4411 = (1'h0);
  reg [(4'h8):(1'h0)] reg4410 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4408 = (1'h0);
  reg [(2'h3):(1'h0)] reg4406 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4405 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4404 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4403 = (1'h0);
  reg [(3'h7):(1'h0)] reg4401 = (1'h0);
  reg [(3'h7):(1'h0)] reg4400 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4399 = (1'h0);
  reg [(3'h4):(1'h0)] reg4398 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4397 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4396 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4395 = (1'h0);
  reg [(4'ha):(1'h0)] reg4394 = (1'h0);
  reg [(4'h8):(1'h0)] reg4393 = (1'h0);
  reg [(3'h6):(1'h0)] reg4392 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4391 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4390 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4389 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4388 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4387 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4386 = (1'h0);
  reg [(4'he):(1'h0)] reg4385 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4384 = (1'h0);
  reg [(4'ha):(1'h0)] reg4383 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4380 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4379 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4378 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4377 = (1'h0);
  reg [(4'h9):(1'h0)] reg4373 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4367 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4364 = (1'h0);
  reg [(3'h6):(1'h0)] reg4362 = (1'h0);
  reg [(4'ha):(1'h0)] reg4376 = (1'h0);
  reg [(5'h10):(1'h0)] reg4375 = (1'h0);
  reg [(3'h7):(1'h0)] reg4374 = (1'h0);
  reg [(4'h8):(1'h0)] reg4372 = (1'h0);
  reg [(4'h8):(1'h0)] reg4371 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4370 = (1'h0);
  reg [(4'h9):(1'h0)] reg4369 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4368 = (1'h0);
  reg [(3'h6):(1'h0)] reg4360 = (1'h0);
  reg [(4'hb):(1'h0)] reg4366 = (1'h0);
  reg [(3'h7):(1'h0)] reg4365 = (1'h0);
  reg [(4'hb):(1'h0)] reg4363 = (1'h0);
  reg [(4'he):(1'h0)] reg4361 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4358 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4357 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4356 = (1'h0);
  reg [(4'hc):(1'h0)] reg4355 = (1'h0);
  reg [(4'h8):(1'h0)] reg4354 = (1'h0);
  reg [(4'hd):(1'h0)] reg4352 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4351 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4350 = (1'h0);
  reg [(4'h8):(1'h0)] reg4349 = (1'h0);
  reg [(4'ha):(1'h0)] reg4348 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4347 = (1'h0);
  reg [(5'h10):(1'h0)] reg4346 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4345 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4340 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4344 = (1'h0);
  reg [(4'he):(1'h0)] reg4343 = (1'h0);
  reg [(4'he):(1'h0)] reg4342 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4341 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4323 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4320 = (1'h0);
  reg [(4'ha):(1'h0)] reg4338 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4337 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4336 = (1'h0);
  reg [(2'h2):(1'h0)] reg4335 = (1'h0);
  reg [(4'h8):(1'h0)] reg4334 = (1'h0);
  reg [(4'ha):(1'h0)] reg4332 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4331 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4330 = (1'h0);
  reg [(2'h3):(1'h0)] reg4329 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4328 = (1'h0);
  reg [(4'hd):(1'h0)] reg4327 = (1'h0);
  reg [(4'hb):(1'h0)] reg4326 = (1'h0);
  reg [(3'h4):(1'h0)] reg4325 = (1'h0);
  reg [(4'hb):(1'h0)] reg4324 = (1'h0);
  reg [(4'he):(1'h0)] reg4322 = (1'h0);
  reg [(4'hc):(1'h0)] reg4321 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4319 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4318 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4317 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4316 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4315 = (1'h0);
  reg [(2'h2):(1'h0)] reg4314 = (1'h0);
  reg [(4'h8):(1'h0)] reg4313 = (1'h0);
  reg [(3'h7):(1'h0)] reg4312 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4311 = (1'h0);
  reg [(4'hf):(1'h0)] reg4310 = (1'h0);
  reg [(2'h3):(1'h0)] reg4309 = (1'h0);
  reg [(4'hf):(1'h0)] reg4308 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4307 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4306 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4305 = (1'h0);
  reg [(3'h5):(1'h0)] reg4304 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4302 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4300 = (1'h0);
  reg [(5'h10):(1'h0)] reg4299 = (1'h0);
  reg [(4'h8):(1'h0)] reg4298 = (1'h0);
  reg [(4'h9):(1'h0)] reg4297 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4296 = (1'h0);
  reg [(4'ha):(1'h0)] reg4295 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4294 = (1'h0);
  reg [(4'h9):(1'h0)] reg4292 = (1'h0);
  reg [(4'he):(1'h0)] reg4291 = (1'h0);
  reg [(3'h6):(1'h0)] reg4290 = (1'h0);
  reg [(3'h5):(1'h0)] reg4289 = (1'h0);
  reg [(4'hc):(1'h0)] reg4287 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4286 = (1'h0);
  reg [(4'ha):(1'h0)] reg4285 = (1'h0);
  reg [(4'he):(1'h0)] reg4284 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4283 = (1'h0);
  reg [(4'ha):(1'h0)] reg4282 = (1'h0);
  reg [(5'h10):(1'h0)] reg4281 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4279 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4278 = (1'h0);
  reg [(5'h10):(1'h0)] reg4276 = (1'h0);
  reg [(4'hb):(1'h0)] reg4275 = (1'h0);
  reg [(4'hc):(1'h0)] reg4274 = (1'h0);
  reg [(5'h10):(1'h0)] reg4269 = (1'h0);
  reg [(4'hd):(1'h0)] reg4268 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4267 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4266 = (1'h0);
  reg [(3'h7):(1'h0)] reg4264 = (1'h0);
  reg [(2'h3):(1'h0)] reg4263 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4262 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4257 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4253 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4245 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4261 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4260 = (1'h0);
  reg [(4'h8):(1'h0)] reg4259 = (1'h0);
  reg [(4'h9):(1'h0)] reg4256 = (1'h0);
  reg [(4'hb):(1'h0)] reg4255 = (1'h0);
  reg [(3'h5):(1'h0)] reg4254 = (1'h0);
  reg [(4'he):(1'h0)] reg4252 = (1'h0);
  reg [(2'h3):(1'h0)] reg4251 = (1'h0);
  reg [(4'hd):(1'h0)] reg4250 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4249 = (1'h0);
  reg [(4'hc):(1'h0)] reg4247 = (1'h0);
  reg [(4'ha):(1'h0)] reg4248 = (1'h0);
  reg [(4'hf):(1'h0)] reg4246 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4243 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4242 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4234 = (1'h0);
  reg [(3'h4):(1'h0)] reg4229 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4222 = (1'h0);
  reg [(4'hf):(1'h0)] reg4241 = (1'h0);
  reg [(4'hb):(1'h0)] reg4240 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4239 = (1'h0);
  reg [(2'h2):(1'h0)] reg4238 = (1'h0);
  reg [(4'ha):(1'h0)] reg4237 = (1'h0);
  reg [(4'ha):(1'h0)] reg4236 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4235 = (1'h0);
  reg [(4'ha):(1'h0)] reg4233 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4232 = (1'h0);
  reg [(3'h5):(1'h0)] reg4231 = (1'h0);
  reg [(3'h4):(1'h0)] reg4228 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4227 = (1'h0);
  reg [(3'h6):(1'h0)] reg4226 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4225 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4224 = (1'h0);
  reg [(4'h9):(1'h0)] reg4223 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4219 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4529 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4520 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4514 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4510 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4506 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4507 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4504 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4501 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4500 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4495 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4487 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4488 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4486 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4482 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4481 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4480 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4476 = (1'h0);
  reg [(4'he):(1'h0)] forvar4473 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4472 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4466 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4462 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4459 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4458 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4457 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4456 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4442 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4440 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4439 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4437 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4436 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4449 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4452 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4445 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4441 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4435 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4433 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4432 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4431 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4422 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4423 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4409 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4407 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4402 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4401 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4396 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4393 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4382 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4381 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4376 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4371 = (1'h0);
  reg [(4'he):(1'h0)] forvar4370 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4363 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4373 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4367 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4364 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4362 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4360 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4359 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4353 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4343 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4340 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4339 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4325 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4321 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4312 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4307 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4333 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4323 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4320 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4313 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4306 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4303 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4301 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4293 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4288 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4280 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4277 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4273 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4272 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4271 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4265 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4260 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4255 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4251 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4246 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4258 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4257 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4253 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4248 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4247 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4245 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4244 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4235 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4228 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4227 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4234 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4230 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4229 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4222 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4221 = (1'h0);
  reg [(4'he):(1'h0)] forvar4220 = (1'h0);
  assign y = {wire4532,
                 wire4430,
                 wire4270,
                 reg4531,
                 reg4530,
                 reg4528,
                 reg4527,
                 reg4526,
                 reg4525,
                 reg4524,
                 reg4523,
                 reg4522,
                 reg4521,
                 reg4514,
                 reg4519,
                 reg4518,
                 reg4517,
                 reg4516,
                 reg4515,
                 reg4513,
                 reg4512,
                 reg4511,
                 reg4507,
                 reg4504,
                 reg4501,
                 reg4500,
                 reg4510,
                 reg4509,
                 reg4508,
                 reg4506,
                 reg4505,
                 reg4503,
                 reg4502,
                 reg4499,
                 reg4498,
                 reg4497,
                 reg4496,
                 reg4494,
                 reg4493,
                 reg4492,
                 reg4491,
                 reg4490,
                 reg4489,
                 reg4488,
                 reg4487,
                 reg4485,
                 reg4484,
                 reg4483,
                 reg4479,
                 reg4478,
                 reg4477,
                 reg4476,
                 reg4475,
                 reg4474,
                 reg4473,
                 reg4462,
                 reg4471,
                 reg4470,
                 reg4469,
                 reg4468,
                 reg4467,
                 reg4465,
                 reg4464,
                 reg4463,
                 reg4461,
                 reg4460,
                 reg4445,
                 reg4455,
                 reg4454,
                 reg4453,
                 reg4451,
                 reg4450,
                 reg4449,
                 reg4448,
                 reg4447,
                 reg4446,
                 reg4435,
                 reg4444,
                 reg4443,
                 reg4433,
                 reg4442,
                 reg4441,
                 reg4440,
                 reg4439,
                 reg4438,
                 reg4437,
                 reg4436,
                 reg4434,
                 reg4429,
                 reg4428,
                 reg4427,
                 reg4423,
                 reg4426,
                 reg4425,
                 reg4424,
                 reg4422,
                 reg4421,
                 reg4420,
                 reg4419,
                 reg4418,
                 reg4417,
                 reg4416,
                 reg4415,
                 reg4414,
                 reg4413,
                 reg4412,
                 reg4411,
                 reg4410,
                 reg4408,
                 reg4406,
                 reg4405,
                 reg4404,
                 reg4403,
                 reg4401,
                 reg4400,
                 reg4399,
                 reg4398,
                 reg4397,
                 reg4396,
                 reg4395,
                 reg4394,
                 reg4393,
                 reg4392,
                 reg4391,
                 reg4390,
                 reg4389,
                 reg4388,
                 reg4387,
                 reg4386,
                 reg4385,
                 reg4384,
                 reg4383,
                 reg4380,
                 reg4379,
                 reg4378,
                 reg4377,
                 reg4373,
                 reg4367,
                 reg4364,
                 reg4362,
                 reg4376,
                 reg4375,
                 reg4374,
                 reg4372,
                 reg4371,
                 reg4370,
                 reg4369,
                 reg4368,
                 reg4360,
                 reg4366,
                 reg4365,
                 reg4363,
                 reg4361,
                 reg4358,
                 reg4357,
                 reg4356,
                 reg4355,
                 reg4354,
                 reg4352,
                 reg4351,
                 reg4350,
                 reg4349,
                 reg4348,
                 reg4347,
                 reg4346,
                 reg4345,
                 reg4340,
                 reg4344,
                 reg4343,
                 reg4342,
                 reg4341,
                 reg4323,
                 reg4320,
                 reg4338,
                 reg4337,
                 reg4336,
                 reg4335,
                 reg4334,
                 reg4332,
                 reg4331,
                 reg4330,
                 reg4329,
                 reg4328,
                 reg4327,
                 reg4326,
                 reg4325,
                 reg4324,
                 reg4322,
                 reg4321,
                 reg4319,
                 reg4318,
                 reg4317,
                 reg4316,
                 reg4315,
                 reg4314,
                 reg4313,
                 reg4312,
                 reg4311,
                 reg4310,
                 reg4309,
                 reg4308,
                 reg4307,
                 reg4306,
                 reg4305,
                 reg4304,
                 reg4302,
                 reg4300,
                 reg4299,
                 reg4298,
                 reg4297,
                 reg4296,
                 reg4295,
                 reg4294,
                 reg4292,
                 reg4291,
                 reg4290,
                 reg4289,
                 reg4287,
                 reg4286,
                 reg4285,
                 reg4284,
                 reg4283,
                 reg4282,
                 reg4281,
                 reg4279,
                 reg4278,
                 reg4276,
                 reg4275,
                 reg4274,
                 reg4269,
                 reg4268,
                 reg4267,
                 reg4266,
                 reg4264,
                 reg4263,
                 reg4262,
                 reg4258,
                 reg4257,
                 reg4253,
                 reg4245,
                 reg4261,
                 reg4260,
                 reg4259,
                 reg4256,
                 reg4255,
                 reg4254,
                 reg4252,
                 reg4251,
                 reg4250,
                 reg4249,
                 reg4247,
                 reg4248,
                 reg4246,
                 reg4243,
                 reg4242,
                 reg4234,
                 reg4229,
                 reg4222,
                 reg4241,
                 reg4240,
                 reg4239,
                 reg4238,
                 reg4237,
                 reg4236,
                 reg4235,
                 reg4233,
                 reg4232,
                 reg4231,
                 reg4228,
                 reg4227,
                 reg4226,
                 reg4225,
                 reg4224,
                 reg4223,
                 reg4219,
                 forvar4529,
                 forvar4520,
                 forvar4514,
                 forvar4510,
                 forvar4506,
                 forvar4507,
                 forvar4504,
                 forvar4501,
                 forvar4500,
                 forvar4495,
                 forvar4487,
                 forvar4488,
                 forvar4486,
                 forvar4482,
                 forvar4481,
                 forvar4480,
                 forvar4476,
                 forvar4473,
                 forvar4472,
                 forvar4466,
                 forvar4462,
                 forvar4459,
                 forvar4458,
                 forvar4457,
                 forvar4456,
                 forvar4442,
                 forvar4440,
                 forvar4439,
                 forvar4437,
                 forvar4436,
                 forvar4449,
                 forvar4452,
                 forvar4445,
                 forvar4441,
                 forvar4435,
                 forvar4433,
                 forvar4432,
                 forvar4431,
                 forvar4422,
                 forvar4423,
                 forvar4409,
                 forvar4407,
                 forvar4402,
                 forvar4401,
                 forvar4396,
                 forvar4393,
                 forvar4382,
                 forvar4381,
                 forvar4376,
                 forvar4371,
                 forvar4370,
                 forvar4363,
                 forvar4373,
                 forvar4367,
                 forvar4364,
                 forvar4362,
                 forvar4360,
                 forvar4359,
                 forvar4353,
                 forvar4343,
                 forvar4340,
                 forvar4339,
                 forvar4325,
                 forvar4321,
                 forvar4312,
                 forvar4307,
                 forvar4333,
                 forvar4323,
                 forvar4320,
                 forvar4313,
                 forvar4306,
                 forvar4303,
                 forvar4301,
                 forvar4293,
                 forvar4288,
                 forvar4280,
                 forvar4277,
                 forvar4273,
                 forvar4272,
                 forvar4271,
                 forvar4265,
                 forvar4260,
                 forvar4255,
                 forvar4251,
                 forvar4246,
                 forvar4258,
                 forvar4257,
                 forvar4253,
                 forvar4248,
                 forvar4247,
                 forvar4245,
                 forvar4244,
                 forvar4235,
                 forvar4228,
                 forvar4227,
                 forvar4234,
                 forvar4230,
                 forvar4229,
                 forvar4222,
                 forvar4221,
                 forvar4220,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4219 <= {($unsigned($signed(wire4215)) ?
              wire4217 : (wire4215[(1'h1):(1'h0)] <= $unsigned(wire4216)))};
      for (forvar4220 = (1'h0); (forvar4220 < (1'h1)); forvar4220 = (forvar4220 + (1'h1)))
        begin
          if ((wire4218 && (-forvar4220)))
            begin
              for (forvar4221 = (1'h0); (forvar4221 < (2'h2)); forvar4221 = (forvar4221 + (1'h1)))
                begin
                  for (forvar4222 = (1'h0); (forvar4222 < (1'h1)); forvar4222 = (forvar4222 + (1'h1)))
                    begin
                      reg4223 <= (wire4218[(3'h7):(3'h7)] ?
                          ({$unsigned(wire4215)} * wire4217[(2'h3):(2'h3)]) : wire4215);
                      reg4224 <= wire4216[(3'h5):(1'h0)];
                      reg4225 <= (~reg4223);
                      reg4226 <= ($signed($unsigned(((8'hb9) ?
                          reg4225 : reg4224))) && (&$signed(wire4217[(2'h2):(2'h2)])));
                    end
                  if (wire4216)
                    begin
                      reg4227 <= (+wire4217[(2'h2):(1'h0)]);
                      reg4228 <= (&(&(reg4224[(1'h0):(1'h0)] ?
                          wire4215[(3'h7):(3'h7)] : (reg4223 & wire4216))));
                    end
                  else
                    begin
                      reg4227 <= (~wire4216[(3'h5):(2'h2)]);
                      reg4228 <= $signed((|reg4227[(3'h4):(2'h2)]));
                    end
                end
              for (forvar4229 = (1'h0); (forvar4229 < (2'h3)); forvar4229 = (forvar4229 + (1'h1)))
                begin
                  for (forvar4230 = (1'h0); (forvar4230 < (2'h2)); forvar4230 = (forvar4230 + (1'h1)))
                    begin
                      reg4231 <= $unsigned((({reg4219} == (|(8'ha3))) ?
                          reg4224 : (forvar4230[(3'h5):(3'h4)] ?
                              (wire4216 << reg4226) : reg4227[(2'h2):(1'h1)])));
                      reg4232 <= {reg4223};
                      reg4233 <= $unsigned(reg4219);
                    end
                  for (forvar4234 = (1'h0); (forvar4234 < (2'h3)); forvar4234 = (forvar4234 + (1'h1)))
                    begin
                      reg4235 <= reg4231;
                      reg4236 <= wire4216;
                      reg4237 <= ($unsigned(forvar4229) ?
                          (+$signed(reg4226)) : wire4217[(1'h0):(1'h0)]);
                    end
                  reg4238 <= $unsigned(forvar4234);
                  if ((-reg4237[(4'h8):(3'h4)]))
                    begin
                      reg4239 <= ($signed(forvar4222[(3'h5):(3'h5)]) ?
                          (!$signed($unsigned((8'hb4)))) : {(8'ha0)});
                      reg4240 <= reg4228;
                      reg4241 <= $signed(reg4236[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg4239 <= $unsigned((reg4225[(1'h0):(1'h0)] ?
                          $unsigned(reg4224[(1'h1):(1'h0)]) : $unsigned((&forvar4234))));
                      reg4240 <= forvar4230;
                    end
                end
            end
          else
            begin
              for (forvar4221 = (1'h0); (forvar4221 < (1'h0)); forvar4221 = (forvar4221 + (1'h1)))
                begin
                  if ($signed(reg4238[(1'h1):(1'h1)]))
                    begin
                      reg4222 <= reg4226;
                      reg4223 <= (({$unsigned(reg4226)} ? (8'h9f) : wire4218) ?
                          $unsigned(((reg4228 << reg4228) == {forvar4220})) : reg4241);
                      reg4224 <= ((reg4219[(4'ha):(1'h0)] ^~ {(^reg4232)}) ?
                          (^~{reg4219[(4'hf):(3'h6)]}) : ((forvar4229[(3'h5):(1'h0)] ?
                                  $signed(reg4219) : $unsigned(reg4240)) ?
                              ($unsigned(reg4228) & reg4239) : $signed((reg4239 ?
                                  forvar4222 : wire4218))));
                    end
                  else
                    begin
                      reg4222 <= (^~$signed({$unsigned(wire4218)}));
                    end
                  if ($unsigned((8'ha0)))
                    begin
                      reg4225 <= (((8'haf) & {reg4227}) ?
                          $unsigned((~&reg4223)) : $unsigned($signed(reg4224[(2'h2):(1'h0)])));
                      reg4226 <= ((($signed(wire4217) ?
                          reg4240[(2'h2):(1'h0)] : (reg4222 >>> wire4215)) ~^ reg4235[(3'h7):(3'h6)]) - ((&(reg4235 ~^ reg4219)) - $signed((~^reg4227))));
                    end
                  else
                    begin
                      reg4225 <= $signed(($signed(reg4241) != (wire4216 <= (reg4219 <<< wire4215))));
                      reg4226 <= (~|{$signed(reg4232[(1'h0):(1'h0)])});
                    end
                end
              for (forvar4227 = (1'h0); (forvar4227 < (1'h0)); forvar4227 = (forvar4227 + (1'h1)))
                begin
                  for (forvar4228 = (1'h0); (forvar4228 < (1'h0)); forvar4228 = (forvar4228 + (1'h1)))
                    begin
                      reg4229 <= ((forvar4221[(1'h1):(1'h0)] ?
                          ($signed(reg4223) <<< (reg4235 ?
                              wire4217 : reg4235)) : (+$signed((8'hb0)))) && (wire4217 ^~ $unsigned($unsigned(forvar4229))));
                    end
                  for (forvar4230 = (1'h0); (forvar4230 < (1'h1)); forvar4230 = (forvar4230 + (1'h1)))
                    begin
                      reg4231 <= $signed(reg4239[(3'h4):(2'h2)]);
                      reg4232 <= (-(^$unsigned($unsigned(reg4227))));
                      reg4233 <= forvar4228[(3'h4):(1'h0)];
                    end
                end
              if ($signed(((~wire4215[(4'ha):(3'h5)]) != (~reg4219[(1'h0):(1'h0)]))))
                begin
                  reg4234 <= reg4228;
                  for (forvar4235 = (1'h0); (forvar4235 < (1'h0)); forvar4235 = (forvar4235 + (1'h1)))
                    begin
                      reg4236 <= $signed({($unsigned((8'hb2)) >= {wire4216})});
                      reg4237 <= reg4241[(4'hf):(4'hd)];
                      reg4238 <= $unsigned((|((|reg4241) ?
                          $unsigned((8'hb8)) : ((8'h9c) >= reg4231))));
                      reg4239 <= ($unsigned(reg4231[(3'h4):(2'h3)]) ?
                          $signed($unsigned((^~reg4229))) : (({(8'ha1)} ^ reg4233[(4'h8):(3'h7)]) && $unsigned((forvar4234 > forvar4220))));
                    end
                end
              else
                begin
                  if (forvar4230)
                    begin
                      reg4234 <= (^~$unsigned($unsigned(wire4215)));
                      reg4235 <= (!(wire4215 ^ $unsigned((wire4216 || reg4222))));
                    end
                  else
                    begin
                      reg4234 <= $unsigned($unsigned((^$unsigned(reg4240))));
                      reg4235 <= ($signed($unsigned((reg4227 ?
                              reg4237 : reg4233))) ?
                          reg4234 : reg4236[(3'h5):(3'h5)]);
                      reg4236 <= (+$unsigned($unsigned(reg4224[(1'h1):(1'h1)])));
                    end
                  if (($signed(((reg4232 || reg4236) ?
                          reg4240[(2'h3):(1'h0)] : (wire4216 > reg4239))) ?
                      {{(forvar4227 ?
                                  wire4217 : wire4217)}} : $signed($signed(reg4241))))
                    begin
                      reg4237 <= (-$signed((forvar4220[(1'h0):(1'h0)] != {reg4239})));
                    end
                  else
                    begin
                      reg4237 <= reg4231;
                    end
                  if ({reg4227})
                    begin
                      reg4238 <= (~&(^~$unsigned(reg4232)));
                    end
                  else
                    begin
                      reg4238 <= (reg4235[(2'h2):(2'h2)] ?
                          ((|$unsigned((8'hb4))) ?
                              reg4241[(4'hd):(2'h2)] : $signed(forvar4221)) : ({reg4238} < (((8'ha1) >> forvar4221) != {forvar4227})));
                      reg4239 <= ((({reg4229} ?
                              $signed(reg4239) : (reg4223 ?
                                  reg4237 : forvar4221)) ?
                          $unsigned((wire4216 ?
                              wire4215 : wire4215)) : (|(~(8'h9c)))) >= reg4223[(4'h9):(1'h1)]);
                    end
                end
            end
          reg4242 <= forvar4221;
          reg4243 <= {$unsigned($unsigned($signed(reg4241)))};
        end
      for (forvar4244 = (1'h0); (forvar4244 < (1'h1)); forvar4244 = (forvar4244 + (1'h1)))
        begin
          if (reg4225)
            begin
              if ((!reg4227))
                begin
                  for (forvar4245 = (1'h0); (forvar4245 < (2'h3)); forvar4245 = (forvar4245 + (1'h1)))
                    begin
                      reg4246 <= $signed($signed(((forvar4222 < forvar4227) ~^ (8'hb0))));
                    end
                  for (forvar4247 = (1'h0); (forvar4247 < (1'h1)); forvar4247 = (forvar4247 + (1'h1)))
                    begin
                      reg4248 <= {$signed(((forvar4244 ?
                              forvar4221 : forvar4245) - $unsigned(reg4231)))};
                    end
                end
              else
                begin
                  for (forvar4245 = (1'h0); (forvar4245 < (2'h2)); forvar4245 = (forvar4245 + (1'h1)))
                    begin
                      reg4246 <= forvar4245[(2'h3):(2'h2)];
                      reg4247 <= ((~^{$unsigned(wire4216)}) && $unsigned($signed((+forvar4221))));
                    end
                  for (forvar4248 = (1'h0); (forvar4248 < (2'h2)); forvar4248 = (forvar4248 + (1'h1)))
                    begin
                      reg4249 <= forvar4228[(3'h5):(3'h5)];
                      reg4250 <= ($signed($unsigned({reg4240})) ?
                          ({(~^forvar4228)} ?
                              $unsigned((reg4225 >= forvar4227)) : $signed((reg4247 ?
                                  (8'ha4) : reg4247))) : $unsigned(($signed(reg4219) > forvar4235)));
                      reg4251 <= $unsigned(reg4234);
                    end
                  reg4252 <= $signed((!reg4246));
                  for (forvar4253 = (1'h0); (forvar4253 < (1'h0)); forvar4253 = (forvar4253 + (1'h1)))
                    begin
                      reg4254 <= forvar4230[(3'h6):(1'h0)];
                      reg4255 <= (+$signed(forvar4235[(3'h6):(3'h6)]));
                      reg4256 <= (~({$signed((8'hb9))} ^ (8'ha6)));
                    end
                end
              for (forvar4257 = (1'h0); (forvar4257 < (1'h1)); forvar4257 = (forvar4257 + (1'h1)))
                begin
                  for (forvar4258 = (1'h0); (forvar4258 < (1'h0)); forvar4258 = (forvar4258 + (1'h1)))
                    begin
                      reg4259 <= reg4249;
                      reg4260 <= reg4251[(2'h2):(2'h2)];
                      reg4261 <= $signed(((reg4254[(2'h3):(1'h0)] >>> (~&reg4231)) ?
                          $signed({(8'hba)}) : $signed(reg4227)));
                    end
                end
            end
          else
            begin
              reg4245 <= {reg4250[(3'h5):(2'h3)]};
              for (forvar4246 = (1'h0); (forvar4246 < (2'h3)); forvar4246 = (forvar4246 + (1'h1)))
                begin
                  if ((+$signed(forvar4229[(3'h4):(2'h3)])))
                    begin
                      reg4247 <= $signed(reg4255);
                    end
                  else
                    begin
                      reg4247 <= (((+(wire4216 && reg4251)) > (~|$unsigned((8'haa)))) ^~ ({wire4216[(1'h0):(1'h0)]} != $signed($signed((8'hb1)))));
                    end
                  if (($unsigned($signed((~&reg4245))) >> (&forvar4257)))
                    begin
                      reg4248 <= (8'ha5);
                      reg4249 <= (8'ha7);
                    end
                  else
                    begin
                      reg4248 <= ((^($signed(forvar4230) + $signed(reg4240))) ?
                          ($signed({forvar4247}) ?
                              ($unsigned(reg4241) ?
                                  {reg4229} : reg4240[(4'h9):(1'h0)]) : $unsigned($unsigned((8'ha8)))) : reg4223[(1'h0):(1'h0)]);
                      reg4249 <= (~&(8'hac));
                      reg4250 <= ((($unsigned(reg4240) ?
                              $unsigned(forvar4258) : (~reg4228)) ?
                          ((!reg4225) ?
                              {reg4238} : forvar4245) : $signed((|forvar4221))) > (reg4241 ?
                          forvar4222 : ((|reg4238) ?
                              forvar4248[(4'hb):(2'h3)] : $unsigned((8'ha2)))));
                    end
                  for (forvar4251 = (1'h0); (forvar4251 < (1'h0)); forvar4251 = (forvar4251 + (1'h1)))
                    begin
                      reg4252 <= (8'hb4);
                      reg4253 <= (~|reg4243);
                    end
                  reg4254 <= $signed($unsigned((+$unsigned(reg4246))));
                end
              if ($unsigned($signed((^(^reg4219)))))
                begin
                  for (forvar4255 = (1'h0); (forvar4255 < (2'h3)); forvar4255 = (forvar4255 + (1'h1)))
                    begin
                      reg4256 <= $unsigned(forvar4221[(3'h5):(2'h2)]);
                      reg4257 <= ((^~reg4239[(1'h1):(1'h0)]) ?
                          $signed(((forvar4222 ?
                              (8'ha3) : reg4233) < (reg4248 >>> wire4218))) : (forvar4244[(4'hd):(1'h0)] - ({(8'ha1)} ?
                              reg4225[(2'h2):(2'h2)] : (reg4229 ?
                                  reg4222 : reg4248))));
                      reg4258 <= {forvar4253[(3'h4):(2'h3)]};
                      reg4259 <= (({forvar4227} > ((~^forvar4255) & (reg4243 < forvar4246))) ?
                          $signed($unsigned($unsigned(reg4257))) : $signed((reg4255 ?
                              ((8'ha3) <<< forvar4230) : reg4242[(1'h0):(1'h0)])));
                    end
                  for (forvar4260 = (1'h0); (forvar4260 < (1'h0)); forvar4260 = (forvar4260 + (1'h1)))
                    begin
                      reg4261 <= ($signed(forvar4251[(2'h2):(1'h0)]) + $signed(($signed(reg4261) ?
                          {reg4237} : (wire4216 < reg4242))));
                      reg4262 <= {(~$signed(((8'hb5) ? reg4238 : reg4253)))};
                      reg4263 <= forvar4221[(1'h1):(1'h0)];
                      reg4264 <= ($unsigned((wire4217 ?
                              {(8'had)} : forvar4227)) ?
                          $signed(({reg4258} || reg4261)) : (8'ha3));
                    end
                  for (forvar4265 = (1'h0); (forvar4265 < (2'h2)); forvar4265 = (forvar4265 + (1'h1)))
                    begin
                      reg4266 <= (|$unsigned(forvar4258[(1'h1):(1'h0)]));
                      reg4267 <= (~^(8'hb4));
                      reg4268 <= $signed(forvar4234[(3'h7):(2'h2)]);
                      reg4269 <= reg4250;
                    end
                end
              else
                begin
                  reg4255 <= {$signed(reg4226[(1'h1):(1'h1)])};
                  reg4256 <= $unsigned($unsigned(reg4259));
                end
            end
        end
    end
  assign wire4270 = ((((reg4229 || reg4249) ?
                        (&reg4250) : {reg4248}) ^~ $signed($signed(reg4263))) * $signed($signed((8'hb2))));
  always
    @(posedge clk) begin
      for (forvar4271 = (1'h0); (forvar4271 < (2'h3)); forvar4271 = (forvar4271 + (1'h1)))
        begin
          for (forvar4272 = (1'h0); (forvar4272 < (2'h2)); forvar4272 = (forvar4272 + (1'h1)))
            begin
              for (forvar4273 = (1'h0); (forvar4273 < (1'h0)); forvar4273 = (forvar4273 + (1'h1)))
                begin
                  if (reg4254[(3'h5):(1'h1)])
                    begin
                      reg4274 <= wire4217[(1'h1):(1'h1)];
                      reg4275 <= {$unsigned($unsigned($signed((8'h9d))))};
                      reg4276 <= ((((reg4267 ^ forvar4273) > {reg4269}) >= reg4263[(1'h0):(1'h0)]) - $signed(reg4232));
                    end
                  else
                    begin
                      reg4274 <= reg4248[(4'h8):(4'h8)];
                      reg4275 <= reg4262[(1'h1):(1'h0)];
                      reg4276 <= $unsigned($signed((~^(reg4276 && reg4275))));
                    end
                  for (forvar4277 = (1'h0); (forvar4277 < (2'h3)); forvar4277 = (forvar4277 + (1'h1)))
                    begin
                      reg4278 <= (reg4243[(2'h2):(2'h2)] ?
                          $signed($signed(reg4264)) : {{$unsigned(reg4249)}});
                      reg4279 <= reg4260[(2'h2):(1'h0)];
                    end
                  for (forvar4280 = (1'h0); (forvar4280 < (1'h1)); forvar4280 = (forvar4280 + (1'h1)))
                    begin
                      reg4281 <= $signed(reg4254[(3'h4):(1'h0)]);
                      reg4282 <= $signed(reg4226[(1'h0):(1'h0)]);
                      reg4283 <= $unsigned(reg4266[(2'h2):(1'h0)]);
                    end
                  if ($signed({(~&$signed(reg4253))}))
                    begin
                      reg4284 <= ($unsigned({(~&wire4270)}) ?
                          $unsigned($unsigned($unsigned(reg4258))) : reg4239[(3'h6):(1'h0)]);
                    end
                  else
                    begin
                      reg4284 <= reg4222[(2'h3):(1'h1)];
                      reg4285 <= reg4243;
                      reg4286 <= (^~(($unsigned(reg4283) | forvar4277) > forvar4271));
                      reg4287 <= ($unsigned($signed((forvar4277 <<< wire4215))) * (-$signed(reg4255)));
                    end
                end
              for (forvar4288 = (1'h0); (forvar4288 < (1'h0)); forvar4288 = (forvar4288 + (1'h1)))
                begin
                  if ($unsigned(reg4237))
                    begin
                      reg4289 <= (reg4253 ?
                          reg4262[(4'h9):(4'h8)] : ($signed(forvar4277) ?
                              ((reg4243 >= reg4243) ?
                                  $signed((8'h9f)) : $signed(reg4274)) : $unsigned((~&forvar4288))));
                      reg4290 <= $signed((({reg4246} ?
                          {(8'hae)} : {reg4240}) >= reg4251));
                    end
                  else
                    begin
                      reg4289 <= reg4255;
                      reg4290 <= {(|($unsigned(reg4274) ?
                              (reg4252 ? (8'hab) : reg4263) : {forvar4288}))};
                      reg4291 <= {{{((8'h9d) ? reg4249 : reg4283)}}};
                      reg4292 <= $unsigned(((reg4253 ?
                          reg4255[(2'h2):(1'h1)] : $signed(reg4246)) ^~ reg4268[(4'hb):(3'h7)]));
                    end
                  for (forvar4293 = (1'h0); (forvar4293 < (2'h2)); forvar4293 = (forvar4293 + (1'h1)))
                    begin
                      reg4294 <= reg4266[(2'h2):(2'h2)];
                      reg4295 <= $unsigned(((reg4285 ?
                          (reg4260 ? (8'hab) : reg4253) : (forvar4273 ?
                              reg4245 : (8'ha3))) != reg4235));
                      reg4296 <= (^~(+((reg4275 <= reg4231) ?
                          wire4217 : $signed((8'hb9)))));
                    end
                  if ((wire4215 ^~ reg4227))
                    begin
                      reg4297 <= ($unsigned(((~&reg4236) ?
                              (reg4251 ?
                                  forvar4273 : reg4274) : $unsigned(wire4216))) ?
                          reg4249[(2'h3):(2'h3)] : (forvar4280 ?
                              $unsigned(forvar4280) : ($signed(reg4295) ?
                                  reg4263[(1'h1):(1'h1)] : (~&reg4295))));
                    end
                  else
                    begin
                      reg4297 <= reg4242[(4'h9):(1'h0)];
                      reg4298 <= $unsigned($unsigned((!reg4219)));
                      reg4299 <= $unsigned(($signed(forvar4272[(2'h2):(2'h2)]) <<< (8'hb9)));
                      reg4300 <= $unsigned((^$signed(reg4296[(3'h6):(2'h3)])));
                    end
                end
              for (forvar4301 = (1'h0); (forvar4301 < (1'h0)); forvar4301 = (forvar4301 + (1'h1)))
                begin
                  reg4302 <= (($unsigned(forvar4277[(1'h1):(1'h1)]) > $signed((reg4255 ?
                          wire4218 : forvar4293))) ?
                      reg4228[(1'h1):(1'h1)] : reg4233);
                  for (forvar4303 = (1'h0); (forvar4303 < (1'h1)); forvar4303 = (forvar4303 + (1'h1)))
                    begin
                      reg4304 <= (~^(^~reg4297));
                      reg4305 <= {forvar4280};
                    end
                end
            end
          if ({$signed(reg4243)})
            begin
              if ($signed({(8'h9d)}))
                begin
                  if (forvar4288)
                    begin
                      reg4306 <= {forvar4303[(2'h3):(1'h1)]};
                      reg4307 <= reg4290[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg4306 <= reg4304[(3'h4):(2'h2)];
                      reg4307 <= $unsigned($signed(({reg4274} || $signed((8'ha3)))));
                      reg4308 <= reg4258;
                      reg4309 <= (+(8'hb6));
                    end
                end
              else
                begin
                  for (forvar4306 = (1'h0); (forvar4306 < (2'h3)); forvar4306 = (forvar4306 + (1'h1)))
                    begin
                      reg4307 <= $signed((((reg4243 & reg4267) ?
                              reg4219[(4'hd):(4'hc)] : $signed(reg4219)) ?
                          (reg4237[(4'h8):(4'h8)] & $signed(reg4247)) : reg4257));
                      reg4308 <= $unsigned(reg4260);
                      reg4309 <= (^($unsigned($signed(forvar4277)) * ($unsigned(reg4245) ?
                          {wire4215} : $signed(reg4269))));
                    end
                end
              if ($unsigned(reg4250))
                begin
                  if ($unsigned(reg4250[(3'h7):(3'h6)]))
                    begin
                      reg4310 <= reg4290[(3'h5):(1'h1)];
                      reg4311 <= reg4225;
                      reg4312 <= (reg4269 ? {(|$signed(reg4294))} : reg4232);
                    end
                  else
                    begin
                      reg4310 <= ({(reg4253 ?
                              (wire4215 ? forvar4288 : reg4260) : (reg4246 ?
                                  (8'hae) : reg4310))} ^ reg4219[(4'h9):(3'h6)]);
                      reg4311 <= reg4226;
                      reg4312 <= reg4264[(2'h3):(1'h0)];
                      reg4313 <= ($unsigned(reg4253[(1'h0):(1'h0)]) && {reg4242});
                    end
                  if ($unsigned((((reg4307 * reg4257) ? (8'hac) : (&reg4292)) ?
                      (~&$unsigned(reg4242)) : ((~|forvar4293) >> $unsigned(reg4312)))))
                    begin
                      reg4314 <= $signed({reg4308});
                      reg4315 <= $signed(reg4224);
                      reg4316 <= (~&(|(reg4258 < (reg4302 >= reg4219))));
                    end
                  else
                    begin
                      reg4314 <= $signed(reg4259[(3'h7):(1'h0)]);
                    end
                end
              else
                begin
                  if ((reg4286[(2'h2):(1'h1)] ?
                      $unsigned($signed($unsigned(reg4253))) : (reg4229 ?
                          forvar4293[(4'he):(2'h2)] : reg4294)))
                    begin
                      reg4310 <= (((reg4314 > (~reg4259)) + $signed($signed(reg4267))) <<< $unsigned($unsigned({reg4263})));
                    end
                  else
                    begin
                      reg4310 <= forvar4293;
                      reg4311 <= ($unsigned($unsigned(forvar4271[(3'h5):(2'h2)])) ~^ $signed(((reg4266 ?
                              reg4255 : (8'h9c)) ?
                          (^reg4283) : (!reg4315))));
                      reg4312 <= $unsigned(reg4253);
                    end
                  for (forvar4313 = (1'h0); (forvar4313 < (2'h2)); forvar4313 = (forvar4313 + (1'h1)))
                    begin
                      reg4314 <= $signed(($signed(forvar4303[(1'h1):(1'h0)]) * (reg4245 >>> reg4284[(2'h2):(1'h0)])));
                      reg4315 <= $unsigned($unsigned(forvar4280[(1'h0):(1'h0)]));
                      reg4316 <= {reg4224[(1'h0):(1'h0)]};
                      reg4317 <= reg4225[(2'h2):(2'h2)];
                    end
                  if ($unsigned((($unsigned(reg4315) || (&(8'h9f))) * reg4316[(3'h7):(3'h6)])))
                    begin
                      reg4318 <= reg4262[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg4318 <= forvar4306[(2'h3):(2'h2)];
                      reg4319 <= $signed(($unsigned($unsigned((8'ha4))) ?
                          reg4236[(4'ha):(4'ha)] : (8'hb8)));
                    end
                  for (forvar4320 = (1'h0); (forvar4320 < (1'h1)); forvar4320 = (forvar4320 + (1'h1)))
                    begin
                      reg4321 <= ({{reg4232[(3'h7):(3'h7)]}} ?
                          $signed(reg4227) : reg4239[(4'hb):(4'hb)]);
                      reg4322 <= forvar4313;
                    end
                end
              for (forvar4323 = (1'h0); (forvar4323 < (2'h3)); forvar4323 = (forvar4323 + (1'h1)))
                begin
                  if (reg4283[(3'h5):(3'h5)])
                    begin
                      reg4324 <= ((reg4241[(4'hf):(3'h4)] ?
                          reg4295[(3'h7):(1'h1)] : (~reg4279[(2'h2):(2'h2)])) ^ $unsigned((reg4307 & reg4228[(2'h3):(1'h0)])));
                      reg4325 <= (8'hb2);
                      reg4326 <= $signed($unsigned($unsigned((reg4238 ?
                          forvar4277 : reg4259))));
                      reg4327 <= (~|$unsigned(reg4298[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg4324 <= (&$unsigned((|$unsigned(reg4243))));
                      reg4325 <= {($signed(((8'hb5) ? wire4270 : (8'hb3))) ?
                              $unsigned((reg4304 ?
                                  wire4218 : reg4231)) : $unsigned($unsigned(reg4274)))};
                    end
                end
              if ((reg4304 << (!(~&reg4279[(3'h5):(1'h1)]))))
                begin
                  if ((reg4307 <<< reg4324))
                    begin
                      reg4328 <= $signed((8'ha3));
                      reg4329 <= reg4228;
                      reg4330 <= {($unsigned($signed(reg4254)) && $signed((|(8'hb0))))};
                    end
                  else
                    begin
                      reg4328 <= $signed(reg4322[(4'hd):(4'h8)]);
                      reg4329 <= reg4255[(4'h9):(3'h5)];
                      reg4330 <= $signed(($signed(((8'hba) ?
                          reg4327 : reg4278)) < reg4309[(2'h2):(2'h2)]));
                    end
                end
              else
                begin
                  if ($signed({$unsigned({forvar4293})}))
                    begin
                      reg4328 <= (|($signed({reg4254}) >>> (+(reg4283 ?
                          (8'ha3) : (8'had)))));
                      reg4329 <= (reg4225 ?
                          $unsigned(((+reg4283) <= {(8'ha5)})) : reg4219[(1'h1):(1'h0)]);
                      reg4330 <= (reg4251 <<< reg4319);
                      reg4331 <= $signed($unsigned($signed($signed(reg4249))));
                    end
                  else
                    begin
                      reg4328 <= (8'ha9);
                      reg4329 <= {($signed((~&reg4261)) ?
                              $signed(((8'h9f) ?
                                  reg4252 : reg4242)) : ((~&reg4224) ?
                                  ((8'hb6) ?
                                      reg4286 : reg4237) : forvar4301[(1'h0):(1'h0)]))};
                      reg4330 <= $unsigned($signed({reg4313}));
                    end
                  reg4332 <= $signed(reg4282[(3'h6):(3'h4)]);
                  for (forvar4333 = (1'h0); (forvar4333 < (2'h2)); forvar4333 = (forvar4333 + (1'h1)))
                    begin
                      reg4334 <= reg4257;
                      reg4335 <= $signed(($signed((reg4318 ?
                          (8'haa) : reg4250)) << reg4298));
                      reg4336 <= (~^((^{reg4326}) ?
                          reg4242[(3'h4):(2'h3)] : (+{(8'ha2)})));
                      reg4337 <= (&$signed($unsigned(reg4219[(2'h2):(1'h0)])));
                    end
                  reg4338 <= (^$unsigned(reg4275));
                end
            end
          else
            begin
              for (forvar4306 = (1'h0); (forvar4306 < (2'h3)); forvar4306 = (forvar4306 + (1'h1)))
                begin
                  for (forvar4307 = (1'h0); (forvar4307 < (2'h3)); forvar4307 = (forvar4307 + (1'h1)))
                    begin
                      reg4308 <= (((8'haa) ^~ (^(reg4232 ?
                              reg4278 : reg4297))) ?
                          $unsigned($unsigned((reg4266 > reg4312))) : $signed(forvar4323));
                      reg4309 <= forvar4333;
                      reg4310 <= ($signed($signed(reg4255[(2'h2):(2'h2)])) <<< $unsigned(($unsigned(wire4218) ?
                          (~&reg4263) : ((8'h9e) < reg4268))));
                      reg4311 <= reg4234[(2'h3):(2'h2)];
                    end
                  for (forvar4312 = (1'h0); (forvar4312 < (1'h0)); forvar4312 = (forvar4312 + (1'h1)))
                    begin
                      reg4313 <= ({(8'hb1)} ?
                          (reg4247[(4'h9):(2'h3)] ~^ {reg4286}) : forvar4307);
                      reg4314 <= (~^$signed($signed((reg4281 || reg4331))));
                      reg4315 <= reg4239[(3'h4):(2'h3)];
                    end
                  if (reg4245)
                    begin
                      reg4316 <= reg4236;
                      reg4317 <= reg4252;
                      reg4318 <= $unsigned((~$signed(reg4223[(3'h7):(3'h4)])));
                      reg4319 <= reg4318;
                    end
                  else
                    begin
                      reg4316 <= (~^{{$unsigned(reg4260)}});
                    end
                end
              reg4320 <= $signed(reg4236);
              if ({$signed(reg4292[(1'h1):(1'h0)])})
                begin
                  if (((^$signed($signed(reg4316))) ?
                      {(~^(reg4251 ?
                              (8'hba) : forvar4323))} : $signed($unsigned(reg4337))))
                    begin
                      reg4321 <= reg4251[(1'h0):(1'h0)];
                      reg4322 <= ((!$signed(forvar4312)) ^ forvar4306[(3'h7):(1'h0)]);
                      reg4323 <= {reg4259[(2'h3):(1'h0)]};
                      reg4324 <= ($unsigned(((|reg4235) ?
                          reg4276 : (forvar4312 ?
                              reg4322 : (8'ha7)))) - $signed(reg4237));
                    end
                  else
                    begin
                      reg4321 <= reg4245[(2'h2):(1'h1)];
                      reg4322 <= $signed((reg4329 ?
                          (reg4327 ?
                              (reg4254 > wire4217) : $signed(reg4307)) : (&(forvar4293 ?
                              reg4304 : reg4256))));
                      reg4323 <= reg4330;
                    end
                  if ((reg4274[(2'h3):(1'h1)] ?
                      reg4326[(4'h8):(3'h7)] : (!$unsigned(((8'hac) ?
                          reg4234 : reg4252)))))
                    begin
                      reg4325 <= reg4299[(3'h6):(2'h3)];
                      reg4326 <= (($signed((reg4291 >= (8'hb7))) ?
                          reg4284[(2'h3):(2'h3)] : ($unsigned(reg4308) == $unsigned((8'hb1)))) - ($signed($unsigned(reg4224)) ?
                          $signed($signed(reg4314)) : reg4287[(3'h6):(1'h1)]));
                      reg4327 <= ($signed($signed((+forvar4320))) | ($signed(reg4269) ?
                          {$unsigned(reg4308)} : reg4250));
                      reg4328 <= (-$unsigned(({reg4264} ?
                          (~forvar4301) : $signed(reg4254))));
                    end
                  else
                    begin
                      reg4325 <= (reg4283[(3'h7):(3'h6)] >= (reg4226 ?
                          reg4269[(4'h9):(3'h5)] : reg4295));
                      reg4326 <= (((&(~^forvar4303)) >>> (wire4218 >>> reg4289[(2'h2):(2'h2)])) & {$unsigned(reg4248[(2'h3):(2'h3)])});
                      reg4327 <= $unsigned((!reg4313[(3'h6):(2'h2)]));
                      reg4328 <= ($signed((reg4219[(2'h3):(2'h3)] ?
                          ((8'haa) <<< reg4263) : {reg4223})) && (forvar4272 ?
                          reg4250 : ((8'haf) || $signed((8'ha6)))));
                    end
                  if ((forvar4271 ? reg4282 : reg4257))
                    begin
                      reg4329 <= {reg4334};
                    end
                  else
                    begin
                      reg4329 <= (({(reg4302 ?
                              reg4279 : reg4334)} + ((forvar4320 ?
                          reg4260 : reg4304) >> (reg4282 < reg4323))) << $signed($unsigned({(8'haa)})));
                    end
                end
              else
                begin
                  for (forvar4321 = (1'h0); (forvar4321 < (2'h3)); forvar4321 = (forvar4321 + (1'h1)))
                    begin
                      reg4322 <= reg4316;
                      reg4323 <= $unsigned(reg4247);
                      reg4324 <= reg4286;
                    end
                  for (forvar4325 = (1'h0); (forvar4325 < (1'h0)); forvar4325 = (forvar4325 + (1'h1)))
                    begin
                      reg4326 <= $unsigned({{(reg4245 >= reg4286)}});
                      reg4327 <= {reg4336[(1'h0):(1'h0)]};
                      reg4328 <= wire4217[(1'h1):(1'h0)];
                      reg4329 <= wire4270[(4'ha):(3'h4)];
                    end
                end
            end
          for (forvar4339 = (1'h0); (forvar4339 < (2'h3)); forvar4339 = (forvar4339 + (1'h1)))
            begin
              if ((((^~$unsigned(reg4222)) <<< reg4308[(1'h1):(1'h1)]) ?
                  reg4320 : $signed(reg4242[(3'h4):(1'h1)])))
                begin
                  for (forvar4340 = (1'h0); (forvar4340 < (1'h1)); forvar4340 = (forvar4340 + (1'h1)))
                    begin
                      reg4341 <= reg4294[(3'h5):(1'h0)];
                      reg4342 <= ($unsigned((forvar4271[(1'h0):(1'h0)] ?
                          $signed(reg4286) : {(8'hae)})) - ($unsigned(reg4228[(2'h2):(1'h1)]) ~^ (reg4341[(1'h0):(1'h0)] ^~ reg4320[(4'h8):(2'h3)])));
                      reg4343 <= (reg4222[(1'h1):(1'h0)] - reg4325[(1'h0):(1'h0)]);
                    end
                  reg4344 <= ($unsigned(reg4327) != reg4252[(3'h4):(1'h1)]);
                end
              else
                begin
                  if ({$unsigned(reg4343)})
                    begin
                      reg4340 <= reg4266[(2'h2):(1'h0)];
                      reg4341 <= (((reg4324[(4'ha):(3'h4)] ?
                              $signed(forvar4323) : reg4279) ?
                          $unsigned($signed(reg4228)) : reg4231) <<< wire4217[(1'h0):(1'h0)]);
                      reg4342 <= ({(~^$signed((8'hae)))} - $signed((^(reg4319 ?
                          forvar4293 : reg4317))));
                    end
                  else
                    begin
                      reg4340 <= reg4319[(2'h2):(2'h2)];
                      reg4341 <= (((~|wire4216) ? reg4243 : (^(~reg4343))) ?
                          $signed((8'ha1)) : reg4289[(2'h3):(1'h1)]);
                    end
                  for (forvar4343 = (1'h0); (forvar4343 < (2'h2)); forvar4343 = (forvar4343 + (1'h1)))
                    begin
                      reg4344 <= reg4267[(3'h7):(3'h6)];
                      reg4345 <= reg4260[(1'h1):(1'h0)];
                    end
                end
              if (reg4331)
                begin
                  if ((^~$signed($signed(reg4307[(2'h2):(1'h1)]))))
                    begin
                      reg4346 <= (8'ha0);
                      reg4347 <= reg4298[(3'h7):(3'h4)];
                      reg4348 <= $signed($unsigned(reg4298));
                      reg4349 <= forvar4333[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg4346 <= (reg4294[(3'h5):(2'h3)] - (8'haa));
                      reg4347 <= ($signed((^~$unsigned((8'hb2)))) - $unsigned((|reg4256)));
                      reg4348 <= ((reg4299[(4'hf):(2'h3)] >> $signed(reg4231)) ?
                          reg4256[(2'h3):(1'h1)] : $signed($signed($unsigned(reg4297))));
                    end
                  if ((($signed($signed(forvar4271)) == $signed($unsigned((8'hb6)))) ?
                      reg4294 : reg4316[(3'h4):(2'h2)]))
                    begin
                      reg4350 <= reg4279[(1'h0):(1'h0)];
                      reg4351 <= ((~forvar4288[(4'h9):(1'h1)]) ?
                          $unsigned({reg4347}) : reg4331[(3'h6):(3'h5)]);
                    end
                  else
                    begin
                      reg4350 <= reg4338;
                      reg4351 <= ((($unsigned(reg4222) | $signed(reg4319)) >>> ({reg4299} < $unsigned((8'ha7)))) ?
                          (($signed(reg4322) ?
                              forvar4313 : (reg4334 ?
                                  forvar4303 : reg4263)) & $unsigned((+reg4297))) : {(((8'hb2) ?
                                      forvar4312 : (8'hb2)) ?
                                  (reg4263 ?
                                      forvar4313 : forvar4306) : reg4234[(2'h2):(1'h0)])});
                    end
                  reg4352 <= ($unsigned((&reg4306)) ~^ reg4315);
                end
              else
                begin
                  if (($unsigned(reg4252) | reg4304[(3'h4):(2'h2)]))
                    begin
                      reg4346 <= ($signed($unsigned(reg4254[(1'h0):(1'h0)])) | $signed(reg4268));
                    end
                  else
                    begin
                      reg4346 <= forvar4272;
                    end
                  reg4347 <= (-reg4233);
                  if ((~&(|forvar4339)))
                    begin
                      reg4348 <= ((reg4326[(4'h8):(3'h7)] ?
                              ((^(8'h9f)) ?
                                  reg4313 : reg4264[(3'h6):(3'h4)]) : (reg4234[(3'h5):(1'h1)] ?
                                  (&reg4328) : $unsigned(reg4235))) ?
                          $unsigned($unsigned((reg4228 && forvar4320))) : reg4350[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg4348 <= (((reg4311 ?
                              (reg4294 == reg4281) : (reg4313 ?
                                  (8'hb1) : (8'hab))) + $unsigned(reg4308[(3'h5):(3'h4)])) ?
                          ({$unsigned((8'hae))} <= $signed((reg4347 < reg4341))) : $unsigned((^(reg4324 - reg4249))));
                      reg4349 <= $unsigned(reg4255[(1'h1):(1'h1)]);
                    end
                end
              for (forvar4353 = (1'h0); (forvar4353 < (2'h3)); forvar4353 = (forvar4353 + (1'h1)))
                begin
                  if (((8'ha6) ~^ reg4266))
                    begin
                      reg4354 <= $signed($signed((^~reg4295)));
                      reg4355 <= reg4222;
                    end
                  else
                    begin
                      reg4354 <= (~^((8'ha2) <<< $unsigned($unsigned(reg4345))));
                      reg4355 <= reg4317[(2'h2):(1'h1)];
                    end
                end
              reg4356 <= ($unsigned((!(reg4225 ? reg4330 : reg4332))) ?
                  (-$signed(reg4337[(3'h4):(3'h4)])) : (!reg4321));
            end
          reg4357 <= ($unsigned((reg4347[(4'ha):(1'h0)] < (8'hb3))) ?
              (~^reg4315[(1'h0):(1'h0)]) : (reg4290[(3'h5):(2'h2)] ?
                  $signed(reg4285) : ((!reg4356) ?
                      (|reg4324) : (reg4225 ? reg4263 : reg4298))));
        end
      reg4358 <= reg4236;
      for (forvar4359 = (1'h0); (forvar4359 < (1'h1)); forvar4359 = (forvar4359 + (1'h1)))
        begin
          if ((reg4337[(2'h3):(2'h3)] ?
              ($signed((wire4215 ?
                  (8'ha1) : (8'ha0))) * reg4299[(4'hd):(3'h7)]) : $signed((8'hb5))))
            begin
              if (reg4342)
                begin
                  for (forvar4360 = (1'h0); (forvar4360 < (1'h0)); forvar4360 = (forvar4360 + (1'h1)))
                    begin
                      reg4361 <= $unsigned(($signed($signed(reg4259)) ?
                          (|$unsigned(reg4336)) : reg4232[(3'h5):(2'h2)]));
                    end
                  for (forvar4362 = (1'h0); (forvar4362 < (2'h2)); forvar4362 = (forvar4362 + (1'h1)))
                    begin
                      reg4363 <= (~&$signed(reg4309[(2'h3):(1'h0)]));
                    end
                  for (forvar4364 = (1'h0); (forvar4364 < (2'h3)); forvar4364 = (forvar4364 + (1'h1)))
                    begin
                      reg4365 <= ((&((reg4224 && reg4232) >> $signed(reg4283))) ?
                          reg4276 : reg4250[(1'h0):(1'h0)]);
                      reg4366 <= reg4242[(3'h4):(2'h2)];
                    end
                end
              else
                begin
                  reg4360 <= reg4296;
                end
              for (forvar4367 = (1'h0); (forvar4367 < (1'h0)); forvar4367 = (forvar4367 + (1'h1)))
                begin
                  reg4368 <= (~|reg4223);
                  if ($signed($signed((~^$signed(reg4321)))))
                    begin
                      reg4369 <= (reg4242 ?
                          ((!((8'hb2) - (8'hb1))) ?
                              ((&reg4315) < (^reg4323)) : $signed((forvar4320 != (8'hb1)))) : $signed(reg4259[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg4369 <= reg4322[(4'hc):(3'h6)];
                      reg4370 <= reg4297;
                      reg4371 <= ($unsigned($unsigned($unsigned((8'hb1)))) ^ (~&(~^reg4291)));
                      reg4372 <= ($unsigned(reg4232[(4'h9):(4'h8)]) & $signed(((reg4267 | reg4285) - (^reg4233))));
                    end
                  for (forvar4373 = (1'h0); (forvar4373 < (1'h0)); forvar4373 = (forvar4373 + (1'h1)))
                    begin
                      reg4374 <= (^$signed($unsigned((forvar4359 ?
                          reg4340 : reg4231))));
                      reg4375 <= ((~$signed($signed(reg4259))) ?
                          $signed((reg4337 ?
                              (!reg4306) : $unsigned(reg4237))) : {($unsigned((8'h9c)) > (reg4357 ?
                                  forvar4280 : (8'hb3)))});
                      reg4376 <= $unsigned($unsigned(($signed(forvar4321) <= (reg4253 ?
                          reg4307 : forvar4343))));
                    end
                end
            end
          else
            begin
              if ($unsigned(reg4371[(3'h4):(2'h3)]))
                begin
                  if ((8'hb1))
                    begin
                      reg4360 <= {reg4346};
                      reg4361 <= $signed({(~&reg4291)});
                      reg4362 <= ((~reg4257) <= forvar4373);
                    end
                  else
                    begin
                      reg4360 <= reg4248[(4'h8):(3'h5)];
                      reg4361 <= $signed($signed({{reg4287}}));
                      reg4362 <= {((((8'ha5) & reg4274) ?
                              $unsigned(reg4253) : {reg4248}) + ($signed(reg4287) ?
                              forvar4313[(2'h2):(2'h2)] : reg4287))};
                    end
                  for (forvar4363 = (1'h0); (forvar4363 < (1'h0)); forvar4363 = (forvar4363 + (1'h1)))
                    begin
                      reg4364 <= $unsigned((!$unsigned(reg4283)));
                      reg4365 <= reg4369;
                      reg4366 <= $signed((~^($signed(reg4241) ?
                          (reg4235 ^ reg4266) : $unsigned(reg4250))));
                    end
                  reg4367 <= $unsigned($signed($signed(reg4351)));
                  if (forvar4293[(4'hc):(1'h0)])
                    begin
                      reg4368 <= $unsigned((($unsigned(reg4298) ^~ $unsigned(reg4255)) + (reg4334 < (reg4334 ~^ forvar4301))));
                    end
                  else
                    begin
                      reg4368 <= (^~($signed(forvar4277[(1'h0):(1'h0)]) >= reg4226[(3'h5):(1'h0)]));
                      reg4369 <= $signed($unsigned((8'ha0)));
                    end
                end
              else
                begin
                  for (forvar4360 = (1'h0); (forvar4360 < (1'h1)); forvar4360 = (forvar4360 + (1'h1)))
                    begin
                      reg4361 <= reg4259;
                    end
                  for (forvar4362 = (1'h0); (forvar4362 < (1'h0)); forvar4362 = (forvar4362 + (1'h1)))
                    begin
                      reg4363 <= {{((reg4251 ~^ reg4349) ?
                                  $unsigned((8'h9e)) : (reg4327 ?
                                      reg4233 : reg4263))}};
                      reg4364 <= {($signed(reg4342[(4'hd):(4'hb)]) >= reg4260)};
                      reg4365 <= {(~&(8'ha1))};
                      reg4366 <= $signed(wire4216[(2'h2):(1'h0)]);
                    end
                  for (forvar4367 = (1'h0); (forvar4367 < (2'h3)); forvar4367 = (forvar4367 + (1'h1)))
                    begin
                      reg4368 <= (reg4365 != $unsigned($signed(reg4292)));
                    end
                end
              for (forvar4370 = (1'h0); (forvar4370 < (1'h0)); forvar4370 = (forvar4370 + (1'h1)))
                begin
                  for (forvar4371 = (1'h0); (forvar4371 < (2'h2)); forvar4371 = (forvar4371 + (1'h1)))
                    begin
                      reg4372 <= {((((8'hab) ?
                              reg4225 : reg4330) ^~ reg4324) >> $unsigned(((8'hac) ?
                              reg4264 : reg4367)))};
                      reg4373 <= reg4354[(2'h2):(2'h2)];
                      reg4374 <= reg4344[(2'h3):(2'h3)];
                      reg4375 <= {(~|reg4361[(1'h1):(1'h1)])};
                    end
                  for (forvar4376 = (1'h0); (forvar4376 < (1'h0)); forvar4376 = (forvar4376 + (1'h1)))
                    begin
                      reg4377 <= $signed((8'hba));
                      reg4378 <= reg4323[(2'h2):(2'h2)];
                    end
                  reg4379 <= (~^$unsigned(reg4219[(4'hb):(2'h2)]));
                  reg4380 <= $signed(reg4324[(1'h1):(1'h1)]);
                end
              for (forvar4381 = (1'h0); (forvar4381 < (1'h0)); forvar4381 = (forvar4381 + (1'h1)))
                begin
                  for (forvar4382 = (1'h0); (forvar4382 < (1'h0)); forvar4382 = (forvar4382 + (1'h1)))
                    begin
                      reg4383 <= $signed((-(reg4299[(4'hc):(4'hb)] ?
                          reg4253 : (reg4380 ? forvar4301 : reg4250))));
                      reg4384 <= ({($signed(reg4334) ?
                                  $unsigned(reg4274) : (reg4350 ?
                                      (8'hb4) : reg4344))} ?
                          {reg4276[(4'h9):(3'h6)]} : $signed($signed(((8'hb3) ?
                              (8'ha5) : (8'hb6)))));
                      reg4385 <= $unsigned(reg4322[(3'h6):(1'h0)]);
                      reg4386 <= $signed($signed($unsigned((~|reg4319))));
                    end
                  if ((8'h9e))
                    begin
                      reg4387 <= (+forvar4301[(1'h0):(1'h0)]);
                      reg4388 <= $unsigned($signed(($unsigned(reg4238) ?
                          (8'had) : (~|reg4298))));
                    end
                  else
                    begin
                      reg4387 <= $unsigned(reg4252[(4'hc):(2'h3)]);
                    end
                  if ((^$unsigned(($unsigned(reg4365) + (forvar4293 ?
                      reg4358 : reg4349)))))
                    begin
                      reg4389 <= reg4274;
                      reg4390 <= reg4361[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg4389 <= (8'hac);
                      reg4390 <= forvar4360;
                      reg4391 <= forvar4321[(2'h3):(2'h3)];
                    end
                end
              if ((forvar4306 << $unsigned((reg4278[(4'h9):(1'h0)] <= ((8'ha8) ?
                  forvar4373 : reg4285)))))
                begin
                  if (reg4222)
                    begin
                      reg4392 <= (reg4233 ?
                          $unsigned(((+reg4307) ?
                              forvar4360[(2'h3):(1'h1)] : $unsigned(reg4372))) : (~&$unsigned((reg4334 != reg4232))));
                      reg4393 <= $signed($unsigned({$unsigned(forvar4382)}));
                      reg4394 <= $unsigned(reg4224[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg4392 <= $signed(reg4289[(3'h4):(1'h0)]);
                      reg4393 <= $signed((^($unsigned(reg4266) ^~ (forvar4382 << reg4315))));
                      reg4394 <= ((($unsigned(reg4347) <<< $signed(reg4266)) ?
                          ($unsigned(reg4380) ?
                              (+reg4239) : $unsigned((8'hb0))) : (forvar4359 + {forvar4306})) >= (|reg4321[(2'h2):(1'h1)]));
                    end
                  if ((reg4324[(2'h3):(2'h3)] * (!$signed((|reg4275)))))
                    begin
                      reg4395 <= {$unsigned((~|(forvar4320 >> reg4231)))};
                    end
                  else
                    begin
                      reg4395 <= (!reg4313[(4'h8):(3'h7)]);
                      reg4396 <= $signed((~$unsigned(reg4298[(4'h8):(3'h6)])));
                      reg4397 <= $signed(((8'haf) > ((reg4243 ?
                              reg4386 : reg4281) ?
                          (reg4310 <= reg4223) : ((8'ha1) ?
                              forvar4343 : reg4266))));
                    end
                end
              else
                begin
                  reg4392 <= reg4363[(1'h1):(1'h0)];
                  for (forvar4393 = (1'h0); (forvar4393 < (1'h1)); forvar4393 = (forvar4393 + (1'h1)))
                    begin
                      reg4394 <= reg4369;
                      reg4395 <= $signed((($signed(wire4270) ?
                              (+reg4372) : $signed(reg4311)) ?
                          reg4395[(3'h5):(3'h5)] : {(^~reg4358)}));
                    end
                  for (forvar4396 = (1'h0); (forvar4396 < (1'h0)); forvar4396 = (forvar4396 + (1'h1)))
                    begin
                      reg4397 <= $signed((reg4222 ?
                          (reg4380 ?
                              reg4237 : (reg4275 ?
                                  reg4306 : forvar4340)) : (|(reg4317 ?
                              reg4370 : (8'hb3)))));
                      reg4398 <= reg4356[(3'h7):(1'h0)];
                      reg4399 <= ($unsigned(($signed(reg4326) ?
                              (reg4338 >>> reg4307) : (reg4224 ?
                                  reg4310 : forvar4382))) ?
                          $unsigned(($unsigned(reg4313) >>> reg4396)) : (~|reg4336));
                      reg4400 <= $signed(forvar4271[(2'h3):(2'h3)]);
                    end
                end
            end
        end
      if ((($signed((reg4324 >> reg4316)) ? forvar4343 : reg4254) ?
          (-reg4350) : reg4343))
        begin
          reg4401 <= $signed({$unsigned(((8'h9d) ? reg4364 : reg4385))});
        end
      else
        begin
          for (forvar4401 = (1'h0); (forvar4401 < (2'h2)); forvar4401 = (forvar4401 + (1'h1)))
            begin
              for (forvar4402 = (1'h0); (forvar4402 < (2'h2)); forvar4402 = (forvar4402 + (1'h1)))
                begin
                  reg4403 <= $unsigned((reg4349 && $signed({reg4313})));
                  if (reg4387[(3'h5):(3'h4)])
                    begin
                      reg4404 <= $signed((reg4310 ?
                          (reg4363[(1'h1):(1'h1)] ?
                              (reg4249 ?
                                  reg4373 : reg4219) : $unsigned(reg4389)) : $signed((reg4312 ?
                              reg4321 : forvar4307))));
                      reg4405 <= reg4375;
                    end
                  else
                    begin
                      reg4404 <= (reg4393[(2'h2):(1'h1)] ^~ (~($unsigned(reg4342) >> reg4257)));
                      reg4405 <= $unsigned($unsigned($signed((~&reg4264))));
                      reg4406 <= $signed(reg4338[(2'h3):(1'h0)]);
                    end
                end
            end
          for (forvar4407 = (1'h0); (forvar4407 < (1'h0)); forvar4407 = (forvar4407 + (1'h1)))
            begin
              reg4408 <= (~(reg4300 ?
                  ((!reg4348) ? reg4269 : reg4344[(1'h1):(1'h1)]) : ((reg4384 ?
                      reg4251 : reg4324) == reg4335)));
            end
          for (forvar4409 = (1'h0); (forvar4409 < (1'h0)); forvar4409 = (forvar4409 + (1'h1)))
            begin
              if ($unsigned((-(-(reg4311 ^~ forvar4272)))))
                begin
                  reg4410 <= (reg4378 == ((8'ha1) * ((^reg4389) >= (^~reg4314))));
                end
              else
                begin
                  if ((8'hb3))
                    begin
                      reg4410 <= {($signed((|reg4345)) ?
                              ((-(8'h9c)) << reg4392) : $unsigned($unsigned(forvar4323)))};
                    end
                  else
                    begin
                      reg4410 <= $signed(forvar4382[(3'h6):(1'h1)]);
                      reg4411 <= $signed(({(~&forvar4364)} << (&$unsigned(reg4260))));
                    end
                end
              if (reg4406[(2'h3):(1'h0)])
                begin
                  reg4412 <= (reg4395 ?
                      $unsigned($signed((~&forvar4306))) : {reg4304});
                  if ((((&(&reg4297)) ?
                      ({reg4313} ?
                          (reg4401 ?
                              reg4241 : (8'hac)) : (^~wire4217)) : reg4317) || $signed($signed(reg4337[(2'h2):(2'h2)]))))
                    begin
                      reg4413 <= $signed((-forvar4393[(2'h3):(1'h0)]));
                      reg4414 <= ((~^$unsigned($signed(reg4393))) + forvar4343);
                      reg4415 <= (8'h9c);
                    end
                  else
                    begin
                      reg4413 <= reg4309;
                    end
                end
              else
                begin
                  reg4412 <= forvar4402[(4'h8):(1'h0)];
                  reg4413 <= $signed(forvar4325);
                end
              if ({(-$signed((&reg4318)))})
                begin
                  reg4416 <= $signed({(8'haa)});
                end
              else
                begin
                  if (($unsigned($unsigned((8'ha8))) ?
                      {((~&reg4268) > $unsigned(reg4396))} : (forvar4364[(1'h1):(1'h1)] <<< reg4400[(3'h6):(3'h4)])))
                    begin
                      reg4416 <= (({$unsigned(reg4226)} && reg4326[(3'h4):(1'h1)]) ^~ reg4389[(1'h0):(1'h0)]);
                      reg4417 <= (|(($unsigned(forvar4362) ?
                              (reg4296 >= (8'ha2)) : (|reg4246)) ?
                          ($unsigned(reg4283) >> $signed(reg4374)) : $signed(reg4274)));
                    end
                  else
                    begin
                      reg4416 <= ($unsigned(reg4392) ^ (~|((~reg4252) ~^ {forvar4364})));
                      reg4417 <= (~&reg4390);
                      reg4418 <= {$unsigned((reg4251 ?
                              forvar4401 : $signed(reg4352)))};
                    end
                  reg4419 <= (&(reg4336 ?
                      ((reg4314 - (8'hb8)) * $signed(forvar4353)) : (~^(8'hb6))));
                  reg4420 <= (((8'hb4) & (~&(reg4335 < reg4274))) && ((|reg4269[(4'hb):(2'h3)]) > (|(reg4329 - (8'hae)))));
                  reg4421 <= $unsigned($unsigned((reg4259 ^~ ((8'ha9) & (8'ha3)))));
                end
              if ($unsigned((((^forvar4320) >> $unsigned(reg4346)) ^ $signed((reg4256 || reg4419)))))
                begin
                  reg4422 <= reg4219;
                  for (forvar4423 = (1'h0); (forvar4423 < (2'h3)); forvar4423 = (forvar4423 + (1'h1)))
                    begin
                      reg4424 <= $signed(reg4420);
                      reg4425 <= ((~|(~{forvar4359})) ^~ reg4238[(2'h2):(2'h2)]);
                      reg4426 <= (($signed(((8'ha1) ? reg4403 : reg4262)) ?
                          ($signed(forvar4271) + forvar4312) : ($unsigned(reg4404) * (reg4281 <<< (8'ha0)))) - reg4305);
                    end
                end
              else
                begin
                  for (forvar4422 = (1'h0); (forvar4422 < (2'h3)); forvar4422 = (forvar4422 + (1'h1)))
                    begin
                      reg4423 <= ((^~$unsigned(reg4275)) ?
                          (((forvar4359 ? (8'hb2) : (8'had)) ?
                              $unsigned((8'ha3)) : (&(8'h9c))) | $signed(reg4308)) : $signed((((8'hb2) ^~ forvar4340) ?
                              reg4312 : (reg4400 ? reg4253 : wire4218))));
                    end
                  if (((^$unsigned(wire4216)) ?
                      reg4368 : (reg4306[(1'h0):(1'h0)] ?
                          $signed((reg4263 << reg4282)) : (!(~&(8'hb4))))))
                    begin
                      reg4424 <= (~$signed(reg4305));
                      reg4425 <= $signed(reg4302);
                    end
                  else
                    begin
                      reg4424 <= (~^(8'h9c));
                      reg4425 <= ((8'ha3) ?
                          (&$unsigned(reg4413[(4'hb):(3'h6)])) : wire4216[(1'h1):(1'h1)]);
                    end
                  if ((reg4294 ?
                      reg4370[(1'h0):(1'h0)] : ($unsigned(reg4367) & (-(forvar4293 ?
                          reg4413 : (8'ha8))))))
                    begin
                      reg4426 <= {((((8'hb0) - reg4354) ?
                                  reg4267 : (reg4377 ? reg4332 : forvar4312)) ?
                              $signed(reg4352[(4'hb):(4'hb)]) : $unsigned((|reg4264)))};
                      reg4427 <= $unsigned((~(~&(reg4350 ^ reg4372))));
                    end
                  else
                    begin
                      reg4426 <= (~|(~$signed((forvar4360 ?
                          (8'hae) : reg4289))));
                      reg4427 <= $signed($signed(((!reg4389) * (reg4369 * (8'h9e)))));
                      reg4428 <= $signed(reg4354);
                      reg4429 <= {{({reg4414} < reg4313[(1'h1):(1'h1)])}};
                    end
                end
            end
        end
    end
  assign wire4430 = reg4290;
  always
    @(posedge clk) begin
      if ({(($signed((8'hac)) >= (reg4384 | reg4420)) ?
              reg4269[(2'h3):(1'h0)] : reg4263[(1'h0):(1'h0)])})
        begin
          for (forvar4431 = (1'h0); (forvar4431 < (1'h0)); forvar4431 = (forvar4431 + (1'h1)))
            begin
              for (forvar4432 = (1'h0); (forvar4432 < (1'h0)); forvar4432 = (forvar4432 + (1'h1)))
                begin
                  for (forvar4433 = (1'h0); (forvar4433 < (2'h3)); forvar4433 = (forvar4433 + (1'h1)))
                    begin
                      reg4434 <= $signed(reg4318);
                    end
                  for (forvar4435 = (1'h0); (forvar4435 < (1'h1)); forvar4435 = (forvar4435 + (1'h1)))
                    begin
                      reg4436 <= $signed((((reg4241 >>> (8'hb6)) ?
                              $signed(reg4319) : $signed(reg4225)) ?
                          reg4389[(1'h1):(1'h1)] : (!(reg4298 + reg4284))));
                      reg4437 <= $signed(reg4352[(4'hc):(4'h8)]);
                      reg4438 <= reg4240;
                    end
                  if ({(!((reg4314 ? reg4321 : (8'had)) ?
                          (reg4232 != (8'ha0)) : (!reg4232)))})
                    begin
                      reg4439 <= {$unsigned(($signed((8'ha1)) ?
                              $signed((8'hb2)) : reg4268))};
                      reg4440 <= (((!forvar4435[(2'h3):(1'h0)]) >> reg4347) >= ($unsigned(reg4403[(2'h2):(2'h2)]) ?
                          ((reg4358 ~^ reg4242) ?
                              (8'had) : $signed(reg4306)) : $unsigned(((8'h9c) ?
                              reg4317 : reg4237))));
                      reg4441 <= ((8'hb8) ?
                          (|reg4360[(1'h1):(1'h0)]) : reg4390[(3'h6):(3'h6)]);
                    end
                  else
                    begin
                      reg4439 <= (&reg4332);
                      reg4440 <= (8'hb6);
                    end
                  reg4442 <= (^$unsigned(({(8'haa)} <<< reg4398)));
                end
            end
        end
      else
        begin
          for (forvar4431 = (1'h0); (forvar4431 < (1'h1)); forvar4431 = (forvar4431 + (1'h1)))
            begin
              for (forvar4432 = (1'h0); (forvar4432 < (1'h0)); forvar4432 = (forvar4432 + (1'h1)))
                begin
                  reg4433 <= ($signed((+reg4250)) - $signed((-(8'h9c))));
                end
            end
          reg4434 <= $signed(reg4427);
          if (reg4400)
            begin
              if (((^(~|$signed(reg4406))) ?
                  (~&reg4300[(1'h1):(1'h0)]) : ($unsigned((reg4341 ?
                          (8'haf) : (8'ha8))) ?
                      $unsigned(reg4246) : reg4361)))
                begin
                  for (forvar4435 = (1'h0); (forvar4435 < (1'h0)); forvar4435 = (forvar4435 + (1'h1)))
                    begin
                      reg4436 <= $signed($unsigned((reg4222 >> (reg4373 ?
                          reg4440 : reg4335))));
                    end
                  if ($signed(reg4294[(1'h0):(1'h0)]))
                    begin
                      reg4437 <= $signed(reg4234);
                      reg4438 <= reg4370[(3'h4):(2'h2)];
                      reg4439 <= (~^reg4254);
                      reg4440 <= reg4355[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg4437 <= $unsigned(reg4248[(3'h4):(2'h3)]);
                      reg4438 <= $signed((8'haa));
                      reg4439 <= ((+(~(~reg4268))) > ($unsigned((reg4401 ?
                          reg4328 : reg4330)) > ($signed(reg4314) ?
                          (reg4264 ? reg4344 : reg4355) : $unsigned(reg4243))));
                    end
                  for (forvar4441 = (1'h0); (forvar4441 < (1'h1)); forvar4441 = (forvar4441 + (1'h1)))
                    begin
                      reg4442 <= reg4403[(2'h3):(2'h3)];
                      reg4443 <= ($signed(($signed(reg4256) ?
                              (^~reg4302) : reg4442[(3'h5):(2'h3)])) ?
                          $unsigned($unsigned(reg4376)) : $signed($unsigned((reg4380 ?
                              (8'ha0) : reg4440))));
                      reg4444 <= (reg4369 && ($unsigned((|reg4219)) * $signed($signed(reg4375))));
                    end
                end
              else
                begin
                  reg4435 <= $unsigned($unsigned((^(&reg4441))));
                  if (forvar4433)
                    begin
                      reg4436 <= reg4264;
                      reg4437 <= (&(|reg4349));
                    end
                  else
                    begin
                      reg4436 <= ($unsigned($signed({reg4345})) ?
                          $unsigned((-$unsigned((8'ha9)))) : (!((wire4217 & reg4285) - reg4234)));
                    end
                end
              if ($signed((reg4292 ?
                  ($signed(reg4227) ? $signed(reg4383) : {reg4329}) : reg4423)))
                begin
                  for (forvar4445 = (1'h0); (forvar4445 < (2'h2)); forvar4445 = (forvar4445 + (1'h1)))
                    begin
                      reg4446 <= (~(($unsigned(reg4246) < reg4379) > $unsigned((reg4240 <= reg4269))));
                      reg4447 <= ({wire4217[(1'h0):(1'h0)]} ?
                          $signed((^~(reg4357 << reg4404))) : reg4385);
                      reg4448 <= reg4362;
                    end
                  if ($unsigned({(&reg4427[(2'h2):(2'h2)])}))
                    begin
                      reg4449 <= reg4329[(2'h2):(1'h0)];
                      reg4450 <= $unsigned(reg4347);
                      reg4451 <= reg4300;
                    end
                  else
                    begin
                      reg4449 <= {($signed($unsigned(reg4447)) == ($signed(reg4390) - reg4310))};
                    end
                  for (forvar4452 = (1'h0); (forvar4452 < (1'h0)); forvar4452 = (forvar4452 + (1'h1)))
                    begin
                      reg4453 <= (^$unsigned((reg4249[(2'h2):(1'h0)] ?
                          (|reg4433) : reg4429[(1'h1):(1'h0)])));
                      reg4454 <= reg4429;
                      reg4455 <= ($signed(reg4366[(4'h9):(3'h5)]) <<< wire4430);
                    end
                end
              else
                begin
                  for (forvar4445 = (1'h0); (forvar4445 < (2'h2)); forvar4445 = (forvar4445 + (1'h1)))
                    begin
                      reg4446 <= reg4329[(2'h2):(1'h0)];
                      reg4447 <= (($signed(((8'ha5) - reg4390)) << (^~(-reg4231))) ?
                          (8'ha7) : (((reg4411 ~^ reg4365) <<< (8'hb2)) ?
                              {(reg4362 >= reg4286)} : reg4314));
                      reg4448 <= reg4239;
                    end
                  for (forvar4449 = (1'h0); (forvar4449 < (1'h0)); forvar4449 = (forvar4449 + (1'h1)))
                    begin
                      reg4450 <= reg4225[(2'h2):(1'h0)];
                      reg4451 <= $signed(reg4444);
                    end
                end
            end
          else
            begin
              reg4435 <= $unsigned(reg4310[(4'hd):(1'h1)]);
              for (forvar4436 = (1'h0); (forvar4436 < (1'h1)); forvar4436 = (forvar4436 + (1'h1)))
                begin
                  for (forvar4437 = (1'h0); (forvar4437 < (1'h1)); forvar4437 = (forvar4437 + (1'h1)))
                    begin
                      reg4438 <= $unsigned((reg4363[(4'h8):(3'h5)] >> $signed((+reg4340))));
                    end
                end
              for (forvar4439 = (1'h0); (forvar4439 < (2'h3)); forvar4439 = (forvar4439 + (1'h1)))
                begin
                  for (forvar4440 = (1'h0); (forvar4440 < (1'h0)); forvar4440 = (forvar4440 + (1'h1)))
                    begin
                      reg4441 <= ($signed((((8'hae) ? (8'ha9) : reg4397) ?
                          {reg4287} : {reg4322})) != forvar4452[(1'h0):(1'h0)]);
                    end
                  for (forvar4442 = (1'h0); (forvar4442 < (2'h3)); forvar4442 = (forvar4442 + (1'h1)))
                    begin
                      reg4443 <= reg4406;
                      reg4444 <= (+$signed(reg4390[(4'h9):(3'h6)]));
                      reg4445 <= reg4255[(4'h8):(2'h3)];
                    end
                end
            end
        end
      for (forvar4456 = (1'h0); (forvar4456 < (2'h3)); forvar4456 = (forvar4456 + (1'h1)))
        begin
          for (forvar4457 = (1'h0); (forvar4457 < (1'h1)); forvar4457 = (forvar4457 + (1'h1)))
            begin
              for (forvar4458 = (1'h0); (forvar4458 < (1'h1)); forvar4458 = (forvar4458 + (1'h1)))
                begin
                  for (forvar4459 = (1'h0); (forvar4459 < (1'h1)); forvar4459 = (forvar4459 + (1'h1)))
                    begin
                      reg4460 <= reg4433;
                      reg4461 <= (((reg4323 != (reg4311 ?
                              wire4217 : reg4258)) | {(reg4376 ?
                                  (8'hb0) : wire4270)}) ?
                          (-$signed((reg4245 ?
                              reg4362 : reg4327))) : reg4246[(4'hd):(3'h6)]);
                    end
                end
              if ((reg4454[(4'h9):(3'h5)] || (($signed(reg4385) >> (reg4368 ^ reg4337)) ?
                  (8'ha7) : ((reg4281 ?
                      reg4411 : (8'hb6)) >>> $unsigned(reg4416)))))
                begin
                  for (forvar4462 = (1'h0); (forvar4462 < (2'h3)); forvar4462 = (forvar4462 + (1'h1)))
                    begin
                      reg4463 <= $unsigned((~|((reg4305 ? reg4328 : reg4400) ?
                          reg4281[(4'hd):(1'h1)] : {reg4314})));
                    end
                  if ((reg4222 > $unsigned((~&((8'h9e) ? (8'haf) : reg4461)))))
                    begin
                      reg4464 <= (8'hac);
                    end
                  else
                    begin
                      reg4464 <= $unsigned(({reg4348} ?
                          reg4448 : $unsigned((reg4363 ^ reg4325))));
                      reg4465 <= reg4347[(4'h9):(3'h7)];
                    end
                  for (forvar4466 = (1'h0); (forvar4466 < (2'h2)); forvar4466 = (forvar4466 + (1'h1)))
                    begin
                      reg4467 <= {((((8'hac) << reg4238) ?
                              (8'hb7) : $unsigned(reg4315)) || (8'hb7))};
                      reg4468 <= $signed($signed({(8'ha3)}));
                    end
                  if ((+reg4397[(1'h1):(1'h0)]))
                    begin
                      reg4469 <= ((+($unsigned(reg4226) + (~|reg4370))) ?
                          (forvar4456[(4'ha):(2'h2)] < {reg4415}) : reg4398[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg4469 <= reg4235[(2'h3):(2'h3)];
                      reg4470 <= (reg4239[(4'h9):(3'h5)] * (reg4239 ?
                          reg4454[(4'h8):(4'h8)] : ($unsigned(forvar4449) ?
                              $unsigned(reg4341) : {reg4308})));
                      reg4471 <= ((((reg4330 ?
                              (8'ha5) : reg4378) | $signed(reg4428)) ?
                          (reg4276[(5'h10):(4'hc)] <= (-reg4410)) : {reg4380[(2'h3):(2'h3)]}) >= ((~{reg4435}) ?
                          $unsigned((reg4440 ?
                              reg4254 : reg4380)) : $signed($signed(reg4377))));
                    end
                end
              else
                begin
                  reg4462 <= {(reg4354 ?
                          reg4439[(3'h5):(3'h5)] : ((reg4311 ?
                              reg4403 : reg4464) & reg4310[(3'h4):(1'h1)]))};
                end
            end
          for (forvar4472 = (1'h0); (forvar4472 < (1'h0)); forvar4472 = (forvar4472 + (1'h1)))
            begin
              if ({reg4424})
                begin
                  if (reg4361)
                    begin
                      reg4473 <= $unsigned(reg4249);
                      reg4474 <= reg4380;
                      reg4475 <= $unsigned(($unsigned((^~reg4313)) ?
                          $unsigned((+(8'hb5))) : reg4282[(2'h3):(2'h2)]));
                      reg4476 <= $signed($signed((~reg4447[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg4473 <= (reg4404 ?
                          (!({reg4241} ? reg4224 : reg4246)) : ((8'h9e) ?
                              {((8'hb9) ?
                                      reg4285 : (8'hb1))} : ($signed((8'hb5)) >> $unsigned(reg4435))));
                      reg4474 <= reg4400[(3'h6):(1'h1)];
                      reg4475 <= reg4420;
                      reg4476 <= wire4218;
                    end
                  if ($signed((reg4260 ?
                      (^~$signed(reg4377)) : $signed((reg4444 || (8'hb3))))))
                    begin
                      reg4477 <= {$signed(reg4373)};
                    end
                  else
                    begin
                      reg4477 <= ($unsigned((^(reg4388 << reg4348))) > reg4312);
                      reg4478 <= ($signed(reg4389[(1'h0):(1'h0)]) ?
                          (reg4226 ?
                              (-reg4419[(1'h0):(1'h0)]) : $unsigned(reg4318)) : {$signed($signed(reg4474))});
                    end
                end
              else
                begin
                  for (forvar4473 = (1'h0); (forvar4473 < (2'h3)); forvar4473 = (forvar4473 + (1'h1)))
                    begin
                      reg4474 <= (-$signed((~|(|reg4219))));
                    end
                  if ({(8'hb9)})
                    begin
                      reg4475 <= (($unsigned((8'hac)) << (~(~|reg4247))) ^ ((~|$signed(reg4429)) ?
                          ((^forvar4462) ?
                              (forvar4473 && reg4281) : (reg4447 > reg4234)) : reg4367));
                    end
                  else
                    begin
                      reg4475 <= (((~&reg4362[(1'h0):(1'h0)]) << ($signed((8'hb9)) ?
                              $signed(reg4308) : (reg4415 ^~ reg4260))) ?
                          ($unsigned(((8'ha5) ? (8'ha6) : reg4453)) ?
                              reg4371 : (&$unsigned(reg4285))) : reg4401[(1'h0):(1'h0)]);
                    end
                  for (forvar4476 = (1'h0); (forvar4476 < (1'h0)); forvar4476 = (forvar4476 + (1'h1)))
                    begin
                      reg4477 <= ((reg4439[(4'h9):(4'h9)] ?
                          $unsigned(wire4270[(3'h7):(1'h0)]) : reg4423) ~^ $signed($unsigned((reg4302 ?
                          reg4307 : reg4222))));
                      reg4478 <= $unsigned((8'haf));
                    end
                  reg4479 <= $signed((reg4453[(2'h3):(1'h0)] ?
                      reg4401[(2'h3):(2'h2)] : reg4314[(2'h2):(1'h1)]));
                end
            end
          for (forvar4480 = (1'h0); (forvar4480 < (2'h2)); forvar4480 = (forvar4480 + (1'h1)))
            begin
              for (forvar4481 = (1'h0); (forvar4481 < (2'h2)); forvar4481 = (forvar4481 + (1'h1)))
                begin
                  for (forvar4482 = (1'h0); (forvar4482 < (1'h1)); forvar4482 = (forvar4482 + (1'h1)))
                    begin
                      reg4483 <= $signed($unsigned(reg4376));
                      reg4484 <= ($unsigned((((8'hb4) != reg4323) ?
                          (reg4340 == reg4358) : {(8'ha9)})) << reg4256);
                      reg4485 <= ($signed($signed(reg4363)) ?
                          $signed($unsigned((reg4247 < (8'hba)))) : reg4413);
                    end
                end
            end
        end
      if (reg4427)
        begin
          for (forvar4486 = (1'h0); (forvar4486 < (2'h2)); forvar4486 = (forvar4486 + (1'h1)))
            begin
              reg4487 <= reg4415[(3'h7):(1'h1)];
            end
          reg4488 <= ($signed($signed((reg4485 ? reg4416 : reg4295))) ?
              reg4375 : ((reg4388 ?
                  $unsigned(reg4304) : $signed(reg4310)) ^~ (!reg4465)));
          reg4489 <= (&(^~$unsigned($unsigned(reg4390))));
        end
      else
        begin
          for (forvar4486 = (1'h0); (forvar4486 < (2'h3)); forvar4486 = (forvar4486 + (1'h1)))
            begin
              if (((!(reg4474[(2'h2):(1'h0)] - ((8'haf) && reg4225))) ?
                  ($unsigned({(8'ha7)}) <= $unsigned({forvar4431})) : (reg4233[(3'h6):(3'h6)] == {(forvar4457 || reg4477)})))
                begin
                  reg4487 <= reg4489;
                  for (forvar4488 = (1'h0); (forvar4488 < (2'h2)); forvar4488 = (forvar4488 + (1'h1)))
                    begin
                      reg4489 <= $signed((~(~|(~|reg4294))));
                      reg4490 <= {((~(~&reg4317)) > {(-reg4399)})};
                      reg4491 <= $signed((8'hae));
                      reg4492 <= $signed($signed(({reg4296} ?
                          ((8'ha4) | reg4298) : (reg4283 ?
                              reg4260 : (8'haa)))));
                    end
                  reg4493 <= $unsigned(($unsigned(forvar4476) ?
                      reg4348 : $unsigned($signed((8'hb8)))));
                end
              else
                begin
                  for (forvar4487 = (1'h0); (forvar4487 < (2'h2)); forvar4487 = (forvar4487 + (1'h1)))
                    begin
                      reg4488 <= $unsigned($signed(({(8'ha5)} ?
                          $unsigned(reg4358) : $unsigned((8'hb2)))));
                    end
                  if (((~&reg4239[(2'h2):(1'h0)]) != reg4455[(1'h0):(1'h0)]))
                    begin
                      reg4489 <= $unsigned(($unsigned(reg4298[(3'h6):(3'h5)]) <<< $unsigned((^reg4233))));
                      reg4490 <= $signed((&$unsigned((~reg4299))));
                      reg4491 <= (8'h9f);
                    end
                  else
                    begin
                      reg4489 <= $unsigned((reg4256[(1'h0):(1'h0)] > ((~reg4266) ?
                          reg4380 : reg4461[(2'h3):(1'h1)])));
                      reg4490 <= $unsigned((reg4327[(4'hd):(2'h2)] ?
                          reg4267 : ((reg4319 & reg4417) > $signed(reg4283))));
                      reg4491 <= (^~(-reg4355));
                    end
                  if (reg4393)
                    begin
                      reg4492 <= (^reg4356[(4'h9):(2'h3)]);
                      reg4493 <= (8'hac);
                      reg4494 <= reg4331[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg4492 <= $signed($unsigned($unsigned($unsigned(reg4255))));
                      reg4493 <= $unsigned({$signed(reg4462[(2'h2):(1'h0)])});
                    end
                end
            end
          if (reg4337[(2'h2):(1'h0)])
            begin
              for (forvar4495 = (1'h0); (forvar4495 < (2'h2)); forvar4495 = (forvar4495 + (1'h1)))
                begin
                  if (($signed((((8'haa) ? reg4485 : wire4215) ?
                      (reg4423 + forvar4472) : reg4401)) | $unsigned((~&(~|reg4306)))))
                    begin
                      reg4496 <= $unsigned((($signed(reg4358) ?
                              (!reg4449) : (-reg4435)) ?
                          (8'hb4) : reg4238));
                      reg4497 <= (-((-{reg4400}) ?
                          reg4405 : (&$unsigned(reg4379))));
                      reg4498 <= reg4469;
                      reg4499 <= $unsigned((~|($signed(reg4370) >> (8'hab))));
                    end
                  else
                    begin
                      reg4496 <= $signed(reg4282[(3'h5):(2'h2)]);
                      reg4497 <= reg4366[(3'h6):(3'h5)];
                      reg4498 <= reg4492[(1'h0):(1'h0)];
                      reg4499 <= $unsigned(($signed($signed(reg4370)) ?
                          reg4237 : reg4378[(1'h1):(1'h1)]));
                    end
                end
              for (forvar4500 = (1'h0); (forvar4500 < (2'h3)); forvar4500 = (forvar4500 + (1'h1)))
                begin
                  for (forvar4501 = (1'h0); (forvar4501 < (2'h2)); forvar4501 = (forvar4501 + (1'h1)))
                    begin
                      reg4502 <= ((reg4488 + (8'hab)) ?
                          $signed($signed($unsigned((8'ha3)))) : reg4233[(3'h7):(3'h7)]);
                      reg4503 <= (~$signed({(forvar4466 && wire4215)}));
                    end
                  for (forvar4504 = (1'h0); (forvar4504 < (1'h0)); forvar4504 = (forvar4504 + (1'h1)))
                    begin
                      reg4505 <= ((~(-{reg4426})) ?
                          ((8'ha0) ?
                              ((reg4297 != reg4479) ?
                                  (&(8'ha0)) : $signed(reg4453)) : {(reg4309 ?
                                      reg4417 : reg4497)}) : ((~^$unsigned(reg4326)) | $signed(reg4369)));
                    end
                  reg4506 <= (8'ha2);
                  for (forvar4507 = (1'h0); (forvar4507 < (1'h0)); forvar4507 = (forvar4507 + (1'h1)))
                    begin
                      reg4508 <= (((&reg4468) ?
                              reg4423 : (reg4440 ?
                                  $signed(reg4474) : (forvar4441 >>> (8'hb6)))) ?
                          (!reg4314) : (8'ha0));
                      reg4509 <= reg4340;
                      reg4510 <= $signed(reg4329[(2'h2):(1'h0)]);
                    end
                end
            end
          else
            begin
              for (forvar4495 = (1'h0); (forvar4495 < (1'h0)); forvar4495 = (forvar4495 + (1'h1)))
                begin
                  if (({(+(reg4469 ? reg4287 : reg4388))} ?
                      {{forvar4487[(3'h5):(3'h4)]}} : reg4295[(4'h8):(3'h4)]))
                    begin
                      reg4496 <= reg4370;
                      reg4497 <= $unsigned(reg4429);
                      reg4498 <= (-($unsigned((reg4219 * (8'h9e))) ?
                          (^~{reg4314}) : (-((8'hae) ^~ (8'hb8)))));
                      reg4499 <= reg4411;
                    end
                  else
                    begin
                      reg4496 <= $signed({$signed(reg4324)});
                    end
                  if (((&$unsigned($unsigned(reg4479))) == $unsigned((((8'hac) ?
                      (8'ha1) : reg4418) | (8'ha7)))))
                    begin
                      reg4500 <= $unsigned({((&reg4508) ?
                              $unsigned((8'ha6)) : $unsigned(reg4366))});
                      reg4501 <= reg4290;
                      reg4502 <= $unsigned(reg4372[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg4500 <= reg4440;
                      reg4501 <= (reg4373[(4'h9):(4'h9)] ?
                          $signed({reg4435}) : (~(reg4421 ?
                              (reg4502 ?
                                  reg4509 : reg4476) : ((8'ha2) <= reg4420))));
                    end
                  if (($unsigned($signed(wire4270)) ?
                      ((forvar4507[(2'h2):(1'h0)] ?
                              (reg4229 & reg4377) : (^~reg4335)) ?
                          $signed(((8'ha5) ?
                              (8'hb6) : reg4227)) : (~|$unsigned(reg4484))) : ((reg4332 ^ $signed(reg4444)) <<< (!$unsigned(reg4391)))))
                    begin
                      reg4503 <= $unsigned((8'h9c));
                      reg4504 <= {(^((reg4335 ?
                              reg4493 : reg4307) && reg4291[(2'h3):(2'h3)]))};
                    end
                  else
                    begin
                      reg4503 <= ($signed($unsigned((^reg4414))) < ({$unsigned(reg4450)} >> $signed((-reg4485))));
                      reg4504 <= reg4231;
                      reg4505 <= (8'ha6);
                    end
                end
              for (forvar4506 = (1'h0); (forvar4506 < (2'h3)); forvar4506 = (forvar4506 + (1'h1)))
                begin
                  if ((+reg4228[(1'h1):(1'h0)]))
                    begin
                      reg4507 <= (reg4418[(4'ha):(4'h8)] <<< $unsigned(((!(8'ha0)) << (~&(8'h9c)))));
                      reg4508 <= $unsigned(reg4255);
                    end
                  else
                    begin
                      reg4507 <= reg4334;
                      reg4508 <= (($unsigned({reg4237}) ?
                              $signed((^~reg4447)) : $unsigned((8'h9f))) ?
                          reg4326 : reg4240);
                    end
                  reg4509 <= reg4240[(3'h5):(1'h0)];
                  for (forvar4510 = (1'h0); (forvar4510 < (2'h2)); forvar4510 = (forvar4510 + (1'h1)))
                    begin
                      reg4511 <= (+$signed({reg4300[(2'h3):(2'h2)]}));
                      reg4512 <= reg4250;
                      reg4513 <= (8'h9d);
                    end
                end
              if ($signed(reg4364))
                begin
                  for (forvar4514 = (1'h0); (forvar4514 < (2'h3)); forvar4514 = (forvar4514 + (1'h1)))
                    begin
                      reg4515 <= {$signed({{reg4494}})};
                      reg4516 <= reg4499;
                      reg4517 <= $unsigned((~$unsigned(reg4471[(3'h4):(3'h4)])));
                      reg4518 <= reg4323[(4'ha):(3'h5)];
                    end
                  reg4519 <= $signed($signed($unsigned($unsigned((8'ha1)))));
                end
              else
                begin
                  reg4514 <= {($unsigned(forvar4510[(3'h6):(2'h2)]) ?
                          ((reg4388 || (8'had)) ?
                              reg4264 : $signed(reg4415)) : $unsigned($signed(reg4414)))};
                  if (reg4513)
                    begin
                      reg4515 <= $signed($unsigned(reg4389));
                      reg4516 <= $unsigned(reg4249[(3'h5):(2'h2)]);
                      reg4517 <= (8'ha5);
                      reg4518 <= (reg4313[(3'h5):(1'h1)] ?
                          (($unsigned(reg4276) ?
                              reg4444 : $unsigned(reg4398)) & {(wire4218 ?
                                  reg4343 : (8'ha7))}) : $unsigned({$unsigned(wire4218)}));
                    end
                  else
                    begin
                      reg4515 <= ((!($signed(reg4281) >>> (forvar4514 ^ (8'ha3)))) ?
                          $signed(reg4375[(3'h6):(2'h2)]) : reg4471[(3'h6):(3'h4)]);
                      reg4516 <= reg4367[(1'h0):(1'h0)];
                      reg4517 <= (reg4503[(2'h2):(1'h1)] ?
                          ($signed((reg4332 >= reg4290)) | {$signed(reg4435)}) : {$unsigned(reg4463[(1'h0):(1'h0)])});
                      reg4518 <= (((-$signed(reg4427)) ?
                          reg4460 : forvar4432[(3'h4):(1'h1)]) ^ {(8'hb3)});
                    end
                end
              for (forvar4520 = (1'h0); (forvar4520 < (2'h2)); forvar4520 = (forvar4520 + (1'h1)))
                begin
                  if ($signed((!$signed($signed((8'h9d))))))
                    begin
                      reg4521 <= (($unsigned((reg4267 - reg4405)) || (reg4274 ?
                              $signed((8'hb5)) : {(8'hb4)})) ?
                          $unsigned((~^forvar4458)) : reg4500);
                      reg4522 <= {(!({forvar4473} ?
                              reg4268[(4'h9):(3'h6)] : $unsigned(reg4502)))};
                      reg4523 <= (8'hae);
                      reg4524 <= $signed((({reg4510} ?
                              $signed(reg4268) : $unsigned(reg4279)) ?
                          reg4229 : (forvar4481 > forvar4440[(2'h3):(2'h3)])));
                    end
                  else
                    begin
                      reg4521 <= ($signed((|(reg4358 || forvar4510))) ^~ (-reg4504));
                    end
                  if ($signed(reg4508[(4'ha):(2'h3)]))
                    begin
                      reg4525 <= (&((+(forvar4458 >= reg4347)) ?
                          $unsigned(reg4351) : (~^reg4357)));
                      reg4526 <= (forvar4487 ?
                          reg4343[(2'h3):(2'h3)] : {(-(^~reg4468))});
                    end
                  else
                    begin
                      reg4525 <= reg4396[(3'h4):(2'h2)];
                      reg4526 <= $signed($signed($signed((reg4438 ?
                          reg4254 : reg4243))));
                      reg4527 <= (forvar4481 ?
                          reg4499 : reg4329[(1'h1):(1'h0)]);
                      reg4528 <= (({$signed(reg4254)} < (|$unsigned(reg4377))) ?
                          $unsigned(reg4441) : $unsigned($unsigned($signed(forvar4449))));
                    end
                  for (forvar4529 = (1'h0); (forvar4529 < (2'h3)); forvar4529 = (forvar4529 + (1'h1)))
                    begin
                      reg4530 <= ($unsigned(reg4226[(3'h6):(1'h1)]) * $signed(($signed(reg4369) ?
                          {reg4375} : (reg4222 ? wire4217 : reg4246))));
                    end
                end
            end
        end
      reg4531 <= {{((reg4367 ? reg4511 : forvar4452) ?
                  $signed(reg4337) : (reg4369 ? reg4279 : (8'h9e)))}};
    end
  assign wire4532 = $signed(((reg4428 ?
                            $unsigned((8'ha6)) : reg4422[(1'h0):(1'h0)]) ?
                        ((reg4234 ? reg4320 : reg4394) ?
                            (^~reg4342) : $signed(reg4269)) : (reg4343 ?
                            (~&reg4453) : (reg4479 ? reg4335 : reg4464))));
endmodule