(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param237 = (+(({(8'ha8)} || ((8'hb8) ~^ (8'h9f))) * (8'hba))))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'hacf):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire3;
  input wire signed [(5'h10):(1'h0)] wire2;
  input wire [(3'h6):(1'h0)] wire1;
  input wire [(4'hb):(1'h0)] wire0;
  wire signed [(3'h5):(1'h0)] wire236;
  wire [(4'ha):(1'h0)] wire235;
  wire signed [(2'h2):(1'h0)] wire234;
  wire signed [(5'h10):(1'h0)] wire233;
  reg [(4'hb):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg182 = (1'h0);
  reg [(4'ha):(1'h0)] reg170 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg169 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg158 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg150 = (1'h0);
  reg [(3'h6):(1'h0)] reg143 = (1'h0);
  reg [(3'h5):(1'h0)] reg137 = (1'h0);
  reg signed [(4'he):(1'h0)] reg135 = (1'h0);
  reg [(4'h8):(1'h0)] reg232 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg231 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg230 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg229 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg228 = (1'h0);
  reg [(4'hf):(1'h0)] reg225 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg227 = (1'h0);
  reg [(3'h4):(1'h0)] reg226 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg224 = (1'h0);
  reg [(4'hf):(1'h0)] reg223 = (1'h0);
  reg [(4'hb):(1'h0)] reg222 = (1'h0);
  reg signed [(4'he):(1'h0)] reg221 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg219 = (1'h0);
  reg [(3'h6):(1'h0)] reg218 = (1'h0);
  reg [(4'he):(1'h0)] reg217 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg215 = (1'h0);
  reg [(4'he):(1'h0)] reg214 = (1'h0);
  reg [(4'he):(1'h0)] reg212 = (1'h0);
  reg [(4'hb):(1'h0)] reg210 = (1'h0);
  reg [(3'h4):(1'h0)] reg209 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg208 = (1'h0);
  reg [(4'ha):(1'h0)] reg206 = (1'h0);
  reg [(2'h3):(1'h0)] reg204 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg202 = (1'h0);
  reg [(2'h2):(1'h0)] reg201 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg199 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg198 = (1'h0);
  reg [(2'h3):(1'h0)] reg196 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg195 = (1'h0);
  reg [(4'ha):(1'h0)] reg194 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg193 = (1'h0);
  reg [(4'h9):(1'h0)] reg192 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg191 = (1'h0);
  reg [(3'h4):(1'h0)] reg190 = (1'h0);
  reg [(4'hd):(1'h0)] reg189 = (1'h0);
  reg [(3'h5):(1'h0)] reg188 = (1'h0);
  reg [(5'h10):(1'h0)] reg187 = (1'h0);
  reg [(2'h2):(1'h0)] reg186 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg179 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg174 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg183 = (1'h0);
  reg [(2'h2):(1'h0)] reg181 = (1'h0);
  reg [(4'hb):(1'h0)] reg180 = (1'h0);
  reg [(4'hb):(1'h0)] reg178 = (1'h0);
  reg [(4'hf):(1'h0)] reg177 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg176 = (1'h0);
  reg [(3'h7):(1'h0)] reg175 = (1'h0);
  reg [(3'h4):(1'h0)] reg173 = (1'h0);
  reg [(4'hd):(1'h0)] reg172 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg171 = (1'h0);
  reg [(4'hb):(1'h0)] reg168 = (1'h0);
  reg [(3'h5):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg166 = (1'h0);
  reg [(3'h7):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg163 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg161 = (1'h0);
  reg [(4'h8):(1'h0)] reg157 = (1'h0);
  reg [(4'h8):(1'h0)] reg156 = (1'h0);
  reg signed [(4'he):(1'h0)] reg154 = (1'h0);
  reg [(4'h8):(1'h0)] reg153 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg152 = (1'h0);
  reg [(4'hf):(1'h0)] reg151 = (1'h0);
  reg signed [(4'he):(1'h0)] reg149 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg148 = (1'h0);
  reg [(4'h9):(1'h0)] reg145 = (1'h0);
  reg [(4'ha):(1'h0)] reg144 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg142 = (1'h0);
  reg [(4'hf):(1'h0)] reg140 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg139 = (1'h0);
  reg [(4'hd):(1'h0)] reg138 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg136 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg134 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg133 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg132 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg131 = (1'h0);
  reg [(2'h2):(1'h0)] reg130 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg128 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg127 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg126 = (1'h0);
  reg [(4'he):(1'h0)] reg124 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg125 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg123 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg121 = (1'h0);
  reg [(4'hf):(1'h0)] reg120 = (1'h0);
  reg [(4'hd):(1'h0)] reg119 = (1'h0);
  reg [(4'hd):(1'h0)] reg118 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg111 = (1'h0);
  reg [(2'h3):(1'h0)] reg117 = (1'h0);
  reg [(4'h8):(1'h0)] reg116 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg115 = (1'h0);
  reg [(2'h2):(1'h0)] reg114 = (1'h0);
  reg signed [(4'he):(1'h0)] reg113 = (1'h0);
  reg [(3'h7):(1'h0)] reg112 = (1'h0);
  reg [(4'hb):(1'h0)] reg110 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg109 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg108 = (1'h0);
  reg signed [(4'he):(1'h0)] reg107 = (1'h0);
  reg [(4'hb):(1'h0)] reg106 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg104 = (1'h0);
  reg [(5'h10):(1'h0)] reg103 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg86 = (1'h0);
  reg [(5'h10):(1'h0)] reg101 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg100 = (1'h0);
  reg [(3'h6):(1'h0)] reg99 = (1'h0);
  reg [(5'h10):(1'h0)] reg98 = (1'h0);
  reg [(2'h2):(1'h0)] reg94 = (1'h0);
  reg [(4'hb):(1'h0)] reg97 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg96 = (1'h0);
  reg [(4'he):(1'h0)] reg95 = (1'h0);
  reg [(5'h10):(1'h0)] reg93 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg92 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg90 = (1'h0);
  reg [(3'h7):(1'h0)] reg89 = (1'h0);
  reg [(4'he):(1'h0)] reg88 = (1'h0);
  reg [(4'h9):(1'h0)] reg87 = (1'h0);
  reg [(4'h8):(1'h0)] reg85 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg83 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg82 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg79 = (1'h0);
  reg [(4'hc):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg77 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg76 = (1'h0);
  reg [(4'hb):(1'h0)] reg75 = (1'h0);
  reg [(4'ha):(1'h0)] reg74 = (1'h0);
  reg signed [(4'he):(1'h0)] reg73 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg72 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg68 = (1'h0);
  reg [(4'he):(1'h0)] reg67 = (1'h0);
  reg [(4'hb):(1'h0)] reg65 = (1'h0);
  reg [(3'h5):(1'h0)] reg63 = (1'h0);
  reg [(4'ha):(1'h0)] reg58 = (1'h0);
  reg [(4'hb):(1'h0)] reg62 = (1'h0);
  reg [(4'hd):(1'h0)] reg61 = (1'h0);
  reg [(4'h9):(1'h0)] reg60 = (1'h0);
  reg [(3'h5):(1'h0)] reg59 = (1'h0);
  reg [(4'h9):(1'h0)] reg56 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg54 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg53 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg52 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg51 = (1'h0);
  reg [(4'hd):(1'h0)] reg50 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg49 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg48 = (1'h0);
  reg [(4'h9):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg42 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg38 = (1'h0);
  reg [(3'h6):(1'h0)] reg45 = (1'h0);
  reg [(4'ha):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg43 = (1'h0);
  reg [(4'h8):(1'h0)] reg41 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg40 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg39 = (1'h0);
  reg signed [(4'he):(1'h0)] reg37 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg36 = (1'h0);
  reg [(3'h7):(1'h0)] reg35 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg34 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5 = (1'h0);
  reg [(4'he):(1'h0)] reg15 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg12 = (1'h0);
  reg [(5'h10):(1'h0)] reg11 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg32 = (1'h0);
  reg [(2'h2):(1'h0)] reg31 = (1'h0);
  reg [(4'h8):(1'h0)] reg30 = (1'h0);
  reg [(3'h6):(1'h0)] reg29 = (1'h0);
  reg [(3'h7):(1'h0)] reg28 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg27 = (1'h0);
  reg [(4'hc):(1'h0)] reg26 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg23 = (1'h0);
  reg [(4'he):(1'h0)] reg22 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg21 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg18 = (1'h0);
  reg [(3'h7):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg16 = (1'h0);
  reg [(4'hb):(1'h0)] reg14 = (1'h0);
  reg [(3'h6):(1'h0)] reg13 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg10 = (1'h0);
  reg [(4'hf):(1'h0)] reg9 = (1'h0);
  reg [(4'hc):(1'h0)] reg8 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7 = (1'h0);
  reg [(4'hb):(1'h0)] reg6 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar191 = (1'h0);
  reg [(4'he):(1'h0)] forvar187 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar186 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar181 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar176 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar175 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar171 = (1'h0);
  reg [(4'hf):(1'h0)] forvar166 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar163 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar145 = (1'h0);
  reg [(3'h5):(1'h0)] forvar136 = (1'h0);
  reg [(4'hf):(1'h0)] forvar226 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar225 = (1'h0);
  reg [(4'he):(1'h0)] forvar220 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar216 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar213 = (1'h0);
  reg [(5'h10):(1'h0)] forvar211 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar207 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar205 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar203 = (1'h0);
  reg [(3'h7):(1'h0)] forvar200 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar197 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar185 = (1'h0);
  reg [(4'h8):(1'h0)] forvar177 = (1'h0);
  reg [(5'h10):(1'h0)] forvar182 = (1'h0);
  reg [(4'hb):(1'h0)] forvar179 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar174 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar170 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar169 = (1'h0);
  reg [(3'h7):(1'h0)] forvar165 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar160 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar159 = (1'h0);
  reg [(3'h7):(1'h0)] forvar158 = (1'h0);
  reg [(3'h7):(1'h0)] forvar155 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar150 = (1'h0);
  reg [(4'ha):(1'h0)] forvar147 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar146 = (1'h0);
  reg [(4'hf):(1'h0)] forvar143 = (1'h0);
  reg [(5'h10):(1'h0)] forvar141 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar137 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar135 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar131 = (1'h0);
  reg [(4'hd):(1'h0)] forvar125 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar129 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar124 = (1'h0);
  reg [(4'hc):(1'h0)] forvar121 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar110 = (1'h0);
  reg [(4'hf):(1'h0)] forvar111 = (1'h0);
  reg [(4'hf):(1'h0)] forvar105 = (1'h0);
  reg [(4'ha):(1'h0)] forvar102 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar96 = (1'h0);
  reg [(4'hb):(1'h0)] forvar94 = (1'h0);
  reg [(4'ha):(1'h0)] forvar91 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar86 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar81 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar71 = (1'h0);
  reg [(4'hb):(1'h0)] forvar70 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar66 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar64 = (1'h0);
  reg [(4'hd):(1'h0)] forvar61 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar58 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar57 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar47 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar39 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar34 = (1'h0);
  reg [(4'h9):(1'h0)] forvar42 = (1'h0);
  reg [(4'h9):(1'h0)] forvar38 = (1'h0);
  reg [(4'hb):(1'h0)] forvar33 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar13 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar8 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar25 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar24 = (1'h0);
  reg [(3'h4):(1'h0)] forvar20 = (1'h0);
  reg [(4'he):(1'h0)] forvar15 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar12 = (1'h0);
  reg [(3'h5):(1'h0)] forvar11 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4 = (1'h0);
  assign y = {wire236,
                 wire235,
                 wire234,
                 wire233,
                 reg185,
                 reg182,
                 reg170,
                 reg169,
                 reg158,
                 reg150,
                 reg143,
                 reg137,
                 reg135,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg225,
                 reg227,
                 reg226,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg219,
                 reg218,
                 reg217,
                 reg215,
                 reg214,
                 reg212,
                 reg210,
                 reg209,
                 reg208,
                 reg206,
                 reg204,
                 reg202,
                 reg201,
                 reg199,
                 reg198,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg179,
                 reg174,
                 reg184,
                 reg183,
                 reg181,
                 reg180,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg173,
                 reg172,
                 reg171,
                 reg168,
                 reg167,
                 reg166,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg157,
                 reg156,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg149,
                 reg148,
                 reg145,
                 reg144,
                 reg142,
                 reg140,
                 reg139,
                 reg138,
                 reg136,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg128,
                 reg127,
                 reg126,
                 reg124,
                 reg125,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg111,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg104,
                 reg103,
                 reg86,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg94,
                 reg97,
                 reg96,
                 reg95,
                 reg93,
                 reg92,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg69,
                 reg68,
                 reg67,
                 reg65,
                 reg63,
                 reg58,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg46,
                 reg42,
                 reg38,
                 reg45,
                 reg44,
                 reg43,
                 reg41,
                 reg40,
                 reg39,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg5,
                 reg15,
                 reg12,
                 reg11,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg23,
                 reg22,
                 reg21,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg14,
                 reg13,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 reg6,
                 forvar191,
                 forvar187,
                 forvar186,
                 forvar181,
                 forvar176,
                 forvar175,
                 forvar171,
                 forvar166,
                 forvar163,
                 forvar145,
                 forvar136,
                 forvar226,
                 forvar225,
                 forvar220,
                 forvar216,
                 forvar213,
                 forvar211,
                 forvar207,
                 forvar205,
                 forvar203,
                 forvar200,
                 forvar197,
                 forvar185,
                 forvar177,
                 forvar182,
                 forvar179,
                 forvar174,
                 forvar170,
                 forvar169,
                 forvar165,
                 forvar160,
                 forvar159,
                 forvar158,
                 forvar155,
                 forvar150,
                 forvar147,
                 forvar146,
                 forvar143,
                 forvar141,
                 forvar137,
                 forvar135,
                 forvar131,
                 forvar125,
                 forvar129,
                 forvar124,
                 forvar121,
                 forvar110,
                 forvar111,
                 forvar105,
                 forvar102,
                 forvar96,
                 forvar94,
                 forvar91,
                 forvar86,
                 forvar81,
                 forvar71,
                 forvar70,
                 forvar66,
                 forvar64,
                 forvar61,
                 forvar58,
                 forvar57,
                 forvar47,
                 forvar39,
                 forvar34,
                 forvar42,
                 forvar38,
                 forvar33,
                 forvar13,
                 forvar8,
                 forvar25,
                 forvar24,
                 forvar20,
                 forvar15,
                 forvar12,
                 forvar11,
                 forvar5,
                 forvar4,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (2'h3)); forvar4 = (forvar4 + (1'h1)))
        begin
          if ({(((~|wire1) ?
                  (wire0 ? wire1 : wire0) : (forvar4 ?
                      forvar4 : wire2)) || wire3)})
            begin
              for (forvar5 = (1'h0); (forvar5 < (2'h2)); forvar5 = (forvar5 + (1'h1)))
                begin
                  if ((((8'ha3) ?
                      $signed(forvar4) : (((8'hab) >> wire0) ?
                          forvar5 : (^wire3))) >>> wire1))
                    begin
                      reg6 <= (8'hb2);
                    end
                  else
                    begin
                      reg6 <= (~&wire3);
                    end
                  if ($signed((!forvar5)))
                    begin
                      reg7 <= (reg6[(4'hb):(1'h1)] | {$unsigned($signed(wire0))});
                      reg8 <= reg6;
                      reg9 <= $unsigned({$signed(reg8)});
                      reg10 <= $signed({reg8});
                    end
                  else
                    begin
                      reg7 <= (~$signed($signed($signed(reg8))));
                      reg8 <= (!forvar5[(3'h5):(2'h3)]);
                      reg9 <= {forvar5[(3'h5):(2'h2)]};
                    end
                end
              for (forvar11 = (1'h0); (forvar11 < (2'h2)); forvar11 = (forvar11 + (1'h1)))
                begin
                  for (forvar12 = (1'h0); (forvar12 < (2'h3)); forvar12 = (forvar12 + (1'h1)))
                    begin
                      reg13 <= $unsigned(({(~&forvar11)} * wire2[(3'h7):(2'h2)]));
                    end
                  reg14 <= (forvar4 ?
                      forvar4 : ($unsigned((^~forvar11)) ?
                          (-wire2[(3'h7):(2'h3)]) : $signed(reg6)));
                  for (forvar15 = (1'h0); (forvar15 < (1'h0)); forvar15 = (forvar15 + (1'h1)))
                    begin
                      reg16 <= reg13[(2'h3):(1'h0)];
                      reg17 <= reg8;
                      reg18 <= reg8[(4'hc):(2'h2)];
                      reg19 <= ($signed($unsigned((forvar4 ? reg6 : wire1))) ?
                          reg7 : $signed(((-reg9) == $unsigned(wire0))));
                    end
                  for (forvar20 = (1'h0); (forvar20 < (1'h0)); forvar20 = (forvar20 + (1'h1)))
                    begin
                      reg21 <= reg8;
                      reg22 <= reg9;
                      reg23 <= $signed($signed(reg9));
                    end
                end
              for (forvar24 = (1'h0); (forvar24 < (2'h3)); forvar24 = (forvar24 + (1'h1)))
                begin
                  for (forvar25 = (1'h0); (forvar25 < (2'h2)); forvar25 = (forvar25 + (1'h1)))
                    begin
                      reg26 <= {((forvar25 != (reg21 & reg10)) == $unsigned((reg21 <= wire0)))};
                      reg27 <= (^~$signed(($unsigned((8'h9d)) ?
                          (+(8'h9f)) : {wire3})));
                      reg28 <= reg9[(4'hf):(1'h1)];
                    end
                  if (reg13[(3'h4):(2'h3)])
                    begin
                      reg29 <= wire2[(2'h3):(1'h1)];
                      reg30 <= (8'hb3);
                      reg31 <= (~^$signed({(~&reg8)}));
                      reg32 <= (8'hba);
                    end
                  else
                    begin
                      reg29 <= reg17[(1'h0):(1'h0)];
                    end
                end
            end
          else
            begin
              if ($unsigned((!{reg18[(3'h5):(3'h5)]})))
                begin
                  for (forvar5 = (1'h0); (forvar5 < (1'h0)); forvar5 = (forvar5 + (1'h1)))
                    begin
                      reg6 <= $unsigned(reg6);
                      reg7 <= reg28;
                    end
                  for (forvar8 = (1'h0); (forvar8 < (1'h1)); forvar8 = (forvar8 + (1'h1)))
                    begin
                      reg9 <= (wire2[(3'h4):(1'h0)] ?
                          wire0 : (reg23[(3'h6):(1'h0)] >>> forvar24));
                      reg10 <= reg27[(1'h0):(1'h0)];
                      reg11 <= ((($signed(reg9) * reg7) | $unsigned({reg13})) ?
                          (~|($unsigned((8'hb2)) ?
                              $unsigned(reg13) : reg18)) : {{{forvar11}}});
                      reg12 <= (8'ha2);
                    end
                  for (forvar13 = (1'h0); (forvar13 < (2'h2)); forvar13 = (forvar13 + (1'h1)))
                    begin
                      reg14 <= (|($unsigned($signed(forvar11)) & $signed((+forvar24))));
                      reg15 <= forvar20;
                      reg16 <= {$unsigned($unsigned((-reg23)))};
                    end
                end
              else
                begin
                  if ((forvar13 ?
                      $unsigned((reg31 == $unsigned(reg30))) : (~^reg18)))
                    begin
                      reg5 <= $unsigned(reg21);
                      reg6 <= {{forvar24}};
                    end
                  else
                    begin
                      reg5 <= reg11;
                      reg6 <= $unsigned($unsigned($signed((wire1 + (8'ha9)))));
                      reg7 <= (^wire2[(4'hc):(2'h2)]);
                    end
                  if (($unsigned(reg7[(3'h5):(2'h3)]) ? forvar13 : wire0))
                    begin
                      reg8 <= reg29[(3'h5):(1'h0)];
                      reg9 <= reg32;
                    end
                  else
                    begin
                      reg8 <= $signed(reg31[(1'h0):(1'h0)]);
                    end
                  if (forvar25[(3'h5):(1'h1)])
                    begin
                      reg10 <= wire1[(2'h3):(1'h1)];
                      reg11 <= (8'hb5);
                      reg12 <= $unsigned((({reg17} || reg31) + reg9));
                      reg13 <= forvar15[(4'hc):(1'h1)];
                    end
                  else
                    begin
                      reg10 <= $signed((8'hb1));
                      reg11 <= {(!reg30[(2'h2):(1'h0)])};
                      reg12 <= (8'ha4);
                      reg13 <= (reg10[(4'hd):(2'h2)] > reg17);
                    end
                  if ($signed((~$signed(reg9[(3'h7):(3'h4)]))))
                    begin
                      reg14 <= $signed(($signed(reg17) > $signed(reg17[(3'h5):(3'h4)])));
                      reg15 <= wire0[(4'ha):(1'h1)];
                      reg16 <= reg21[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg14 <= reg23[(4'hb):(1'h1)];
                    end
                end
            end
          for (forvar33 = (1'h0); (forvar33 < (2'h3)); forvar33 = (forvar33 + (1'h1)))
            begin
              if (reg8[(3'h7):(3'h4)])
                begin
                  if (($signed(forvar15) ?
                      $unsigned($signed(forvar25)) : reg8[(4'h8):(1'h1)]))
                    begin
                      reg34 <= reg7;
                      reg35 <= ($signed(reg18[(1'h1):(1'h0)]) ?
                          forvar33[(3'h4):(1'h0)] : wire3[(1'h1):(1'h0)]);
                      reg36 <= (^~{$signed($signed((8'ha1)))});
                      reg37 <= (((((8'ha3) ? wire2 : (8'ha8)) ?
                                  reg11[(4'h8):(1'h1)] : (reg7 ?
                                      reg28 : reg15)) ?
                              forvar4[(2'h3):(2'h2)] : $unsigned(((8'ha8) ?
                                  reg36 : reg18))) ?
                          {reg16[(3'h4):(2'h3)]} : $unsigned((~|(reg5 ?
                              reg21 : forvar11))));
                    end
                  else
                    begin
                      reg34 <= reg30;
                      reg35 <= (~|{(reg36 ?
                              $signed(reg12) : $unsigned(reg29))});
                      reg36 <= $unsigned(reg28);
                    end
                  for (forvar38 = (1'h0); (forvar38 < (2'h3)); forvar38 = (forvar38 + (1'h1)))
                    begin
                      reg39 <= (8'ha9);
                      reg40 <= (!$signed(((reg8 <<< reg6) * forvar38)));
                      reg41 <= $signed($unsigned($signed($unsigned(reg26))));
                    end
                  for (forvar42 = (1'h0); (forvar42 < (2'h3)); forvar42 = (forvar42 + (1'h1)))
                    begin
                      reg43 <= $unsigned((~|(+reg28)));
                      reg44 <= reg19;
                      reg45 <= (($signed($signed(reg17)) ? (8'hac) : reg26) ?
                          $unsigned({$signed(forvar20)}) : reg5[(3'h4):(3'h4)]);
                    end
                end
              else
                begin
                  for (forvar34 = (1'h0); (forvar34 < (1'h0)); forvar34 = (forvar34 + (1'h1)))
                    begin
                      reg35 <= reg32[(4'hb):(3'h7)];
                      reg36 <= {((!{forvar15}) ?
                              reg14[(3'h5):(3'h5)] : ({reg15} >>> ((8'hae) - (8'hb1))))};
                      reg37 <= {(~|forvar20[(2'h3):(1'h1)])};
                      reg38 <= $unsigned((&($unsigned(reg28) ?
                          ((8'hb3) ? reg16 : forvar12) : $signed(reg18))));
                    end
                  for (forvar39 = (1'h0); (forvar39 < (2'h3)); forvar39 = (forvar39 + (1'h1)))
                    begin
                      reg40 <= $signed(reg19);
                      reg41 <= forvar33[(3'h4):(1'h0)];
                      reg42 <= ((!reg23) ?
                          (|$signed({reg12})) : ((~|(forvar13 | (8'hb7))) ?
                              reg37[(2'h3):(1'h1)] : ((forvar15 ~^ reg12) ^~ $unsigned(forvar15))));
                    end
                  reg43 <= reg39[(4'h9):(2'h2)];
                end
            end
          if ($signed(({forvar12[(2'h2):(2'h2)]} ?
              (^(reg19 ? reg39 : reg41)) : ($unsigned(wire0) ?
                  (reg16 ? reg8 : (8'ha2)) : reg9[(4'he):(4'hc)]))))
            begin
              reg46 <= forvar5;
              for (forvar47 = (1'h0); (forvar47 < (2'h2)); forvar47 = (forvar47 + (1'h1)))
                begin
                  reg48 <= (forvar24[(4'ha):(4'h9)] ^~ ((-$signed((8'ha1))) ?
                      forvar25 : reg16[(2'h2):(2'h2)]));
                  if ((8'had))
                    begin
                      reg49 <= reg12[(4'h9):(2'h3)];
                      reg50 <= $unsigned((!reg38));
                      reg51 <= ($signed(forvar25) ?
                          (-((&(8'hb5)) ? reg29 : $signed(reg22))) : (8'ha4));
                    end
                  else
                    begin
                      reg49 <= reg21;
                      reg50 <= ($unsigned((+$signed(reg26))) ?
                          reg26 : {$signed(reg21[(4'hd):(3'h6)])});
                      reg51 <= $unsigned((|forvar47[(1'h1):(1'h0)]));
                      reg52 <= reg6;
                    end
                  if (forvar39[(2'h3):(1'h1)])
                    begin
                      reg53 <= (8'ha5);
                      reg54 <= reg38;
                      reg55 <= (!forvar13[(1'h1):(1'h1)]);
                      reg56 <= $signed((|reg23[(4'hf):(3'h5)]));
                    end
                  else
                    begin
                      reg53 <= (+(+$signed($unsigned(forvar13))));
                    end
                end
            end
          else
            begin
              reg46 <= $unsigned({(~^$unsigned(wire0))});
            end
        end
      for (forvar57 = (1'h0); (forvar57 < (1'h1)); forvar57 = (forvar57 + (1'h1)))
        begin
          if ({(&$signed((-(8'hb6))))})
            begin
              if ($signed(((^~(reg42 ? reg32 : (8'hab))) ?
                  (reg51 ?
                      reg13 : (forvar33 ?
                          (8'ha0) : reg7)) : ((forvar24 | forvar39) >>> (reg18 * reg5)))))
                begin
                  for (forvar58 = (1'h0); (forvar58 < (1'h1)); forvar58 = (forvar58 + (1'h1)))
                    begin
                      reg59 <= $unsigned((forvar4 || $unsigned((reg15 ?
                          forvar38 : (8'h9f)))));
                      reg60 <= $unsigned((((^~reg40) ?
                              (reg50 ? (8'ha7) : reg48) : {reg27}) ?
                          $signed($signed(reg11)) : ({reg40} != reg28)));
                      reg61 <= (~|$signed(reg5));
                    end
                  reg62 <= ({(~|$unsigned(reg44))} ?
                      (|$signed((forvar57 | forvar38))) : ((&reg51) ^~ {(reg18 && reg55)}));
                end
              else
                begin
                  reg58 <= forvar25;
                end
            end
          else
            begin
              if (reg5)
                begin
                  reg58 <= $signed((~|$signed((~reg14))));
                end
              else
                begin
                  if ((((8'hb2) ? (-{reg8}) : $signed(reg59)) ?
                      $unsigned(((forvar47 ? forvar57 : reg21) ?
                          forvar11[(2'h3):(2'h3)] : (~^reg37))) : $signed(reg42)))
                    begin
                      reg58 <= $unsigned($unsigned(((~&(8'hb6)) ?
                          (reg62 < reg48) : $signed(reg60))));
                      reg59 <= reg35[(1'h1):(1'h0)];
                      reg60 <= (((reg59 ? reg55 : $unsigned(wire3)) ?
                          $unsigned(reg5) : forvar25[(4'he):(2'h2)]) + reg21);
                    end
                  else
                    begin
                      reg58 <= $signed($signed($signed((^~reg50))));
                      reg59 <= (((-((8'hb3) ^~ forvar39)) ?
                              (+(+(8'ha5))) : (reg46[(3'h4):(2'h2)] ^ (reg31 + forvar25))) ?
                          ((^reg11[(4'he):(3'h5)]) ?
                              ($unsigned(forvar24) ~^ reg54[(3'h7):(1'h1)]) : (!$unsigned(reg39))) : (reg9[(2'h2):(2'h2)] | (~|(~&reg11))));
                    end
                  for (forvar61 = (1'h0); (forvar61 < (2'h3)); forvar61 = (forvar61 + (1'h1)))
                    begin
                      reg62 <= reg39[(1'h1):(1'h1)];
                      reg63 <= reg39[(4'h9):(3'h6)];
                    end
                  for (forvar64 = (1'h0); (forvar64 < (1'h1)); forvar64 = (forvar64 + (1'h1)))
                    begin
                      reg65 <= reg13[(1'h0):(1'h0)];
                    end
                  for (forvar66 = (1'h0); (forvar66 < (1'h1)); forvar66 = (forvar66 + (1'h1)))
                    begin
                      reg67 <= ((($signed((8'hb3)) ?
                          $signed(reg6) : $unsigned(reg5)) == {$signed(forvar61)}) >= $signed((reg53 ?
                          reg28 : $unsigned(wire2))));
                      reg68 <= reg39[(2'h2):(1'h1)];
                      reg69 <= forvar42[(3'h4):(1'h1)];
                    end
                end
              for (forvar70 = (1'h0); (forvar70 < (1'h1)); forvar70 = (forvar70 + (1'h1)))
                begin
                  for (forvar71 = (1'h0); (forvar71 < (1'h1)); forvar71 = (forvar71 + (1'h1)))
                    begin
                      reg72 <= $signed(forvar42);
                      reg73 <= {((forvar5[(4'h9):(3'h4)] && forvar25) ?
                              (forvar15[(3'h5):(2'h3)] && $signed((8'ha9))) : ($signed(reg61) ?
                                  (reg37 == reg48) : {reg19}))};
                      reg74 <= (~&($signed($unsigned(reg69)) & (reg39 >>> (reg49 ~^ forvar4))));
                    end
                  if ((~(|(^~forvar39))))
                    begin
                      reg75 <= forvar64[(1'h1):(1'h1)];
                      reg76 <= $signed((((reg49 ? reg15 : reg51) ?
                          {(8'ha3)} : $unsigned(reg5)) == reg74[(2'h3):(1'h1)]));
                      reg77 <= (wire0 ?
                          {{reg67}} : (^(reg32[(1'h0):(1'h0)] ?
                              (reg29 ? forvar24 : reg27) : {(8'hab)})));
                    end
                  else
                    begin
                      reg75 <= ((^(^~(reg68 ?
                          reg17 : (8'hab)))) && $unsigned(reg68));
                      reg76 <= (({reg13[(1'h0):(1'h0)]} + ({reg30} ?
                              $signed(reg41) : $signed(reg76))) ?
                          (reg75[(2'h3):(2'h2)] << ((|reg50) ^~ $unsigned(reg8))) : {(+$signed(reg76))});
                      reg77 <= ((&((forvar70 >>> reg35) != $signed(reg9))) << ($signed((reg41 ^ reg61)) > reg10));
                    end
                  if (((($unsigned(forvar20) ?
                              (&forvar38) : forvar70[(4'h8):(1'h0)]) ?
                          (reg9 ?
                              $signed(reg5) : (forvar42 ?
                                  (8'hb8) : reg67)) : $signed($signed(reg17))) ?
                      (-wire1[(1'h1):(1'h1)]) : (reg76 ?
                          (^forvar34[(4'hb):(3'h4)]) : (8'hb3))))
                    begin
                      reg78 <= $unsigned($signed($signed($unsigned(reg6))));
                      reg79 <= {(+$unsigned(wire3[(3'h5):(2'h2)]))};
                      reg80 <= (forvar15[(4'ha):(3'h5)] ?
                          $signed($signed((reg76 ?
                              forvar42 : reg11))) : (~|forvar12));
                    end
                  else
                    begin
                      reg78 <= (^~(forvar39 <= (reg42 ?
                          $unsigned(forvar33) : $unsigned((8'ha1)))));
                    end
                  for (forvar81 = (1'h0); (forvar81 < (2'h2)); forvar81 = (forvar81 + (1'h1)))
                    begin
                      reg82 <= $unsigned((~$unsigned((^~(8'hb0)))));
                      reg83 <= $signed((~|(forvar81[(1'h0):(1'h0)] ?
                          reg75 : reg21[(3'h5):(3'h5)])));
                      reg84 <= (8'ha0);
                      reg85 <= wire0[(2'h3):(1'h0)];
                    end
                end
            end
          if ($unsigned($signed(((reg54 <= forvar5) ?
              forvar64[(3'h4):(3'h4)] : reg49[(3'h7):(3'h7)]))))
            begin
              for (forvar86 = (1'h0); (forvar86 < (2'h2)); forvar86 = (forvar86 + (1'h1)))
                begin
                  if ((~&($signed((~reg18)) ?
                      {(forvar70 ? wire1 : forvar71)} : $signed((forvar81 ?
                          reg76 : forvar70)))))
                    begin
                      reg87 <= forvar8[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg87 <= $signed((-reg52));
                      reg88 <= reg19;
                      reg89 <= ((((&(8'ha7)) > (reg56 * reg38)) || (forvar5[(3'h4):(2'h2)] <<< {forvar70})) <<< $unsigned(forvar42[(1'h1):(1'h0)]));
                      reg90 <= reg58[(4'h9):(4'h8)];
                    end
                  for (forvar91 = (1'h0); (forvar91 < (1'h1)); forvar91 = (forvar91 + (1'h1)))
                    begin
                      reg92 <= (+(~|reg56[(2'h3):(1'h1)]));
                      reg93 <= reg42;
                    end
                  for (forvar94 = (1'h0); (forvar94 < (2'h3)); forvar94 = (forvar94 + (1'h1)))
                    begin
                      reg95 <= $signed(reg22);
                      reg96 <= ((!forvar8) ?
                          (reg36 << $signed(reg55[(3'h5):(1'h1)])) : (~^forvar64[(1'h0):(1'h0)]));
                    end
                  reg97 <= $signed($unsigned(((reg73 ? forvar8 : reg92) ?
                      (wire1 ? forvar15 : reg62) : (~^reg87))));
                end
            end
          else
            begin
              if (reg23[(2'h2):(1'h1)])
                begin
                  for (forvar86 = (1'h0); (forvar86 < (2'h3)); forvar86 = (forvar86 + (1'h1)))
                    begin
                      reg87 <= $unsigned($unsigned($signed($signed(reg84))));
                      reg88 <= (+$signed(forvar71[(1'h0):(1'h0)]));
                      reg89 <= $unsigned(reg59[(2'h3):(1'h0)]);
                      reg90 <= $unsigned((~^(~^((8'h9e) || reg51))));
                    end
                  for (forvar91 = (1'h0); (forvar91 < (1'h0)); forvar91 = (forvar91 + (1'h1)))
                    begin
                      reg92 <= (~|({(!forvar66)} & $unsigned($unsigned(forvar24))));
                      reg93 <= ((8'hb5) ?
                          $signed(forvar66[(3'h4):(3'h4)]) : reg22[(2'h2):(2'h2)]);
                      reg94 <= (-reg6[(3'h7):(2'h3)]);
                      reg95 <= (&$unsigned((reg35[(1'h0):(1'h0)] ?
                          $unsigned(reg39) : reg89)));
                    end
                  for (forvar96 = (1'h0); (forvar96 < (2'h2)); forvar96 = (forvar96 + (1'h1)))
                    begin
                      reg97 <= {reg31[(2'h2):(1'h1)]};
                      reg98 <= wire3;
                      reg99 <= (^$signed((+(~|forvar61))));
                    end
                  if ($signed((8'hb1)))
                    begin
                      reg100 <= $signed($unsigned($unsigned(reg75)));
                      reg101 <= (((reg100 ~^ $unsigned(reg17)) ?
                          reg92[(4'h8):(1'h0)] : (!$unsigned(reg43))) > ({$unsigned(reg11)} >> $signed((+forvar91))));
                    end
                  else
                    begin
                      reg100 <= $signed(forvar58[(2'h3):(2'h2)]);
                      reg101 <= (8'hb0);
                    end
                end
              else
                begin
                  reg86 <= $signed(({$signed(forvar39)} ?
                      reg43 : reg92[(4'h8):(3'h6)]));
                  if (($signed($unsigned((~^reg8))) <<< forvar64[(2'h2):(2'h2)]))
                    begin
                      reg87 <= (($unsigned(reg22[(4'hb):(3'h5)]) ?
                              (~|reg74) : (+forvar42)) ?
                          (&reg95[(3'h6):(3'h6)]) : ($unsigned(reg99[(3'h5):(2'h3)]) >= $signed($signed(reg36))));
                      reg88 <= $unsigned(reg78[(4'ha):(4'ha)]);
                      reg89 <= reg87[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg87 <= $signed((|(!(reg8 * reg78))));
                      reg88 <= forvar91[(3'h4):(3'h4)];
                    end
                end
              for (forvar102 = (1'h0); (forvar102 < (1'h0)); forvar102 = (forvar102 + (1'h1)))
                begin
                  reg103 <= (~&(forvar64[(4'h8):(2'h3)] ?
                      $unsigned((8'hb0)) : $unsigned($unsigned(reg82))));
                  reg104 <= $unsigned((-$unsigned($unsigned(reg42))));
                  for (forvar105 = (1'h0); (forvar105 < (1'h0)); forvar105 = (forvar105 + (1'h1)))
                    begin
                      reg106 <= $unsigned(((wire1 ~^ (forvar38 ?
                          (8'h9f) : reg92)) > $signed({reg23})));
                      reg107 <= $signed((reg95[(2'h3):(2'h3)] ?
                          $unsigned(forvar4) : reg87[(2'h3):(1'h1)]));
                      reg108 <= (+({{(8'hb1)}} ?
                          {$unsigned((8'hab))} : forvar8));
                      reg109 <= forvar57[(3'h4):(1'h1)];
                    end
                end
              if (forvar47[(3'h7):(1'h0)])
                begin
                  reg110 <= $unsigned(($unsigned($signed(reg18)) ?
                      $signed($signed((8'hb8))) : ((forvar94 > reg87) ?
                          $signed(forvar12) : (reg48 ^ reg30))));
                  for (forvar111 = (1'h0); (forvar111 < (2'h2)); forvar111 = (forvar111 + (1'h1)))
                    begin
                      reg112 <= (8'hb3);
                      reg113 <= ({$signed($unsigned(reg48))} ?
                          $signed({forvar13}) : (^~(~&(8'ha4))));
                      reg114 <= $signed(($signed($unsigned(reg21)) ?
                          {(forvar102 ?
                                  forvar20 : reg38)} : forvar8[(3'h5):(3'h5)]));
                    end
                  reg115 <= wire3;
                  if ((8'ha9))
                    begin
                      reg116 <= wire1;
                      reg117 <= (&(8'hb7));
                    end
                  else
                    begin
                      reg116 <= (($unsigned(reg15[(4'h8):(2'h3)]) ?
                              forvar25 : ({wire3} ?
                                  (+forvar91) : $signed(forvar33))) ?
                          (reg109[(2'h2):(1'h1)] >= (8'had)) : wire3[(2'h3):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar110 = (1'h0); (forvar110 < (2'h3)); forvar110 = (forvar110 + (1'h1)))
                    begin
                      reg111 <= $signed({forvar11[(1'h0):(1'h0)]});
                      reg112 <= (8'hb0);
                      reg113 <= reg7;
                    end
                  if ({($signed($signed((8'ha4))) ?
                          $signed((reg85 ~^ reg38)) : reg101)})
                    begin
                      reg114 <= reg58[(1'h0):(1'h0)];
                      reg115 <= {(!((reg22 ?
                              forvar34 : reg53) == ((8'ha9) >>> (8'hb6))))};
                      reg116 <= (^(reg114 ? reg32 : $signed(forvar81)));
                      reg117 <= $unsigned(reg107);
                    end
                  else
                    begin
                      reg114 <= $unsigned(reg82[(3'h4):(1'h0)]);
                    end
                  if ((8'h9f))
                    begin
                      reg118 <= $unsigned(($signed(reg55) | $unsigned((reg107 ?
                          reg77 : forvar81))));
                    end
                  else
                    begin
                      reg118 <= $signed(forvar39);
                      reg119 <= $signed((((reg103 ?
                          reg75 : reg82) & reg88[(4'hd):(2'h2)]) - ((forvar24 ?
                          forvar12 : (8'hb8)) != (reg117 <= forvar15))));
                      reg120 <= ((~(((8'hb0) ? reg79 : reg51) || (reg87 ?
                          (8'hb7) : reg48))) >> $signed($unsigned($unsigned(forvar94))));
                    end
                end
            end
          if (reg106)
            begin
              if (({reg112[(1'h1):(1'h1)]} ?
                  ($unsigned(reg77) ?
                      (((8'hb9) - reg61) == reg89) : $unsigned((8'ha6))) : $unsigned($unsigned(reg12))))
                begin
                  reg121 <= ($signed(({reg77} ?
                          $signed(reg8) : ((8'haa) ? reg23 : reg8))) ?
                      {$signed($unsigned(reg87))} : (reg93 ?
                          reg60 : reg21[(2'h3):(1'h1)]));
                end
              else
                begin
                  for (forvar121 = (1'h0); (forvar121 < (1'h1)); forvar121 = (forvar121 + (1'h1)))
                    begin
                      reg122 <= (~|{forvar94});
                    end
                  reg123 <= reg63[(1'h0):(1'h0)];
                  for (forvar124 = (1'h0); (forvar124 < (1'h0)); forvar124 = (forvar124 + (1'h1)))
                    begin
                      reg125 <= $signed((((^~reg48) ?
                          reg44 : reg119) == {reg22}));
                    end
                end
            end
          else
            begin
              if ($unsigned({($unsigned(forvar13) && (^~reg62))}))
                begin
                  for (forvar121 = (1'h0); (forvar121 < (1'h0)); forvar121 = (forvar121 + (1'h1)))
                    begin
                      reg122 <= wire3;
                      reg123 <= ((|(~^(reg54 ?
                          reg109 : forvar66))) >>> reg17[(3'h7):(1'h1)]);
                      reg124 <= ({(&{reg51})} ^~ (reg85[(3'h7):(3'h6)] ?
                          (~|wire0[(2'h2):(1'h0)]) : forvar71[(4'hc):(4'hc)]));
                      reg125 <= $unsigned(reg28[(3'h6):(2'h3)]);
                    end
                  if ({$signed((!$signed(reg78)))})
                    begin
                      reg126 <= reg6[(3'h4):(1'h0)];
                      reg127 <= (reg37[(4'he):(1'h0)] ^~ ($signed($signed(reg87)) >> ((+reg32) ?
                          forvar110[(4'ha):(4'h8)] : forvar110)));
                    end
                  else
                    begin
                      reg126 <= (forvar61 < reg52[(1'h1):(1'h0)]);
                      reg127 <= ((reg65[(2'h3):(1'h1)] >>> $signed($signed(reg74))) <<< (^$signed($unsigned(reg116))));
                      reg128 <= forvar121;
                    end
                  for (forvar129 = (1'h0); (forvar129 < (1'h1)); forvar129 = (forvar129 + (1'h1)))
                    begin
                      reg130 <= $unsigned(reg29[(3'h4):(2'h2)]);
                      reg131 <= $signed(reg119[(2'h3):(2'h3)]);
                    end
                end
              else
                begin
                  if (reg108[(1'h1):(1'h0)])
                    begin
                      reg121 <= $unsigned((^reg99[(2'h2):(1'h0)]));
                      reg122 <= $signed({(-$signed(reg75))});
                    end
                  else
                    begin
                      reg121 <= (reg82[(3'h6):(2'h3)] ?
                          ($unsigned(((8'hac) ? forvar71 : reg96)) <= ((reg80 ?
                                  reg8 : reg96) ?
                              $unsigned(forvar70) : {forvar70})) : (~($signed(reg32) ?
                              (!reg35) : $signed(reg17))));
                      reg122 <= $unsigned(reg31);
                      reg123 <= reg106;
                      reg124 <= $signed(({(forvar24 & reg98)} ?
                          ({reg22} != reg98[(2'h2):(2'h2)]) : ($signed((8'ha4)) ?
                              reg83[(4'h9):(3'h5)] : reg26[(1'h1):(1'h0)])));
                    end
                  for (forvar125 = (1'h0); (forvar125 < (1'h0)); forvar125 = (forvar125 + (1'h1)))
                    begin
                      reg126 <= reg67[(1'h0):(1'h0)];
                      reg127 <= (((8'ha2) ?
                              ((8'h9d) ?
                                  forvar110[(2'h2):(2'h2)] : ((8'h9c) ~^ (8'haa))) : ((forvar61 <= forvar42) ?
                                  (forvar47 >= reg119) : $unsigned(reg44))) ?
                          $signed((~|$unsigned(reg107))) : {$unsigned(forvar96[(1'h0):(1'h0)])});
                      reg128 <= forvar25[(4'h8):(3'h6)];
                    end
                  for (forvar129 = (1'h0); (forvar129 < (2'h3)); forvar129 = (forvar129 + (1'h1)))
                    begin
                      reg130 <= ($signed($unsigned(reg14)) ^ (({forvar111} ^ ((8'haa) == forvar86)) ?
                          (8'ha4) : forvar20[(1'h0):(1'h0)]));
                    end
                  for (forvar131 = (1'h0); (forvar131 < (1'h1)); forvar131 = (forvar131 + (1'h1)))
                    begin
                      reg132 <= ((reg92[(4'h9):(2'h3)] ?
                              reg53[(3'h7):(1'h1)] : ($unsigned(reg46) > reg32[(2'h3):(1'h0)])) ?
                          $unsigned(reg111) : {reg106});
                      reg133 <= (-$unsigned(((|reg40) ?
                          reg65[(1'h0):(1'h0)] : reg22[(4'hb):(4'h8)])));
                    end
                end
              reg134 <= ((((&reg7) ? $unsigned((8'haf)) : $unsigned(reg52)) ?
                  $unsigned($unsigned(forvar4)) : ($signed(reg77) && $signed(reg49))) - ((~|reg127) ?
                  reg103 : $signed((forvar125 ? reg113 : (8'hb4)))));
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg110)
        begin
          for (forvar135 = (1'h0); (forvar135 < (1'h0)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 <= wire3;
              if ((reg60[(1'h0):(1'h0)] || (|(reg48[(1'h0):(1'h0)] ?
                  $unsigned((8'ha4)) : reg30))))
                begin
                  for (forvar137 = (1'h0); (forvar137 < (1'h1)); forvar137 = (forvar137 + (1'h1)))
                    begin
                      reg138 <= (^((^(reg83 ? reg76 : reg56)) ?
                          ((reg95 > reg40) > $unsigned(reg49)) : $signed(((8'ha8) & forvar135))));
                      reg139 <= ($signed($unsigned(reg22)) ?
                          $signed(($signed(reg9) >> $unsigned(reg106))) : (reg41[(1'h1):(1'h0)] & $unsigned({reg124})));
                    end
                end
              else
                begin
                  for (forvar137 = (1'h0); (forvar137 < (1'h0)); forvar137 = (forvar137 + (1'h1)))
                    begin
                      reg138 <= (+(8'hb4));
                      reg139 <= reg26[(4'hb):(4'ha)];
                      reg140 <= reg77;
                    end
                  for (forvar141 = (1'h0); (forvar141 < (1'h1)); forvar141 = (forvar141 + (1'h1)))
                    begin
                      reg142 <= $signed($unsigned(((8'ha6) < reg17)));
                    end
                  for (forvar143 = (1'h0); (forvar143 < (1'h1)); forvar143 = (forvar143 + (1'h1)))
                    begin
                      reg144 <= $unsigned({(((8'hba) ? reg28 : (8'hae)) ?
                              reg44[(4'h8):(3'h7)] : $unsigned(reg124))});
                      reg145 <= ((-(reg58[(3'h7):(1'h0)] < $unsigned((8'ha6)))) ^ ($unsigned($signed(reg16)) - wire1));
                    end
                end
              for (forvar146 = (1'h0); (forvar146 < (1'h0)); forvar146 = (forvar146 + (1'h1)))
                begin
                  for (forvar147 = (1'h0); (forvar147 < (1'h1)); forvar147 = (forvar147 + (1'h1)))
                    begin
                      reg148 <= ({$signed(reg119[(2'h3):(2'h2)])} ?
                          $signed(reg6[(4'h9):(2'h2)]) : $unsigned($unsigned(reg110[(2'h2):(1'h0)])));
                      reg149 <= {(!reg18)};
                    end
                end
              for (forvar150 = (1'h0); (forvar150 < (2'h2)); forvar150 = (forvar150 + (1'h1)))
                begin
                  if ($signed((({reg114} ?
                      $signed((8'h9c)) : reg121[(2'h3):(2'h2)]) ^~ reg148[(2'h2):(1'h0)])))
                    begin
                      reg151 <= $signed($unsigned(reg21[(2'h3):(2'h3)]));
                      reg152 <= reg84;
                    end
                  else
                    begin
                      reg151 <= ((~forvar146) ~^ $unsigned((reg26 * reg120)));
                      reg152 <= $signed(($signed((reg10 ?
                          reg62 : reg53)) == (reg69 >> {reg50})));
                    end
                  reg153 <= reg128;
                  if ($signed($unsigned($unsigned((|reg67)))))
                    begin
                      reg154 <= $signed(reg114);
                    end
                  else
                    begin
                      reg154 <= $signed(((&(reg65 != reg21)) * $unsigned((reg111 ?
                          (8'hb0) : reg116))));
                    end
                  for (forvar155 = (1'h0); (forvar155 < (2'h2)); forvar155 = (forvar155 + (1'h1)))
                    begin
                      reg156 <= $unsigned((forvar146[(3'h5):(2'h3)] ?
                          ($unsigned(reg122) ?
                              reg36 : $unsigned(reg6)) : (reg72 ?
                              reg51 : $signed(reg14))));
                      reg157 <= ((-((reg106 ^~ reg149) ?
                              $signed(reg156) : {reg111})) ?
                          $signed($signed({(8'hb5)})) : $unsigned(((8'hb0) >= (-reg6))));
                    end
                end
            end
          for (forvar158 = (1'h0); (forvar158 < (1'h0)); forvar158 = (forvar158 + (1'h1)))
            begin
              for (forvar159 = (1'h0); (forvar159 < (2'h3)); forvar159 = (forvar159 + (1'h1)))
                begin
                  for (forvar160 = (1'h0); (forvar160 < (2'h2)); forvar160 = (forvar160 + (1'h1)))
                    begin
                      reg161 <= (($unsigned((wire3 ^~ reg52)) * forvar146[(1'h1):(1'h1)]) ?
                          ({(reg83 && reg120)} ?
                              $unsigned($unsigned(reg92)) : reg114[(2'h2):(2'h2)]) : reg145[(3'h4):(3'h4)]);
                      reg162 <= {$signed($signed($signed(reg68)))};
                      reg163 <= reg16;
                      reg164 <= (-(-(reg92[(4'he):(4'ha)] == reg28[(2'h3):(1'h0)])));
                    end
                  for (forvar165 = (1'h0); (forvar165 < (2'h2)); forvar165 = (forvar165 + (1'h1)))
                    begin
                      reg166 <= (($signed(reg36[(2'h3):(1'h1)]) & (reg9[(2'h2):(1'h0)] >> $signed(reg98))) ?
                          reg125 : $signed(reg157));
                    end
                  reg167 <= $unsigned((reg53[(3'h7):(1'h0)] ?
                      wire3 : reg94[(1'h1):(1'h0)]));
                end
              reg168 <= (+reg164[(3'h4):(2'h3)]);
            end
          for (forvar169 = (1'h0); (forvar169 < (2'h2)); forvar169 = (forvar169 + (1'h1)))
            begin
              if ($unsigned($signed($signed($unsigned(reg10)))))
                begin
                  for (forvar170 = (1'h0); (forvar170 < (2'h3)); forvar170 = (forvar170 + (1'h1)))
                    begin
                      reg171 <= (reg126 || $signed((8'ha6)));
                      reg172 <= {((reg117[(2'h2):(2'h2)] || $unsigned(reg11)) * reg111)};
                      reg173 <= {(((^~reg168) - (reg112 ? reg5 : (8'had))) ?
                              (reg59 ?
                                  forvar170[(3'h7):(3'h7)] : {reg7}) : reg17[(2'h3):(2'h2)])};
                    end
                  for (forvar174 = (1'h0); (forvar174 < (1'h0)); forvar174 = (forvar174 + (1'h1)))
                    begin
                      reg175 <= forvar169;
                      reg176 <= {(((reg72 <= reg171) >> reg167[(2'h2):(1'h1)]) ?
                              reg37 : $signed(reg149[(4'h8):(3'h6)]))};
                      reg177 <= $signed(reg161);
                      reg178 <= ((((!reg154) < (reg56 ? reg86 : reg28)) ?
                          (~&(reg37 ? reg50 : (8'hb7))) : $unsigned((reg88 ?
                              reg55 : reg76))) * (~&$signed(((8'hae) >>> reg35))));
                    end
                  for (forvar179 = (1'h0); (forvar179 < (1'h1)); forvar179 = (forvar179 + (1'h1)))
                    begin
                      reg180 <= (~^$unsigned(reg41));
                      reg181 <= ({((^reg53) ?
                                  (reg154 || reg68) : (reg11 <<< reg88))} ?
                          $signed((~&forvar170[(4'h8):(2'h2)])) : reg8[(1'h1):(1'h1)]);
                    end
                  for (forvar182 = (1'h0); (forvar182 < (1'h0)); forvar182 = (forvar182 + (1'h1)))
                    begin
                      reg183 <= ((-{$signed(reg78)}) >> reg80[(1'h1):(1'h0)]);
                      reg184 <= reg121[(4'hf):(3'h5)];
                    end
                end
              else
                begin
                  for (forvar170 = (1'h0); (forvar170 < (2'h3)); forvar170 = (forvar170 + (1'h1)))
                    begin
                      reg171 <= $signed((reg44[(3'h4):(1'h1)] >>> reg180));
                      reg172 <= (((-(reg40 || reg6)) ?
                          reg92[(3'h6):(1'h1)] : $unsigned((+reg53))) - ($signed((|reg67)) ?
                          {forvar137[(1'h1):(1'h1)]} : $unsigned({(8'ha4)})));
                      reg173 <= (~&forvar146);
                      reg174 <= reg65[(4'hb):(4'h9)];
                    end
                  if ((~&reg55[(3'h7):(3'h6)]))
                    begin
                      reg175 <= reg83;
                      reg176 <= $signed((8'ha2));
                    end
                  else
                    begin
                      reg175 <= (^(^(reg180[(1'h1):(1'h1)] << reg73[(3'h5):(2'h2)])));
                      reg176 <= $signed((((^~forvar141) > (reg117 ?
                              reg164 : reg108)) ?
                          reg22[(2'h3):(2'h2)] : (~^$signed(reg55))));
                    end
                  for (forvar177 = (1'h0); (forvar177 < (2'h3)); forvar177 = (forvar177 + (1'h1)))
                    begin
                      reg178 <= (((~&(reg38 & (8'hb0))) ?
                          $signed($signed(reg154)) : {(reg16 ?
                                  reg126 : (8'hb5))}) >> reg78);
                      reg179 <= ((^(forvar141[(4'h9):(3'h4)] == (~^reg15))) ?
                          forvar137 : {((+reg183) ?
                                  (^~reg15) : $unsigned(reg171))});
                      reg180 <= reg13;
                    end
                end
              for (forvar185 = (1'h0); (forvar185 < (2'h3)); forvar185 = (forvar185 + (1'h1)))
                begin
                  if ({reg87})
                    begin
                      reg186 <= (^reg72);
                    end
                  else
                    begin
                      reg186 <= $signed((+$signed($signed(reg100))));
                      reg187 <= (reg18 ?
                          ($signed(reg167) != (~|(reg126 ?
                              reg132 : reg126))) : (|reg172));
                    end
                  if ({reg41[(3'h4):(3'h4)]})
                    begin
                      reg188 <= reg41[(4'h8):(2'h2)];
                      reg189 <= (reg120 >>> $signed((^~reg56[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg188 <= reg49;
                      reg189 <= $unsigned(forvar169);
                      reg190 <= reg34[(3'h6):(2'h3)];
                      reg191 <= $signed({(~&(!reg189))});
                    end
                  reg192 <= $unsigned($signed(({reg65} != (8'hae))));
                  if ((^(|reg124[(4'he):(4'hb)])))
                    begin
                      reg193 <= $signed((~|reg86[(3'h7):(3'h6)]));
                      reg194 <= reg134[(2'h3):(2'h2)];
                      reg195 <= $unsigned(reg178[(3'h7):(3'h5)]);
                      reg196 <= $unsigned(((8'h9e) & $signed((reg184 ?
                          reg187 : (8'ha5)))));
                    end
                  else
                    begin
                      reg193 <= ($signed($unsigned(reg133[(3'h6):(3'h5)])) ?
                          ($unsigned((reg95 ? reg175 : reg171)) ?
                              (reg54 ?
                                  (forvar170 ? reg145 : reg27) : (reg82 ?
                                      reg117 : reg49)) : ((reg115 == reg30) >>> $unsigned((8'hb5)))) : (-((reg67 ?
                              reg104 : reg154) << reg118)));
                      reg194 <= {(((reg62 ? reg6 : reg36) << (reg72 ?
                              (8'ha6) : forvar137)) << $signed((reg123 == reg130)))};
                      reg195 <= (+{forvar135});
                      reg196 <= reg43[(2'h3):(2'h2)];
                    end
                end
              for (forvar197 = (1'h0); (forvar197 < (2'h3)); forvar197 = (forvar197 + (1'h1)))
                begin
                  reg198 <= (((8'hb3) ?
                          ((reg157 ?
                              forvar185 : wire2) >> $signed(reg37)) : (((8'hab) ?
                                  forvar141 : (8'h9c)) ?
                              (&forvar177) : reg118)) ?
                      reg49[(4'h9):(3'h5)] : ((reg104[(2'h2):(1'h1)] >>> {(8'ha3)}) == reg175));
                  reg199 <= reg32;
                  for (forvar200 = (1'h0); (forvar200 < (2'h2)); forvar200 = (forvar200 + (1'h1)))
                    begin
                      reg201 <= ((&reg189) ?
                          ($unsigned(reg38) ? reg174 : reg60) : reg58);
                    end
                  reg202 <= (($unsigned(((8'ha9) > reg10)) ^~ (reg180 + reg173)) ?
                      $signed((|(^~reg76))) : reg52);
                end
            end
          for (forvar203 = (1'h0); (forvar203 < (1'h0)); forvar203 = (forvar203 + (1'h1)))
            begin
              reg204 <= reg87[(4'h8):(3'h5)];
              for (forvar205 = (1'h0); (forvar205 < (1'h0)); forvar205 = (forvar205 + (1'h1)))
                begin
                  reg206 <= $signed($unsigned(reg56));
                  for (forvar207 = (1'h0); (forvar207 < (2'h2)); forvar207 = (forvar207 + (1'h1)))
                    begin
                      reg208 <= ({((8'h9f) ?
                                  $signed((8'hac)) : $signed(reg55))} ?
                          (reg12[(3'h7):(2'h3)] ?
                              reg38 : reg122) : ((&$signed(reg172)) ?
                              $unsigned(reg61) : forvar182));
                      reg209 <= ({$unsigned($signed(forvar205))} ?
                          (+($signed(reg22) ?
                              reg188[(1'h1):(1'h0)] : (~^reg178))) : ((reg156 > $signed(reg134)) ?
                              reg140 : $signed($unsigned(reg59))));
                      reg210 <= ($signed((reg117 || $signed(reg77))) ?
                          forvar147[(2'h3):(2'h2)] : $signed($unsigned((reg154 ?
                              reg16 : reg184))));
                    end
                  for (forvar211 = (1'h0); (forvar211 < (1'h1)); forvar211 = (forvar211 + (1'h1)))
                    begin
                      reg212 <= (^~(~reg166[(4'hf):(4'h9)]));
                    end
                end
              for (forvar213 = (1'h0); (forvar213 < (1'h0)); forvar213 = (forvar213 + (1'h1)))
                begin
                  if ($unsigned(reg23[(3'h5):(2'h3)]))
                    begin
                      reg214 <= reg19;
                      reg215 <= reg120;
                    end
                  else
                    begin
                      reg214 <= $signed({reg23});
                      reg215 <= reg130;
                    end
                  for (forvar216 = (1'h0); (forvar216 < (2'h3)); forvar216 = (forvar216 + (1'h1)))
                    begin
                      reg217 <= $unsigned((({reg48} ?
                          $signed(reg157) : {reg194}) || $signed((8'hb1))));
                      reg218 <= $unsigned($signed($signed({reg100})));
                      reg219 <= reg100;
                    end
                  for (forvar220 = (1'h0); (forvar220 < (1'h1)); forvar220 = (forvar220 + (1'h1)))
                    begin
                      reg221 <= reg93[(4'hc):(4'hc)];
                      reg222 <= $signed($signed(((reg78 ?
                          (8'hb7) : (8'hb4)) * (forvar177 ? reg175 : reg52))));
                      reg223 <= (((-(reg72 >> forvar177)) << ($signed((8'haa)) ?
                          (reg188 ~^ wire0) : (8'hb6))) >= reg214[(4'hd):(3'h7)]);
                      reg224 <= (!{$signed(((8'h9c) ? reg46 : reg85))});
                    end
                end
              if ($signed(reg61[(4'hb):(3'h7)]))
                begin
                  for (forvar225 = (1'h0); (forvar225 < (1'h0)); forvar225 = (forvar225 + (1'h1)))
                    begin
                      reg226 <= (-reg40[(4'h9):(3'h7)]);
                      reg227 <= forvar207;
                    end
                end
              else
                begin
                  reg225 <= reg195[(4'h9):(1'h0)];
                  for (forvar226 = (1'h0); (forvar226 < (2'h3)); forvar226 = (forvar226 + (1'h1)))
                    begin
                      reg227 <= ((8'h9e) ?
                          (($signed(reg48) ?
                              reg195[(4'h9):(3'h5)] : forvar226[(4'hd):(4'hb)]) & {(forvar203 > reg8)}) : $signed($signed({reg161})));
                      reg228 <= $signed((forvar165 ?
                          (~reg92[(4'hb):(4'h9)]) : $unsigned(reg97[(4'ha):(3'h6)])));
                      reg229 <= (^~reg34[(4'ha):(3'h6)]);
                    end
                  if ($signed(reg113[(4'h8):(4'h8)]))
                    begin
                      reg230 <= reg6[(1'h1):(1'h0)];
                      reg231 <= (+reg175);
                    end
                  else
                    begin
                      reg230 <= reg212;
                      reg231 <= $unsigned($unsigned((reg109 >>> reg69[(1'h1):(1'h0)])));
                      reg232 <= $unsigned($signed(forvar185[(3'h6):(3'h4)]));
                    end
                end
            end
        end
      else
        begin
          if ((($unsigned(reg195[(4'hc):(4'h9)]) ?
                  (~|((8'ha1) ? reg126 : reg176)) : reg133[(1'h0):(1'h0)]) ?
              reg68 : forvar146[(1'h0):(1'h0)]))
            begin
              reg135 <= {((~&(|reg107)) ? $signed($signed(reg48)) : reg94)};
              if (reg218[(3'h5):(3'h5)])
                begin
                  reg136 <= reg23[(4'hf):(2'h3)];
                  reg137 <= (^~($unsigned(reg50) ? reg101 : reg104));
                end
              else
                begin
                  for (forvar136 = (1'h0); (forvar136 < (1'h1)); forvar136 = (forvar136 + (1'h1)))
                    begin
                      reg137 <= reg11[(3'h7):(2'h2)];
                      reg138 <= (|($signed((!(8'ha7))) ~^ reg56[(2'h2):(1'h1)]));
                      reg139 <= ((($unsigned(reg111) & reg124) >>> $unsigned(reg157)) ?
                          reg130[(2'h2):(1'h0)] : ($signed(forvar226[(3'h6):(3'h4)]) ?
                              ((reg219 + reg5) >= (reg161 ?
                                  reg126 : reg175)) : (~&(reg17 ~^ forvar177))));
                      reg140 <= (8'h9d);
                    end
                  for (forvar141 = (1'h0); (forvar141 < (1'h1)); forvar141 = (forvar141 + (1'h1)))
                    begin
                      reg142 <= (reg14[(3'h5):(3'h5)] >> (-reg89[(1'h0):(1'h0)]));
                      reg143 <= (reg173 ?
                          {((^(8'h9e)) ^ $signed(reg35))} : $unsigned({{reg31}}));
                    end
                end
              reg144 <= $signed($signed(((+(8'hb5)) ?
                  (reg226 ? (8'hb0) : (8'ha7)) : $unsigned((8'hae)))));
            end
          else
            begin
              reg135 <= (!(8'haf));
            end
          for (forvar145 = (1'h0); (forvar145 < (2'h3)); forvar145 = (forvar145 + (1'h1)))
            begin
              for (forvar146 = (1'h0); (forvar146 < (2'h3)); forvar146 = (forvar146 + (1'h1)))
                begin
                  for (forvar147 = (1'h0); (forvar147 < (2'h2)); forvar147 = (forvar147 + (1'h1)))
                    begin
                      reg148 <= $signed(($signed((^~reg41)) ?
                          (^~$signed(reg72)) : $unsigned((reg112 ?
                              forvar174 : reg6))));
                      reg149 <= $unsigned(reg192);
                      reg150 <= $signed($signed(reg120));
                    end
                  reg151 <= ((reg63[(1'h0):(1'h0)] ^~ $unsigned($signed((8'ha4)))) ?
                      forvar200[(1'h0):(1'h0)] : ($unsigned($unsigned(reg179)) ?
                          $unsigned((~reg59)) : (^$unsigned(reg85))));
                  if (reg139)
                    begin
                      reg152 <= ({(((8'hb3) ? reg100 : reg73) ?
                              (reg69 - reg142) : $unsigned(reg191))} <= (((reg90 <<< (8'hb1)) >> (reg60 && reg45)) <<< $unsigned($unsigned(reg13))));
                      reg153 <= ($signed(reg84[(3'h5):(2'h2)]) ?
                          (((~&forvar137) ^ (reg202 < (8'ha1))) ?
                              $signed($unsigned(reg215)) : $signed((reg96 ?
                                  forvar159 : reg79))) : (reg23 ^ (^~(reg103 || (8'hb4)))));
                      reg154 <= $unsigned($signed($unsigned($unsigned(reg67))));
                    end
                  else
                    begin
                      reg152 <= forvar170[(4'hc):(2'h2)];
                      reg153 <= reg151[(3'h7):(2'h3)];
                      reg154 <= reg95;
                    end
                  for (forvar155 = (1'h0); (forvar155 < (2'h2)); forvar155 = (forvar155 + (1'h1)))
                    begin
                      reg156 <= reg219;
                      reg157 <= ($signed(((reg113 ? reg96 : reg5) ?
                              (reg51 ~^ reg229) : $unsigned((8'h9d)))) ?
                          ($unsigned(reg59) ?
                              (^{(8'hb5)}) : ($unsigned(reg21) ?
                                  $signed(reg56) : (~^reg144))) : $signed(forvar207[(4'hb):(3'h6)]));
                      reg158 <= {reg208};
                    end
                end
            end
          for (forvar159 = (1'h0); (forvar159 < (2'h3)); forvar159 = (forvar159 + (1'h1)))
            begin
              for (forvar160 = (1'h0); (forvar160 < (1'h0)); forvar160 = (forvar160 + (1'h1)))
                begin
                  if ($signed((|(forvar141[(4'h9):(1'h0)] ~^ (~^(8'ha7))))))
                    begin
                      reg161 <= {reg63[(1'h1):(1'h1)]};
                      reg162 <= (~|reg65);
                    end
                  else
                    begin
                      reg161 <= $signed(reg164);
                    end
                  for (forvar163 = (1'h0); (forvar163 < (1'h1)); forvar163 = (forvar163 + (1'h1)))
                    begin
                      reg164 <= forvar170[(5'h10):(2'h2)];
                    end
                end
              for (forvar165 = (1'h0); (forvar165 < (1'h0)); forvar165 = (forvar165 + (1'h1)))
                begin
                  for (forvar166 = (1'h0); (forvar166 < (1'h0)); forvar166 = (forvar166 + (1'h1)))
                    begin
                      reg167 <= (reg148 - $unsigned($signed((8'hb9))));
                      reg168 <= {$unsigned(reg126)};
                      reg169 <= $signed(((~reg174) ?
                          (~^$unsigned((8'hb4))) : (reg230[(2'h3):(2'h2)] << (reg195 < (8'haf)))));
                      reg170 <= {(wire0[(3'h7):(1'h1)] ?
                              (forvar135 <<< (reg186 ?
                                  (8'h9f) : (8'hb6))) : ((reg114 <= reg8) ?
                                  {reg69} : reg189))};
                    end
                  for (forvar171 = (1'h0); (forvar171 < (2'h2)); forvar171 = (forvar171 + (1'h1)))
                    begin
                      reg172 <= reg151;
                      reg173 <= ({((!(8'hb3)) || (!reg76))} ?
                          $signed($signed((^~reg111))) : ($signed($signed(reg50)) ?
                              $signed(reg183) : ((reg109 <= (8'h9c)) ?
                                  reg35[(3'h7):(3'h7)] : (-(8'hac)))));
                      reg174 <= reg37[(3'h4):(2'h2)];
                    end
                end
            end
          for (forvar175 = (1'h0); (forvar175 < (1'h0)); forvar175 = (forvar175 + (1'h1)))
            begin
              for (forvar176 = (1'h0); (forvar176 < (2'h3)); forvar176 = (forvar176 + (1'h1)))
                begin
                  for (forvar177 = (1'h0); (forvar177 < (1'h0)); forvar177 = (forvar177 + (1'h1)))
                    begin
                      reg178 <= reg68[(3'h5):(3'h5)];
                      reg179 <= (8'had);
                      reg180 <= $unsigned(reg157[(1'h1):(1'h1)]);
                    end
                  for (forvar181 = (1'h0); (forvar181 < (1'h1)); forvar181 = (forvar181 + (1'h1)))
                    begin
                      reg182 <= reg31[(1'h1):(1'h1)];
                      reg183 <= (($unsigned((!reg109)) ^ ({reg209} ?
                          {forvar169} : (reg110 ?
                              reg90 : forvar160))) >= {{(~reg26)}});
                      reg184 <= $signed(reg29[(3'h4):(1'h1)]);
                      reg185 <= (~&((reg201[(2'h2):(1'h0)] ?
                          reg65[(3'h6):(3'h6)] : (reg61 > reg93)) <<< (^(reg162 ?
                          reg183 : reg230))));
                    end
                end
              for (forvar186 = (1'h0); (forvar186 < (2'h2)); forvar186 = (forvar186 + (1'h1)))
                begin
                  for (forvar187 = (1'h0); (forvar187 < (1'h1)); forvar187 = (forvar187 + (1'h1)))
                    begin
                      reg188 <= forvar207;
                      reg189 <= reg229[(1'h1):(1'h1)];
                      reg190 <= ($unsigned($signed($signed(forvar155))) ^ reg210[(4'h8):(4'h8)]);
                    end
                  for (forvar191 = (1'h0); (forvar191 < (1'h0)); forvar191 = (forvar191 + (1'h1)))
                    begin
                      reg192 <= (reg85 ? (!(^{reg167})) : {reg164});
                    end
                  reg193 <= (reg138 <= (((reg68 >= forvar181) ?
                      reg10[(4'hd):(3'h4)] : $signed(reg182)) - ({reg50} != $signed((8'hb3)))));
                end
            end
        end
    end
  assign wire233 = reg44[(4'h8):(1'h1)];
  assign wire234 = ($signed(reg181[(2'h2):(2'h2)]) >>> ($unsigned(((8'had) <<< reg124)) != reg162));
  assign wire235 = $signed((($unsigned(reg104) ^ reg179[(4'h8):(2'h2)]) ?
                       (reg86[(2'h3):(2'h3)] ?
                           reg92[(3'h6):(2'h2)] : $unsigned(reg37)) : (reg96[(2'h2):(1'h0)] ^ reg29[(3'h4):(3'h4)])));
  assign wire236 = {((reg215[(1'h1):(1'h1)] * $unsigned(reg175)) ~^ ((reg135 ?
                               reg210 : reg136) ?
                           reg13 : $unsigned(reg67)))};
endmodule