(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param4724 = (~|(^~((!(8'had)) ? (~|(8'hb9)) : ((8'hae) ? (8'hb7) : (8'h9d))))))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h10c4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire3;
  input wire signed [(4'hc):(1'h0)] wire2;
  input wire signed [(5'h10):(1'h0)] wire1;
  input wire [(5'h10):(1'h0)] wire0;
  wire [(2'h2):(1'h0)] wire4661;
  wire [(3'h7):(1'h0)] wire4660;
  wire signed [(3'h7):(1'h0)] wire4518;
  wire [(4'hb):(1'h0)] wire4320;
  wire [(4'he):(1'h0)] wire4319;
  wire [(4'hd):(1'h0)] wire4318;
  wire [(4'hd):(1'h0)] wire4316;
  reg signed [(3'h6):(1'h0)] reg4723 = (1'h0);
  reg [(4'he):(1'h0)] reg4722 = (1'h0);
  reg [(4'hb):(1'h0)] reg4721 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4719 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4718 = (1'h0);
  reg [(3'h5):(1'h0)] reg4717 = (1'h0);
  reg [(4'hb):(1'h0)] reg4715 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4714 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4713 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4711 = (1'h0);
  reg [(5'h10):(1'h0)] reg4710 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4709 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4707 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4706 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4702 = (1'h0);
  reg [(3'h6):(1'h0)] reg4701 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4700 = (1'h0);
  reg [(3'h4):(1'h0)] reg4698 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4696 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4695 = (1'h0);
  reg [(4'h9):(1'h0)] reg4694 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4693 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4692 = (1'h0);
  reg [(4'ha):(1'h0)] reg4688 = (1'h0);
  reg [(4'h9):(1'h0)] reg4675 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4680 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4691 = (1'h0);
  reg [(3'h4):(1'h0)] reg4690 = (1'h0);
  reg [(4'ha):(1'h0)] reg4689 = (1'h0);
  reg [(2'h2):(1'h0)] reg4687 = (1'h0);
  reg [(4'h8):(1'h0)] reg4686 = (1'h0);
  reg [(2'h2):(1'h0)] reg4685 = (1'h0);
  reg [(5'h10):(1'h0)] reg4684 = (1'h0);
  reg [(4'he):(1'h0)] reg4683 = (1'h0);
  reg [(2'h3):(1'h0)] reg4682 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4681 = (1'h0);
  reg [(4'h9):(1'h0)] reg4679 = (1'h0);
  reg [(4'h8):(1'h0)] reg4678 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4676 = (1'h0);
  reg [(4'hb):(1'h0)] reg4671 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4670 = (1'h0);
  reg [(4'h9):(1'h0)] reg4663 = (1'h0);
  reg [(3'h7):(1'h0)] reg4662 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4677 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4674 = (1'h0);
  reg [(4'hc):(1'h0)] reg4673 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4672 = (1'h0);
  reg [(3'h6):(1'h0)] reg4669 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4668 = (1'h0);
  reg [(2'h2):(1'h0)] reg4667 = (1'h0);
  reg [(4'ha):(1'h0)] reg4666 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4665 = (1'h0);
  reg [(2'h2):(1'h0)] reg4664 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4659 = (1'h0);
  reg [(4'hb):(1'h0)] reg4657 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4656 = (1'h0);
  reg [(2'h2):(1'h0)] reg4655 = (1'h0);
  reg [(4'hd):(1'h0)] reg4654 = (1'h0);
  reg [(3'h4):(1'h0)] reg4652 = (1'h0);
  reg [(5'h10):(1'h0)] reg4651 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4650 = (1'h0);
  reg [(4'h9):(1'h0)] reg4649 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4648 = (1'h0);
  reg [(5'h10):(1'h0)] reg4647 = (1'h0);
  reg [(4'hb):(1'h0)] reg4645 = (1'h0);
  reg [(4'ha):(1'h0)] reg4644 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4643 = (1'h0);
  reg [(4'h8):(1'h0)] reg4640 = (1'h0);
  reg [(2'h2):(1'h0)] reg4638 = (1'h0);
  reg [(4'hc):(1'h0)] reg4637 = (1'h0);
  reg [(4'he):(1'h0)] reg4635 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4634 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4633 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4631 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4626 = (1'h0);
  reg [(2'h2):(1'h0)] reg4623 = (1'h0);
  reg [(4'he):(1'h0)] reg4630 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4629 = (1'h0);
  reg [(3'h5):(1'h0)] reg4628 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4627 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4625 = (1'h0);
  reg [(4'he):(1'h0)] reg4624 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4622 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4621 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4620 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4613 = (1'h0);
  reg [(5'h10):(1'h0)] reg4608 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4605 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4597 = (1'h0);
  reg [(3'h6):(1'h0)] reg4618 = (1'h0);
  reg [(4'hc):(1'h0)] reg4616 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4615 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4614 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4612 = (1'h0);
  reg [(5'h10):(1'h0)] reg4611 = (1'h0);
  reg [(4'hc):(1'h0)] reg4610 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4603 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4601 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4607 = (1'h0);
  reg [(4'hd):(1'h0)] reg4606 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4604 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4602 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4600 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4599 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4598 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4585 = (1'h0);
  reg [(3'h6):(1'h0)] reg4596 = (1'h0);
  reg [(4'h9):(1'h0)] reg4595 = (1'h0);
  reg [(2'h2):(1'h0)] reg4594 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4593 = (1'h0);
  reg [(2'h3):(1'h0)] reg4592 = (1'h0);
  reg [(3'h5):(1'h0)] reg4591 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4590 = (1'h0);
  reg [(3'h4):(1'h0)] reg4589 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4588 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4587 = (1'h0);
  reg [(2'h2):(1'h0)] reg4586 = (1'h0);
  reg [(5'h10):(1'h0)] reg4583 = (1'h0);
  reg [(4'hd):(1'h0)] reg4581 = (1'h0);
  reg [(3'h6):(1'h0)] reg4575 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4570 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4563 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4580 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4579 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4578 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4577 = (1'h0);
  reg [(3'h4):(1'h0)] reg4576 = (1'h0);
  reg [(3'h5):(1'h0)] reg4574 = (1'h0);
  reg [(4'hb):(1'h0)] reg4573 = (1'h0);
  reg [(3'h5):(1'h0)] reg4572 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4571 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4569 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4568 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4567 = (1'h0);
  reg [(2'h2):(1'h0)] reg4566 = (1'h0);
  reg [(3'h6):(1'h0)] reg4565 = (1'h0);
  reg [(3'h6):(1'h0)] reg4564 = (1'h0);
  reg [(3'h7):(1'h0)] reg4562 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4561 = (1'h0);
  reg [(4'hd):(1'h0)] reg4560 = (1'h0);
  reg [(5'h10):(1'h0)] reg4559 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4558 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4557 = (1'h0);
  reg [(4'h8):(1'h0)] reg4554 = (1'h0);
  reg [(5'h10):(1'h0)] reg4551 = (1'h0);
  reg [(2'h3):(1'h0)] reg4553 = (1'h0);
  reg [(3'h4):(1'h0)] reg4552 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4545 = (1'h0);
  reg [(3'h5):(1'h0)] reg4549 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4548 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4547 = (1'h0);
  reg [(4'h8):(1'h0)] reg4546 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4544 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4543 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4539 = (1'h0);
  reg [(3'h4):(1'h0)] reg4534 = (1'h0);
  reg [(3'h5):(1'h0)] reg4532 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4542 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4541 = (1'h0);
  reg [(4'hb):(1'h0)] reg4540 = (1'h0);
  reg [(4'hd):(1'h0)] reg4538 = (1'h0);
  reg [(4'hf):(1'h0)] reg4537 = (1'h0);
  reg [(4'hc):(1'h0)] reg4536 = (1'h0);
  reg [(3'h7):(1'h0)] reg4535 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4533 = (1'h0);
  reg [(4'hb):(1'h0)] reg4531 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4530 = (1'h0);
  reg [(4'hf):(1'h0)] reg4529 = (1'h0);
  reg [(2'h2):(1'h0)] reg4528 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4521 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4527 = (1'h0);
  reg [(2'h3):(1'h0)] reg4525 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4524 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4523 = (1'h0);
  reg [(3'h4):(1'h0)] reg4522 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4495 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4517 = (1'h0);
  reg [(4'h8):(1'h0)] reg4516 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4515 = (1'h0);
  reg [(3'h4):(1'h0)] reg4514 = (1'h0);
  reg [(4'he):(1'h0)] reg4513 = (1'h0);
  reg [(2'h3):(1'h0)] reg4512 = (1'h0);
  reg [(4'hb):(1'h0)] reg4511 = (1'h0);
  reg [(3'h6):(1'h0)] reg4510 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4509 = (1'h0);
  reg [(4'hb):(1'h0)] reg4507 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4506 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4505 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4504 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4502 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4501 = (1'h0);
  reg [(3'h4):(1'h0)] reg4500 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4499 = (1'h0);
  reg [(2'h3):(1'h0)] reg4497 = (1'h0);
  reg [(4'h9):(1'h0)] reg4496 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4494 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4493 = (1'h0);
  reg [(4'h8):(1'h0)] reg4492 = (1'h0);
  reg [(4'he):(1'h0)] reg4491 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4489 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4487 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4486 = (1'h0);
  reg [(4'hf):(1'h0)] reg4485 = (1'h0);
  reg [(2'h3):(1'h0)] reg4484 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4467 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4465 = (1'h0);
  reg [(4'hc):(1'h0)] reg4483 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4476 = (1'h0);
  reg [(3'h4):(1'h0)] reg4482 = (1'h0);
  reg [(4'h9):(1'h0)] reg4481 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4480 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4479 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4478 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4477 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4472 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4475 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4474 = (1'h0);
  reg [(3'h6):(1'h0)] reg4473 = (1'h0);
  reg [(2'h2):(1'h0)] reg4471 = (1'h0);
  reg [(4'he):(1'h0)] reg4469 = (1'h0);
  reg [(2'h2):(1'h0)] reg4468 = (1'h0);
  reg [(4'hc):(1'h0)] reg4466 = (1'h0);
  reg [(2'h3):(1'h0)] reg4464 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4463 = (1'h0);
  reg [(3'h6):(1'h0)] reg4462 = (1'h0);
  reg [(4'hc):(1'h0)] reg4461 = (1'h0);
  reg [(4'h9):(1'h0)] reg4460 = (1'h0);
  reg [(4'he):(1'h0)] reg4457 = (1'h0);
  reg [(4'ha):(1'h0)] reg4456 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4455 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4453 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4452 = (1'h0);
  reg [(5'h10):(1'h0)] reg4451 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4450 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4449 = (1'h0);
  reg [(4'h8):(1'h0)] reg4447 = (1'h0);
  reg [(3'h7):(1'h0)] reg4446 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4445 = (1'h0);
  reg [(4'h9):(1'h0)] reg4444 = (1'h0);
  reg [(3'h4):(1'h0)] reg4441 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4440 = (1'h0);
  reg [(4'hc):(1'h0)] reg4439 = (1'h0);
  reg [(3'h4):(1'h0)] reg4437 = (1'h0);
  reg [(4'h8):(1'h0)] reg4436 = (1'h0);
  reg [(3'h6):(1'h0)] reg4435 = (1'h0);
  reg [(3'h4):(1'h0)] reg4434 = (1'h0);
  reg [(4'h8):(1'h0)] reg4433 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4432 = (1'h0);
  reg [(4'hd):(1'h0)] reg4431 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4430 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4427 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4426 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4424 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4423 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4422 = (1'h0);
  reg [(4'ha):(1'h0)] reg4421 = (1'h0);
  reg [(4'h8):(1'h0)] reg4419 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4418 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4415 = (1'h0);
  reg [(3'h7):(1'h0)] reg4414 = (1'h0);
  reg [(5'h10):(1'h0)] reg4413 = (1'h0);
  reg [(4'hb):(1'h0)] reg4412 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4411 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4405 = (1'h0);
  reg [(4'h8):(1'h0)] reg4409 = (1'h0);
  reg [(3'h5):(1'h0)] reg4408 = (1'h0);
  reg [(4'he):(1'h0)] reg4407 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4406 = (1'h0);
  reg [(3'h6):(1'h0)] reg4404 = (1'h0);
  reg [(4'ha):(1'h0)] reg4380 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4375 = (1'h0);
  reg [(4'h9):(1'h0)] reg4376 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4401 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4400 = (1'h0);
  reg [(4'hf):(1'h0)] reg4399 = (1'h0);
  reg [(4'hb):(1'h0)] reg4398 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4397 = (1'h0);
  reg [(2'h3):(1'h0)] reg4395 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4394 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4393 = (1'h0);
  reg [(4'hd):(1'h0)] reg4391 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4390 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4389 = (1'h0);
  reg [(4'hc):(1'h0)] reg4388 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4387 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4386 = (1'h0);
  reg [(3'h4):(1'h0)] reg4385 = (1'h0);
  reg [(2'h3):(1'h0)] reg4384 = (1'h0);
  reg [(2'h3):(1'h0)] reg4383 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4382 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4381 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4379 = (1'h0);
  reg [(3'h6):(1'h0)] reg4378 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4377 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4373 = (1'h0);
  reg [(3'h5):(1'h0)] reg4372 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4371 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4366 = (1'h0);
  reg [(4'h8):(1'h0)] reg4370 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4369 = (1'h0);
  reg [(2'h3):(1'h0)] reg4368 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4367 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4365 = (1'h0);
  reg [(4'ha):(1'h0)] reg4364 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4363 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4362 = (1'h0);
  reg [(3'h6):(1'h0)] reg4360 = (1'h0);
  reg [(3'h5):(1'h0)] reg4359 = (1'h0);
  reg [(2'h3):(1'h0)] reg4358 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4357 = (1'h0);
  reg [(4'ha):(1'h0)] reg4356 = (1'h0);
  reg [(4'he):(1'h0)] reg4355 = (1'h0);
  reg [(3'h6):(1'h0)] reg4354 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4353 = (1'h0);
  reg [(2'h2):(1'h0)] reg4352 = (1'h0);
  reg [(4'h9):(1'h0)] reg4348 = (1'h0);
  reg [(4'hc):(1'h0)] reg4344 = (1'h0);
  reg [(4'hf):(1'h0)] reg4343 = (1'h0);
  reg [(3'h5):(1'h0)] reg4351 = (1'h0);
  reg [(4'he):(1'h0)] reg4350 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4349 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4347 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4346 = (1'h0);
  reg [(5'h10):(1'h0)] reg4345 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4339 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4337 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4342 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4341 = (1'h0);
  reg [(4'h8):(1'h0)] reg4340 = (1'h0);
  reg [(4'ha):(1'h0)] reg4338 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4336 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4335 = (1'h0);
  reg [(5'h10):(1'h0)] reg4334 = (1'h0);
  reg [(2'h3):(1'h0)] reg4333 = (1'h0);
  reg [(3'h7):(1'h0)] reg4332 = (1'h0);
  reg [(4'hc):(1'h0)] reg4331 = (1'h0);
  reg [(4'hd):(1'h0)] reg4330 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4328 = (1'h0);
  reg [(2'h3):(1'h0)] reg4327 = (1'h0);
  reg [(3'h6):(1'h0)] reg4324 = (1'h0);
  reg [(3'h5):(1'h0)] reg4322 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4720 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4716 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4712 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4708 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4705 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4704 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4703 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4699 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4697 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4690 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4679 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4686 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4683 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4672 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4688 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4680 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4673 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4664 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4676 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4675 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4671 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4670 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4663 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4662 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4658 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4653 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4646 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4642 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4641 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4639 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4621 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4636 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4632 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4630 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4625 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4620 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4626 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4623 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4619 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4604 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4599 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4617 = (1'h0);
  reg [(4'he):(1'h0)] forvar4613 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4609 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4608 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4605 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4603 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4601 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4597 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4589 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4585 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4584 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4582 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4573 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4572 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4567 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4564 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4561 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4560 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4554 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4575 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4570 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4563 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4556 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4555 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4551 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4550 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4547 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4544 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4545 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4537 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4529 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4539 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4534 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4532 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4528 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4526 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4521 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4520 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4519 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4508 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4503 = (1'h0);
  reg [(4'he):(1'h0)] forvar4498 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4495 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4490 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4488 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4484 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4479 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4478 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4474 = (1'h0);
  reg [(4'he):(1'h0)] forvar4473 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4464 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4462 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4476 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4472 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4470 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4467 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4465 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4461 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4459 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4458 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4454 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4448 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4443 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4442 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4438 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4429 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4428 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4425 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4420 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4417 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4416 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4411 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4410 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4405 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4403 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4402 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4383 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4396 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4392 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4380 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4376 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4375 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4374 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4363 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4366 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4361 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4347 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4346 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4348 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4344 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4343 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4334 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4339 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4337 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4329 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4326 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4325 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4323 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4321 = (1'h0);
  assign y = {wire4661,
                 wire4660,
                 wire4518,
                 wire4320,
                 wire4319,
                 wire4318,
                 wire4316,
                 reg4723,
                 reg4722,
                 reg4721,
                 reg4719,
                 reg4718,
                 reg4717,
                 reg4715,
                 reg4714,
                 reg4713,
                 reg4711,
                 reg4710,
                 reg4709,
                 reg4707,
                 reg4706,
                 reg4702,
                 reg4701,
                 reg4700,
                 reg4698,
                 reg4696,
                 reg4695,
                 reg4694,
                 reg4693,
                 reg4692,
                 reg4688,
                 reg4675,
                 reg4680,
                 reg4691,
                 reg4690,
                 reg4689,
                 reg4687,
                 reg4686,
                 reg4685,
                 reg4684,
                 reg4683,
                 reg4682,
                 reg4681,
                 reg4679,
                 reg4678,
                 reg4676,
                 reg4671,
                 reg4670,
                 reg4663,
                 reg4662,
                 reg4677,
                 reg4674,
                 reg4673,
                 reg4672,
                 reg4669,
                 reg4668,
                 reg4667,
                 reg4666,
                 reg4665,
                 reg4664,
                 reg4659,
                 reg4657,
                 reg4656,
                 reg4655,
                 reg4654,
                 reg4652,
                 reg4651,
                 reg4650,
                 reg4649,
                 reg4648,
                 reg4647,
                 reg4645,
                 reg4644,
                 reg4643,
                 reg4640,
                 reg4638,
                 reg4637,
                 reg4635,
                 reg4634,
                 reg4633,
                 reg4631,
                 reg4626,
                 reg4623,
                 reg4630,
                 reg4629,
                 reg4628,
                 reg4627,
                 reg4625,
                 reg4624,
                 reg4622,
                 reg4621,
                 reg4620,
                 reg4613,
                 reg4608,
                 reg4605,
                 reg4597,
                 reg4618,
                 reg4616,
                 reg4615,
                 reg4614,
                 reg4612,
                 reg4611,
                 reg4610,
                 reg4603,
                 reg4601,
                 reg4607,
                 reg4606,
                 reg4604,
                 reg4602,
                 reg4600,
                 reg4599,
                 reg4598,
                 reg4585,
                 reg4596,
                 reg4595,
                 reg4594,
                 reg4593,
                 reg4592,
                 reg4591,
                 reg4590,
                 reg4589,
                 reg4588,
                 reg4587,
                 reg4586,
                 reg4583,
                 reg4581,
                 reg4575,
                 reg4570,
                 reg4563,
                 reg4580,
                 reg4579,
                 reg4578,
                 reg4577,
                 reg4576,
                 reg4574,
                 reg4573,
                 reg4572,
                 reg4571,
                 reg4569,
                 reg4568,
                 reg4567,
                 reg4566,
                 reg4565,
                 reg4564,
                 reg4562,
                 reg4561,
                 reg4560,
                 reg4559,
                 reg4558,
                 reg4557,
                 reg4554,
                 reg4551,
                 reg4553,
                 reg4552,
                 reg4545,
                 reg4549,
                 reg4548,
                 reg4547,
                 reg4546,
                 reg4544,
                 reg4543,
                 reg4539,
                 reg4534,
                 reg4532,
                 reg4542,
                 reg4541,
                 reg4540,
                 reg4538,
                 reg4537,
                 reg4536,
                 reg4535,
                 reg4533,
                 reg4531,
                 reg4530,
                 reg4529,
                 reg4528,
                 reg4521,
                 reg4527,
                 reg4525,
                 reg4524,
                 reg4523,
                 reg4522,
                 reg4495,
                 reg4517,
                 reg4516,
                 reg4515,
                 reg4514,
                 reg4513,
                 reg4512,
                 reg4511,
                 reg4510,
                 reg4509,
                 reg4507,
                 reg4506,
                 reg4505,
                 reg4504,
                 reg4502,
                 reg4501,
                 reg4500,
                 reg4499,
                 reg4497,
                 reg4496,
                 reg4494,
                 reg4493,
                 reg4492,
                 reg4491,
                 reg4489,
                 reg4487,
                 reg4486,
                 reg4485,
                 reg4484,
                 reg4467,
                 reg4465,
                 reg4483,
                 reg4476,
                 reg4482,
                 reg4481,
                 reg4480,
                 reg4479,
                 reg4478,
                 reg4477,
                 reg4472,
                 reg4475,
                 reg4474,
                 reg4473,
                 reg4471,
                 reg4469,
                 reg4468,
                 reg4466,
                 reg4464,
                 reg4463,
                 reg4462,
                 reg4461,
                 reg4460,
                 reg4457,
                 reg4456,
                 reg4455,
                 reg4453,
                 reg4452,
                 reg4451,
                 reg4450,
                 reg4449,
                 reg4447,
                 reg4446,
                 reg4445,
                 reg4444,
                 reg4441,
                 reg4440,
                 reg4439,
                 reg4437,
                 reg4436,
                 reg4435,
                 reg4434,
                 reg4433,
                 reg4432,
                 reg4431,
                 reg4430,
                 reg4427,
                 reg4426,
                 reg4424,
                 reg4423,
                 reg4422,
                 reg4421,
                 reg4419,
                 reg4418,
                 reg4415,
                 reg4414,
                 reg4413,
                 reg4412,
                 reg4411,
                 reg4405,
                 reg4409,
                 reg4408,
                 reg4407,
                 reg4406,
                 reg4404,
                 reg4380,
                 reg4375,
                 reg4376,
                 reg4401,
                 reg4400,
                 reg4399,
                 reg4398,
                 reg4397,
                 reg4395,
                 reg4394,
                 reg4393,
                 reg4391,
                 reg4390,
                 reg4389,
                 reg4388,
                 reg4387,
                 reg4386,
                 reg4385,
                 reg4384,
                 reg4383,
                 reg4382,
                 reg4381,
                 reg4379,
                 reg4378,
                 reg4377,
                 reg4373,
                 reg4372,
                 reg4371,
                 reg4366,
                 reg4370,
                 reg4369,
                 reg4368,
                 reg4367,
                 reg4365,
                 reg4364,
                 reg4363,
                 reg4362,
                 reg4360,
                 reg4359,
                 reg4358,
                 reg4357,
                 reg4356,
                 reg4355,
                 reg4354,
                 reg4353,
                 reg4352,
                 reg4348,
                 reg4344,
                 reg4343,
                 reg4351,
                 reg4350,
                 reg4349,
                 reg4347,
                 reg4346,
                 reg4345,
                 reg4339,
                 reg4337,
                 reg4342,
                 reg4341,
                 reg4340,
                 reg4338,
                 reg4336,
                 reg4335,
                 reg4334,
                 reg4333,
                 reg4332,
                 reg4331,
                 reg4330,
                 reg4328,
                 reg4327,
                 reg4324,
                 reg4322,
                 forvar4720,
                 forvar4716,
                 forvar4712,
                 forvar4708,
                 forvar4705,
                 forvar4704,
                 forvar4703,
                 forvar4699,
                 forvar4697,
                 forvar4690,
                 forvar4679,
                 forvar4686,
                 forvar4683,
                 forvar4672,
                 forvar4688,
                 forvar4680,
                 forvar4673,
                 forvar4664,
                 forvar4676,
                 forvar4675,
                 forvar4671,
                 forvar4670,
                 forvar4663,
                 forvar4662,
                 forvar4658,
                 forvar4653,
                 forvar4646,
                 forvar4642,
                 forvar4641,
                 forvar4639,
                 forvar4621,
                 forvar4636,
                 forvar4632,
                 forvar4630,
                 forvar4625,
                 forvar4620,
                 forvar4626,
                 forvar4623,
                 forvar4619,
                 forvar4604,
                 forvar4599,
                 forvar4617,
                 forvar4613,
                 forvar4609,
                 forvar4608,
                 forvar4605,
                 forvar4603,
                 forvar4601,
                 forvar4597,
                 forvar4589,
                 forvar4585,
                 forvar4584,
                 forvar4582,
                 forvar4573,
                 forvar4572,
                 forvar4567,
                 forvar4564,
                 forvar4561,
                 forvar4560,
                 forvar4554,
                 forvar4575,
                 forvar4570,
                 forvar4563,
                 forvar4556,
                 forvar4555,
                 forvar4551,
                 forvar4550,
                 forvar4547,
                 forvar4544,
                 forvar4545,
                 forvar4537,
                 forvar4529,
                 forvar4539,
                 forvar4534,
                 forvar4532,
                 forvar4528,
                 forvar4526,
                 forvar4521,
                 forvar4520,
                 forvar4519,
                 forvar4508,
                 forvar4503,
                 forvar4498,
                 forvar4495,
                 forvar4490,
                 forvar4488,
                 forvar4484,
                 forvar4479,
                 forvar4478,
                 forvar4474,
                 forvar4473,
                 forvar4464,
                 forvar4462,
                 forvar4476,
                 forvar4472,
                 forvar4470,
                 forvar4467,
                 forvar4465,
                 forvar4461,
                 forvar4459,
                 forvar4458,
                 forvar4454,
                 forvar4448,
                 forvar4443,
                 forvar4442,
                 forvar4438,
                 forvar4429,
                 forvar4428,
                 forvar4425,
                 forvar4420,
                 forvar4417,
                 forvar4416,
                 forvar4411,
                 forvar4410,
                 forvar4405,
                 forvar4403,
                 forvar4402,
                 forvar4383,
                 forvar4396,
                 forvar4392,
                 forvar4380,
                 forvar4376,
                 forvar4375,
                 forvar4374,
                 forvar4363,
                 forvar4366,
                 forvar4361,
                 forvar4347,
                 forvar4346,
                 forvar4348,
                 forvar4344,
                 forvar4343,
                 forvar4334,
                 forvar4339,
                 forvar4337,
                 forvar4329,
                 forvar4326,
                 forvar4325,
                 forvar4323,
                 forvar4321,
                 (1'h0)};
  module4 #() modinst4317 (.wire5(wire0), .clk(clk), .wire6(wire1), .wire7(wire3), .y(wire4316), .wire8(wire2));
  assign wire4318 = wire0[(4'hd):(4'h9)];
  assign wire4319 = (|(|(~^wire0[(3'h5):(2'h3)])));
  assign wire4320 = ((wire0 == ($signed(wire4316) >= (wire4316 | wire4316))) < (wire4318[(1'h1):(1'h0)] >> (wire3 - $unsigned(wire4318))));
  always
    @(posedge clk) begin
      for (forvar4321 = (1'h0); (forvar4321 < (2'h3)); forvar4321 = (forvar4321 + (1'h1)))
        begin
          reg4322 <= $unsigned(wire4316[(4'hc):(4'h8)]);
          for (forvar4323 = (1'h0); (forvar4323 < (1'h1)); forvar4323 = (forvar4323 + (1'h1)))
            begin
              reg4324 <= (($unsigned((wire4320 ?
                  forvar4321 : (8'hb3))) + wire1) ~^ (wire4320[(3'h7):(3'h5)] ?
                  forvar4321[(4'hd):(4'ha)] : wire0));
              for (forvar4325 = (1'h0); (forvar4325 < (2'h2)); forvar4325 = (forvar4325 + (1'h1)))
                begin
                  for (forvar4326 = (1'h0); (forvar4326 < (2'h3)); forvar4326 = (forvar4326 + (1'h1)))
                    begin
                      reg4327 <= reg4322[(2'h2):(2'h2)];
                      reg4328 <= $signed($unsigned(forvar4321));
                    end
                  for (forvar4329 = (1'h0); (forvar4329 < (2'h3)); forvar4329 = (forvar4329 + (1'h1)))
                    begin
                      reg4330 <= ((($unsigned(reg4327) <= wire0[(3'h5):(2'h3)]) ?
                              (wire4319[(3'h5):(3'h4)] ?
                                  forvar4323 : (~|wire0)) : wire2[(2'h2):(1'h0)]) ?
                          (($signed((8'hb7)) ? reg4322 : wire3) ?
                              $signed((^~wire1)) : forvar4329) : {{{forvar4329}}});
                      reg4331 <= {{(wire1[(5'h10):(1'h1)] ?
                                  wire4318 : (~reg4322))}};
                      reg4332 <= wire4320;
                      reg4333 <= (reg4327 ~^ ((wire4319 ?
                              $unsigned(wire4320) : wire4318[(3'h6):(2'h2)]) ?
                          ($unsigned(wire4320) ?
                              (~&reg4322) : $signed((8'ha7))) : $signed((~^reg4330))));
                    end
                end
              if ((wire4320[(3'h7):(3'h7)] ?
                  (($signed(reg4332) * $unsigned(wire2)) || (+(~|(8'ha1)))) : (!((reg4333 ^ wire4316) * (~(8'ha0))))))
                begin
                  if ($unsigned(reg4328))
                    begin
                      reg4334 <= (forvar4325[(4'ha):(1'h0)] ?
                          (~&forvar4329[(4'ha):(3'h4)]) : $unsigned(reg4322));
                    end
                  else
                    begin
                      reg4334 <= (((wire4318[(4'hb):(4'ha)] ?
                              {forvar4321} : {wire2}) ?
                          ((wire1 ? forvar4325 : wire0) ?
                              $signed(forvar4325) : $signed(wire2)) : $signed(forvar4326)) & $unsigned(($unsigned(forvar4323) << $signed(reg4330))));
                      reg4335 <= (~^($signed(reg4328[(2'h2):(2'h2)]) ?
                          ((reg4334 > wire0) == $unsigned(reg4332)) : forvar4323[(3'h6):(2'h3)]));
                      reg4336 <= wire0;
                    end
                  for (forvar4337 = (1'h0); (forvar4337 < (2'h2)); forvar4337 = (forvar4337 + (1'h1)))
                    begin
                      reg4338 <= $signed(($unsigned($unsigned(wire4319)) < (reg4327[(2'h3):(2'h2)] == forvar4329)));
                    end
                  for (forvar4339 = (1'h0); (forvar4339 < (2'h2)); forvar4339 = (forvar4339 + (1'h1)))
                    begin
                      reg4340 <= $unsigned((|$unsigned((reg4334 ?
                          (8'had) : wire0))));
                      reg4341 <= $signed({reg4332[(3'h7):(2'h3)]});
                      reg4342 <= (($signed($unsigned(forvar4339)) <= wire4318) ?
                          (reg4332[(2'h3):(2'h3)] | $signed($signed(reg4328))) : ($unsigned((reg4341 == (8'ha9))) == (8'hba)));
                    end
                end
              else
                begin
                  for (forvar4334 = (1'h0); (forvar4334 < (2'h3)); forvar4334 = (forvar4334 + (1'h1)))
                    begin
                      reg4335 <= ($unsigned(((wire2 ?
                              wire0 : (8'hb3)) ~^ (reg4331 ?
                              reg4324 : wire4318))) ?
                          (((reg4336 >> reg4330) ?
                              reg4335 : $signed(wire3)) >= $unsigned(reg4324[(3'h4):(1'h0)])) : (reg4334 ?
                              reg4342 : ((forvar4334 ^ reg4327) ?
                                  $unsigned(wire1) : (wire4318 == wire1))));
                    end
                  if (forvar4337)
                    begin
                      reg4336 <= wire4318[(4'h8):(3'h5)];
                      reg4337 <= $signed(($signed((reg4342 != reg4338)) ^ $signed($signed(wire4320))));
                      reg4338 <= $unsigned($signed(wire4319[(4'hc):(3'h6)]));
                    end
                  else
                    begin
                      reg4336 <= $unsigned(reg4322[(1'h1):(1'h0)]);
                      reg4337 <= reg4341[(3'h4):(1'h1)];
                    end
                  if ($unsigned((reg4333 || reg4327[(2'h3):(2'h2)])))
                    begin
                      reg4339 <= wire3;
                      reg4340 <= reg4340[(1'h0):(1'h0)];
                      reg4341 <= ((8'had) ?
                          (&{((8'ha3) ?
                                  (8'ha5) : reg4324)}) : $signed(wire4316));
                      reg4342 <= wire3[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg4339 <= $unsigned(reg4322);
                    end
                end
            end
          if ($unsigned((~wire3)))
            begin
              for (forvar4343 = (1'h0); (forvar4343 < (1'h1)); forvar4343 = (forvar4343 + (1'h1)))
                begin
                  for (forvar4344 = (1'h0); (forvar4344 < (2'h3)); forvar4344 = (forvar4344 + (1'h1)))
                    begin
                      reg4345 <= forvar4339;
                      reg4346 <= $unsigned(forvar4339[(3'h7):(2'h3)]);
                      reg4347 <= reg4337[(1'h1):(1'h1)];
                    end
                  for (forvar4348 = (1'h0); (forvar4348 < (1'h0)); forvar4348 = (forvar4348 + (1'h1)))
                    begin
                      reg4349 <= ($signed(wire4320) ~^ reg4328[(2'h2):(1'h0)]);
                      reg4350 <= wire0;
                      reg4351 <= $signed({forvar4321[(4'h9):(4'h8)]});
                    end
                end
            end
          else
            begin
              if ($signed(reg4339))
                begin
                  reg4343 <= {(((wire4316 ? reg4335 : reg4339) >>> reg4322) ?
                          $signed((forvar4348 << reg4331)) : forvar4329[(1'h1):(1'h0)])};
                  reg4344 <= wire4316[(3'h7):(3'h5)];
                  reg4345 <= reg4346;
                end
              else
                begin
                  reg4343 <= ((^$signed(reg4333[(1'h0):(1'h0)])) & wire4316[(3'h6):(1'h0)]);
                end
              for (forvar4346 = (1'h0); (forvar4346 < (1'h0)); forvar4346 = (forvar4346 + (1'h1)))
                begin
                  for (forvar4347 = (1'h0); (forvar4347 < (2'h3)); forvar4347 = (forvar4347 + (1'h1)))
                    begin
                      reg4348 <= forvar4329[(4'ha):(4'h9)];
                      reg4349 <= (^~$signed($unsigned((~^wire4318))));
                      reg4350 <= (~$unsigned((-$unsigned(forvar4348))));
                      reg4351 <= (8'hab);
                    end
                  if ($unsigned(reg4349[(3'h5):(1'h1)]))
                    begin
                      reg4352 <= $signed(({reg4327[(2'h2):(1'h1)]} != (reg4351 - (reg4327 ?
                          reg4334 : reg4335))));
                    end
                  else
                    begin
                      reg4352 <= ((~|((wire4316 ? reg4330 : reg4337) ?
                          (reg4344 < reg4341) : (8'ha8))) ^ $unsigned(forvar4334));
                      reg4353 <= $unsigned((~&(!$signed(reg4347))));
                      reg4354 <= reg4335;
                      reg4355 <= ({reg4348[(4'h8):(3'h4)]} ?
                          (+forvar4321) : {((^~reg4348) >= forvar4346[(4'hb):(4'ha)])});
                    end
                  if ((reg4341[(3'h5):(3'h4)] ~^ (^($signed(reg4327) <= wire1))))
                    begin
                      reg4356 <= {$signed(((8'had) ?
                              $unsigned(reg4340) : $signed((8'ha1))))};
                      reg4357 <= $unsigned($signed($signed(forvar4329)));
                      reg4358 <= reg4348[(4'h9):(2'h2)];
                      reg4359 <= $signed($unsigned($signed(forvar4346)));
                    end
                  else
                    begin
                      reg4356 <= wire4319;
                      reg4357 <= (~&reg4322);
                      reg4358 <= wire3;
                    end
                end
              if ((-reg4353))
                begin
                  if ($signed(reg4337[(3'h6):(2'h3)]))
                    begin
                      reg4360 <= ({((wire4316 ?
                              reg4354 : reg4344) ^~ {reg4328})} <= forvar4325);
                    end
                  else
                    begin
                      reg4360 <= (~|($signed((wire2 * forvar4347)) ?
                          ($signed(reg4324) ?
                              reg4355 : $signed(reg4351)) : (~^(reg4357 ^ (8'ha1)))));
                    end
                  for (forvar4361 = (1'h0); (forvar4361 < (1'h1)); forvar4361 = (forvar4361 + (1'h1)))
                    begin
                      reg4362 <= reg4322[(2'h2):(1'h1)];
                      reg4363 <= $signed((reg4337 ?
                          $unsigned($unsigned(forvar4348)) : ({(8'ha9)} >= (forvar4325 ^~ (8'h9e)))));
                      reg4364 <= (8'hb8);
                    end
                  reg4365 <= (($unsigned((|reg4333)) && $signed(forvar4346)) ?
                      reg4322 : (8'hb2));
                  for (forvar4366 = (1'h0); (forvar4366 < (2'h3)); forvar4366 = (forvar4366 + (1'h1)))
                    begin
                      reg4367 <= reg4339;
                      reg4368 <= $unsigned(({(^reg4365)} ?
                          ((forvar4321 && reg4331) << reg4337) : $signed(forvar4323[(3'h4):(1'h0)])));
                      reg4369 <= (reg4343 ? wire4316 : reg4342);
                      reg4370 <= ((reg4337[(3'h5):(3'h4)] ?
                              $signed(forvar4325) : (((8'haf) - forvar4361) ?
                                  (8'ha1) : reg4353[(2'h2):(1'h0)])) ?
                          forvar4346 : ($signed((^reg4363)) ?
                              ((&reg4349) ?
                                  (-forvar4325) : forvar4343) : wire4320));
                    end
                end
              else
                begin
                  reg4360 <= $signed((-forvar4366[(4'h8):(2'h2)]));
                  for (forvar4361 = (1'h0); (forvar4361 < (1'h0)); forvar4361 = (forvar4361 + (1'h1)))
                    begin
                      reg4362 <= (forvar4326[(2'h2):(2'h2)] < (|(|(reg4357 ?
                          (8'h9f) : reg4324))));
                    end
                  for (forvar4363 = (1'h0); (forvar4363 < (1'h0)); forvar4363 = (forvar4363 + (1'h1)))
                    begin
                      reg4364 <= ((&(((8'ha6) ?
                              (8'hb2) : forvar4343) >= reg4338)) ?
                          reg4358 : (&reg4339));
                      reg4365 <= ((reg4357[(4'hc):(3'h5)] > reg4362[(2'h3):(1'h1)]) ?
                          ((-reg4332[(3'h5):(2'h2)]) << ({reg4337} ?
                              (forvar4321 ?
                                  reg4364 : reg4346) : wire4316)) : (~|forvar4326));
                      reg4366 <= $signed({($unsigned(reg4359) >> $unsigned(wire2))});
                      reg4367 <= $signed((((reg4351 ?
                          reg4351 : reg4352) << (reg4355 ?
                          reg4345 : reg4343)) ^~ ((reg4347 <<< reg4339) + (~|reg4347))));
                    end
                end
              reg4371 <= ((&$unsigned($signed(reg4349))) << (&(!(forvar4361 ?
                  forvar4337 : reg4345))));
            end
        end
      reg4372 <= $signed((reg4370 ? forvar4346[(4'ha):(2'h2)] : (8'hae)));
      reg4373 <= (((|((8'hba) ?
          forvar4339 : reg4365)) ~^ reg4324) > wire2[(4'h9):(4'h8)]);
    end
  always
    @(posedge clk) begin
      if ({(((-reg4360) ^ reg4350) ?
              ($signed((8'hae)) * (~^reg4346)) : $unsigned((reg4369 <= reg4327)))})
        begin
          for (forvar4374 = (1'h0); (forvar4374 < (1'h0)); forvar4374 = (forvar4374 + (1'h1)))
            begin
              for (forvar4375 = (1'h0); (forvar4375 < (2'h3)); forvar4375 = (forvar4375 + (1'h1)))
                begin
                  for (forvar4376 = (1'h0); (forvar4376 < (2'h3)); forvar4376 = (forvar4376 + (1'h1)))
                    begin
                      reg4377 <= ((|{$signed(forvar4374)}) & ((forvar4375 ?
                              (forvar4374 ? wire4318 : reg4334) : (reg4322 ?
                                  (8'hb0) : reg4359)) ?
                          ((^reg4324) << $unsigned(reg4342)) : reg4371));
                      reg4378 <= (($signed((reg4369 ?
                              reg4336 : reg4341)) ^~ (wire4320[(4'h9):(2'h3)] <<< reg4352[(1'h1):(1'h0)])) ?
                          $unsigned(((reg4337 < reg4341) ?
                              (~^(8'ha7)) : reg4356)) : (8'hb6));
                      reg4379 <= ($unsigned({(~&(8'hab))}) << $unsigned((-$unsigned(reg4373))));
                    end
                  for (forvar4380 = (1'h0); (forvar4380 < (2'h3)); forvar4380 = (forvar4380 + (1'h1)))
                    begin
                      reg4381 <= $unsigned($unsigned($signed((reg4349 || reg4359))));
                      reg4382 <= $signed($signed(((~^wire1) ~^ $signed(reg4381))));
                    end
                  if ({reg4366})
                    begin
                      reg4383 <= forvar4380;
                      reg4384 <= ((~&reg4345[(4'hc):(2'h3)]) >> (reg4369[(3'h5):(3'h4)] ?
                          $unsigned($unsigned((8'h9e))) : (((8'hb2) ?
                                  reg4382 : (8'hb7)) ?
                              (reg4348 ? wire4320 : forvar4376) : reg4332)));
                      reg4385 <= forvar4374;
                    end
                  else
                    begin
                      reg4383 <= reg4338;
                      reg4384 <= forvar4380[(1'h1):(1'h0)];
                      reg4385 <= reg4371[(4'hf):(4'hd)];
                      reg4386 <= reg4354;
                    end
                  if (($unsigned($signed($signed(wire2))) ?
                      ($signed(((8'h9c) && (8'ha2))) < {(forvar4374 ^ (8'h9f))}) : (|((reg4363 <<< reg4330) ?
                          ((8'hb0) > reg4364) : $signed(wire1)))))
                    begin
                      reg4387 <= $unsigned($signed(wire4316));
                      reg4388 <= (~&((reg4381[(4'hd):(3'h7)] >> (~&reg4363)) == $unsigned((reg4322 ?
                          reg4330 : (8'hb3)))));
                      reg4389 <= (reg4382 >>> forvar4380[(1'h0):(1'h0)]);
                      reg4390 <= $unsigned($unsigned({$signed(reg4365)}));
                    end
                  else
                    begin
                      reg4387 <= $unsigned($unsigned(reg4377[(2'h3):(1'h0)]));
                    end
                end
              reg4391 <= $signed(wire0);
              for (forvar4392 = (1'h0); (forvar4392 < (1'h0)); forvar4392 = (forvar4392 + (1'h1)))
                begin
                  if (wire2[(3'h7):(1'h0)])
                    begin
                      reg4393 <= $signed(reg4382[(3'h6):(1'h1)]);
                      reg4394 <= (({forvar4376[(3'h6):(1'h1)]} * $signed((^~reg4332))) ?
                          (($signed(reg4371) ?
                              forvar4376 : (~^reg4331)) <<< ((~(8'ha6)) ?
                              reg4393[(2'h2):(2'h2)] : (&reg4366))) : $signed(wire4319[(4'hd):(2'h3)]));
                      reg4395 <= $unsigned($signed(((reg4349 - wire4318) <<< (reg4335 ^~ reg4358))));
                    end
                  else
                    begin
                      reg4393 <= (({$signed(reg4352)} ?
                              (~|(8'hb9)) : {(reg4369 ? reg4366 : reg4335)}) ?
                          $signed(((~&wire4316) >>> $signed(reg4347))) : wire4316[(3'h7):(3'h5)]);
                    end
                  for (forvar4396 = (1'h0); (forvar4396 < (1'h1)); forvar4396 = (forvar4396 + (1'h1)))
                    begin
                      reg4397 <= reg4360;
                    end
                  reg4398 <= reg4395[(1'h1):(1'h1)];
                  if ($signed({($signed((8'haf)) + $signed((8'hb5)))}))
                    begin
                      reg4399 <= $signed((8'hb8));
                      reg4400 <= $unsigned(wire4318);
                      reg4401 <= ($signed(reg4322[(3'h4):(1'h1)]) && $unsigned(($signed(reg4389) ?
                          $signed(reg4371) : (8'ha7))));
                    end
                  else
                    begin
                      reg4399 <= (|$signed(reg4357));
                    end
                end
            end
        end
      else
        begin
          for (forvar4374 = (1'h0); (forvar4374 < (1'h0)); forvar4374 = (forvar4374 + (1'h1)))
            begin
              if (reg4383[(1'h0):(1'h0)])
                begin
                  for (forvar4375 = (1'h0); (forvar4375 < (2'h2)); forvar4375 = (forvar4375 + (1'h1)))
                    begin
                      reg4376 <= (!{($signed(reg4328) << (reg4381 && reg4357))});
                      reg4377 <= ((8'hb7) * $unsigned((-forvar4375[(1'h1):(1'h1)])));
                      reg4378 <= $unsigned((!((^(8'hb7)) >>> $unsigned(reg4377))));
                      reg4379 <= {{(reg4376[(2'h3):(1'h0)] == (!(8'ha7)))}};
                    end
                  for (forvar4380 = (1'h0); (forvar4380 < (1'h1)); forvar4380 = (forvar4380 + (1'h1)))
                    begin
                      reg4381 <= $signed({$signed($signed((8'ha7)))});
                    end
                  if ((&reg4339))
                    begin
                      reg4382 <= $unsigned(((~reg4367[(3'h5):(3'h5)]) ?
                          $unsigned((reg4348 != reg4351)) : {wire4319}));
                    end
                  else
                    begin
                      reg4382 <= reg4332;
                    end
                  for (forvar4383 = (1'h0); (forvar4383 < (1'h0)); forvar4383 = (forvar4383 + (1'h1)))
                    begin
                      reg4384 <= $unsigned((wire4318 ?
                          reg4337[(4'h9):(3'h5)] : ((&reg4381) >= (wire4319 & forvar4376))));
                      reg4385 <= reg4394[(2'h3):(1'h1)];
                      reg4386 <= ($signed((^~(forvar4376 ?
                          reg4338 : wire2))) * (reg4345[(2'h2):(2'h2)] < ($unsigned(reg4369) && $signed(reg4389))));
                    end
                end
              else
                begin
                  if (reg4355[(1'h0):(1'h0)])
                    begin
                      reg4375 <= ((((&reg4365) ?
                                  reg4367[(2'h2):(2'h2)] : ((8'hb0) >>> reg4394)) ?
                              reg4351[(1'h0):(1'h0)] : reg4381) ?
                          (~&$unsigned($signed(reg4356))) : $signed(((^(8'hb8)) ?
                              $signed(reg4400) : reg4327)));
                      reg4376 <= (+reg4383[(1'h0):(1'h0)]);
                      reg4377 <= (|$signed($unsigned((reg4349 >= forvar4392))));
                    end
                  else
                    begin
                      reg4375 <= ((reg4343 ?
                              ((reg4349 && reg4360) ?
                                  {reg4355} : $signed(reg4356)) : $unsigned($unsigned(reg4322))) ?
                          reg4363 : reg4367[(3'h6):(1'h0)]);
                    end
                  if ($unsigned(reg4375[(4'hf):(3'h5)]))
                    begin
                      reg4378 <= (reg4391 ?
                          ((^$unsigned((8'h9c))) != $signed((~^reg4387))) : reg4360);
                    end
                  else
                    begin
                      reg4378 <= $signed(forvar4383[(1'h1):(1'h1)]);
                      reg4379 <= reg4335[(4'h9):(1'h0)];
                      reg4380 <= $signed(reg4388[(3'h7):(3'h4)]);
                    end
                end
            end
        end
      for (forvar4402 = (1'h0); (forvar4402 < (1'h1)); forvar4402 = (forvar4402 + (1'h1)))
        begin
          for (forvar4403 = (1'h0); (forvar4403 < (1'h1)); forvar4403 = (forvar4403 + (1'h1)))
            begin
              if ($unsigned((~(~&wire4316[(3'h4):(2'h3)]))))
                begin
                  reg4404 <= $unsigned(reg4367[(2'h3):(2'h2)]);
                  for (forvar4405 = (1'h0); (forvar4405 < (1'h0)); forvar4405 = (forvar4405 + (1'h1)))
                    begin
                      reg4406 <= $signed($signed((^~$signed(reg4346))));
                      reg4407 <= reg4357[(1'h0):(1'h0)];
                    end
                  reg4408 <= (-((|reg4330) - $signed($signed(reg4347))));
                  reg4409 <= ($unsigned(wire4316[(4'hd):(1'h0)]) <<< reg4399);
                end
              else
                begin
                  reg4404 <= forvar4396[(4'h9):(2'h3)];
                  reg4405 <= $signed((^~$signed((!reg4365))));
                  reg4406 <= $unsigned({$signed($signed(reg4342))});
                  if ($signed(wire1))
                    begin
                      reg4407 <= reg4375[(4'hc):(4'hc)];
                      reg4408 <= ((reg4393 ?
                              (8'hae) : $signed((forvar4383 << (8'ha6)))) ?
                          $signed(reg4373) : (reg4381[(2'h2):(1'h1)] > ($unsigned((8'ha0)) * forvar4376[(3'h6):(2'h2)])));
                      reg4409 <= $unsigned({((8'hb0) ?
                              wire4316[(4'hc):(1'h0)] : reg4352)});
                    end
                  else
                    begin
                      reg4407 <= (reg4351[(2'h3):(1'h1)] >> (reg4359[(2'h2):(1'h0)] == $signed(reg4377)));
                      reg4408 <= (+(~|$signed($signed(reg4365))));
                      reg4409 <= {(reg4364 + $signed(reg4357))};
                    end
                end
            end
          for (forvar4410 = (1'h0); (forvar4410 < (1'h0)); forvar4410 = (forvar4410 + (1'h1)))
            begin
              if (({reg4334} | $unsigned((|$signed(reg4399)))))
                begin
                  reg4411 <= reg4350[(4'hd):(1'h0)];
                  if (reg4380[(2'h2):(1'h1)])
                    begin
                      reg4412 <= (((((8'ha9) ? reg4349 : reg4355) ~^ reg4387) ?
                          {reg4350[(3'h6):(3'h6)]} : ((reg4409 ^ reg4358) ^ {reg4369})) << (^~$signed((reg4370 ?
                          wire4320 : (8'ha2)))));
                    end
                  else
                    begin
                      reg4412 <= forvar4402;
                      reg4413 <= reg4362[(4'h8):(3'h7)];
                      reg4414 <= $signed((reg4377 == {(reg4327 ?
                              (8'haf) : forvar4375)}));
                    end
                end
              else
                begin
                  for (forvar4411 = (1'h0); (forvar4411 < (1'h0)); forvar4411 = (forvar4411 + (1'h1)))
                    begin
                      reg4412 <= (~^(8'hb4));
                      reg4413 <= ($unsigned(((&reg4342) ?
                              $unsigned((8'ha5)) : forvar4376)) ?
                          (~&((^~wire4318) << (forvar4376 ?
                              reg4339 : reg4365))) : reg4358[(2'h3):(1'h1)]);
                      reg4414 <= $signed(($signed((^reg4376)) >= (~&wire4320[(4'h8):(2'h3)])));
                    end
                  reg4415 <= {$signed((&((8'ha0) <<< reg4356)))};
                end
              for (forvar4416 = (1'h0); (forvar4416 < (1'h0)); forvar4416 = (forvar4416 + (1'h1)))
                begin
                  for (forvar4417 = (1'h0); (forvar4417 < (1'h1)); forvar4417 = (forvar4417 + (1'h1)))
                    begin
                      reg4418 <= reg4333;
                      reg4419 <= forvar4410[(2'h2):(1'h0)];
                    end
                  for (forvar4420 = (1'h0); (forvar4420 < (2'h3)); forvar4420 = (forvar4420 + (1'h1)))
                    begin
                      reg4421 <= (8'ha7);
                      reg4422 <= {(8'hac)};
                      reg4423 <= (({(reg4348 >> reg4366)} > forvar4411[(4'h9):(3'h7)]) >>> $unsigned({reg4405[(1'h0):(1'h0)]}));
                      reg4424 <= ((~&(~(reg4347 <<< reg4379))) ^ (reg4342[(3'h4):(3'h4)] ?
                          ((reg4423 >>> (8'hb0)) ?
                              reg4355[(3'h7):(1'h1)] : (reg4334 ?
                                  (8'hb1) : wire0)) : (^{reg4413})));
                    end
                  for (forvar4425 = (1'h0); (forvar4425 < (2'h3)); forvar4425 = (forvar4425 + (1'h1)))
                    begin
                      reg4426 <= reg4376;
                      reg4427 <= $signed($signed(reg4334[(1'h0):(1'h0)]));
                    end
                end
            end
          for (forvar4428 = (1'h0); (forvar4428 < (1'h1)); forvar4428 = (forvar4428 + (1'h1)))
            begin
              for (forvar4429 = (1'h0); (forvar4429 < (2'h2)); forvar4429 = (forvar4429 + (1'h1)))
                begin
                  if ((reg4414[(3'h7):(3'h4)] ?
                      $unsigned($signed((reg4344 >>> reg4423))) : $signed($unsigned({forvar4375}))))
                    begin
                      reg4430 <= ($signed($signed(reg4352)) >> forvar4410);
                      reg4431 <= reg4330;
                      reg4432 <= ($unsigned(forvar4417[(4'hd):(3'h4)]) ?
                          $signed($signed({forvar4416})) : reg4390);
                    end
                  else
                    begin
                      reg4430 <= ($unsigned(reg4371[(2'h3):(1'h1)]) - reg4404);
                      reg4431 <= reg4373[(4'h8):(3'h5)];
                      reg4432 <= ((((reg4334 ?
                          reg4370 : (8'h9d)) && reg4404) | forvar4403[(4'ha):(3'h5)]) + {(wire4316 - {(8'had)})});
                      reg4433 <= $signed($signed($signed($unsigned(reg4422))));
                    end
                  if ((reg4433[(1'h1):(1'h0)] <= $unsigned(wire3[(3'h7):(3'h6)])))
                    begin
                      reg4434 <= $unsigned((+$unsigned(reg4409[(3'h7):(3'h4)])));
                      reg4435 <= (($unsigned(reg4351[(2'h3):(1'h0)]) ?
                              reg4366 : (8'hb2)) ?
                          (^~{(reg4349 >= reg4328)}) : (reg4341 ?
                              $signed(reg4406[(1'h1):(1'h1)]) : (8'hac)));
                      reg4436 <= (forvar4416[(2'h3):(2'h3)] != reg4336[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg4434 <= reg4393[(3'h4):(2'h2)];
                      reg4435 <= (~&reg4384[(1'h1):(1'h0)]);
                      reg4436 <= (reg4383 ? (8'hb0) : forvar4416);
                      reg4437 <= $signed(((reg4340 * (8'hb8)) ?
                          (~|(reg4409 ?
                              reg4355 : (8'hb0))) : reg4356[(2'h3):(2'h3)]));
                    end
                  for (forvar4438 = (1'h0); (forvar4438 < (1'h0)); forvar4438 = (forvar4438 + (1'h1)))
                    begin
                      reg4439 <= (~($signed((~|reg4345)) ?
                          forvar4396 : ((reg4345 >> forvar4429) > (reg4394 + reg4400))));
                      reg4440 <= reg4380;
                      reg4441 <= ((reg4322 != $unsigned((reg4349 >>> forvar4416))) || wire4320);
                    end
                end
              for (forvar4442 = (1'h0); (forvar4442 < (2'h2)); forvar4442 = (forvar4442 + (1'h1)))
                begin
                  for (forvar4443 = (1'h0); (forvar4443 < (1'h0)); forvar4443 = (forvar4443 + (1'h1)))
                    begin
                      reg4444 <= $signed(reg4331[(2'h2):(1'h1)]);
                      reg4445 <= {reg4411};
                      reg4446 <= ((wire4318[(4'hc):(1'h0)] << $signed((reg4385 ?
                              (8'hb3) : reg4401))) ?
                          reg4322 : ($unsigned((reg4376 - reg4333)) ?
                              ((reg4399 ? forvar4410 : wire4318) ?
                                  (-reg4375) : $signed((8'h9e))) : $unsigned((reg4345 << reg4339))));
                      reg4447 <= (+reg4379[(4'hf):(4'hb)]);
                    end
                  for (forvar4448 = (1'h0); (forvar4448 < (1'h1)); forvar4448 = (forvar4448 + (1'h1)))
                    begin
                      reg4449 <= $unsigned((~|reg4393[(1'h0):(1'h0)]));
                    end
                  if (reg4358)
                    begin
                      reg4450 <= reg4401;
                      reg4451 <= reg4406;
                      reg4452 <= $unsigned(({$signed(reg4409)} > $unsigned({wire4316})));
                      reg4453 <= (((^$unsigned((8'ha0))) - ((~&forvar4402) ?
                          $signed(wire1) : (reg4388 - wire3))) == $unsigned((reg4394 || (reg4419 <= reg4341))));
                    end
                  else
                    begin
                      reg4450 <= ((|(~|(reg4407 | reg4414))) ?
                          (^(8'hb7)) : {(~^$signed(forvar4392))});
                      reg4451 <= ((8'hb3) ? reg4343 : wire2);
                      reg4452 <= reg4362[(3'h7):(3'h7)];
                    end
                  for (forvar4454 = (1'h0); (forvar4454 < (2'h3)); forvar4454 = (forvar4454 + (1'h1)))
                    begin
                      reg4455 <= (((~^reg4332[(3'h5):(1'h0)]) ?
                          $unsigned((!reg4407)) : $unsigned(reg4369[(2'h2):(2'h2)])) | (|(~^(reg4352 ?
                          reg4398 : reg4357))));
                      reg4456 <= $signed(reg4455[(1'h0):(1'h0)]);
                      reg4457 <= ((8'ha9) ^ ($unsigned((~^forvar4403)) >> (|$signed(reg4367))));
                    end
                end
            end
        end
      for (forvar4458 = (1'h0); (forvar4458 < (1'h0)); forvar4458 = (forvar4458 + (1'h1)))
        begin
          for (forvar4459 = (1'h0); (forvar4459 < (2'h3)); forvar4459 = (forvar4459 + (1'h1)))
            begin
              reg4460 <= $unsigned(reg4431[(3'h5):(3'h5)]);
            end
        end
      if ((($unsigned(reg4400) ?
              $signed(((8'hb5) + reg4391)) : (^(reg4419 >= reg4370))) ?
          $signed((!(forvar4402 ? reg4452 : reg4322))) : (((+reg4451) ?
              (~&forvar4403) : reg4408[(1'h0):(1'h0)]) >> {{wire4318}})))
        begin
          if (((~|reg4376) ?
              ((reg4391 <<< reg4359[(2'h2):(2'h2)]) != ((^~reg4452) ?
                  reg4322[(2'h3):(1'h1)] : (reg4419 ?
                      reg4386 : reg4411))) : reg4430[(1'h1):(1'h0)]))
            begin
              if ((&(8'hb8)))
                begin
                  if (forvar4443[(4'hb):(3'h6)])
                    begin
                      reg4461 <= (~reg4328);
                      reg4462 <= reg4431;
                    end
                  else
                    begin
                      reg4461 <= (&reg4336[(2'h3):(2'h2)]);
                      reg4462 <= reg4390[(2'h3):(1'h0)];
                      reg4463 <= (({(reg4342 ? reg4393 : (8'hb1))} ?
                              (reg4342[(3'h4):(2'h2)] >= reg4353[(2'h3):(2'h3)]) : reg4444[(3'h4):(2'h2)]) ?
                          ($signed(wire1) ?
                              ({reg4336} ?
                                  reg4362[(2'h3):(1'h0)] : (8'h9f)) : reg4411[(1'h1):(1'h0)]) : reg4369[(1'h1):(1'h1)]);
                      reg4464 <= reg4373;
                    end
                end
              else
                begin
                  for (forvar4461 = (1'h0); (forvar4461 < (1'h1)); forvar4461 = (forvar4461 + (1'h1)))
                    begin
                      reg4462 <= $signed((-reg4354[(3'h5):(1'h0)]));
                      reg4463 <= forvar4392;
                      reg4464 <= ((reg4390 || reg4324[(1'h1):(1'h1)]) ?
                          reg4342[(1'h1):(1'h0)] : $unsigned(reg4370[(3'h6):(1'h0)]));
                    end
                  for (forvar4465 = (1'h0); (forvar4465 < (2'h2)); forvar4465 = (forvar4465 + (1'h1)))
                    begin
                      reg4466 <= forvar4438[(3'h7):(3'h6)];
                    end
                  for (forvar4467 = (1'h0); (forvar4467 < (2'h3)); forvar4467 = (forvar4467 + (1'h1)))
                    begin
                      reg4468 <= reg4456[(3'h6):(3'h5)];
                      reg4469 <= (~^(!reg4379));
                    end
                  for (forvar4470 = (1'h0); (forvar4470 < (1'h0)); forvar4470 = (forvar4470 + (1'h1)))
                    begin
                      reg4471 <= ((reg4398[(4'h9):(2'h3)] && $signed((8'hb7))) ?
                          ($unsigned($signed(forvar4459)) ?
                              forvar4420 : (~|{wire4319})) : $unsigned($signed({reg4322})));
                    end
                end
              if ($unsigned((^reg4390[(1'h0):(1'h0)])))
                begin
                  for (forvar4472 = (1'h0); (forvar4472 < (2'h2)); forvar4472 = (forvar4472 + (1'h1)))
                    begin
                      reg4473 <= ({reg4453[(3'h7):(3'h6)]} >>> reg4345[(4'ha):(4'h8)]);
                      reg4474 <= ($unsigned($unsigned(reg4460)) ?
                          $signed(((reg4380 <= reg4375) ?
                              {(8'hb4)} : (reg4373 <<< reg4426))) : (((reg4367 && reg4342) ?
                                  {reg4369} : (|reg4327)) ?
                              (+{reg4391}) : $unsigned(reg4435)));
                      reg4475 <= $signed(($signed({reg4364}) ?
                          (^~(|reg4400)) : ((^~reg4415) ?
                              $unsigned(forvar4458) : (~reg4353))));
                    end
                end
              else
                begin
                  if ((8'ha2))
                    begin
                      reg4472 <= $unsigned((reg4348 >> {{reg4348}}));
                      reg4473 <= $unsigned((reg4371[(4'he):(2'h3)] ?
                          (reg4434[(3'h4):(2'h3)] >= (reg4372 ?
                              reg4419 : reg4399)) : reg4457[(3'h6):(1'h0)]));
                      reg4474 <= {($signed((reg4331 ^ reg4357)) > (&reg4337[(5'h10):(4'he)]))};
                      reg4475 <= $signed({$unsigned((8'ha1))});
                    end
                  else
                    begin
                      reg4472 <= (forvar4458 ?
                          reg4418 : $unsigned((^$unsigned(reg4384))));
                    end
                end
              if (({$unsigned((reg4365 << reg4345))} ?
                  $unsigned(reg4352[(2'h2):(1'h0)]) : ((8'h9f) >> reg4340)))
                begin
                  for (forvar4476 = (1'h0); (forvar4476 < (2'h3)); forvar4476 = (forvar4476 + (1'h1)))
                    begin
                      reg4477 <= ((~&reg4334[(4'h9):(3'h5)]) ?
                          reg4358[(2'h3):(2'h2)] : reg4367[(1'h1):(1'h0)]);
                      reg4478 <= $unsigned($unsigned(reg4439));
                      reg4479 <= (-$unsigned(reg4346[(3'h5):(1'h1)]));
                    end
                  reg4480 <= {wire2[(2'h2):(2'h2)]};
                  reg4481 <= reg4426;
                  reg4482 <= (+$unsigned(({reg4408} < $unsigned(reg4456))));
                end
              else
                begin
                  if (forvar4405[(3'h7):(3'h4)])
                    begin
                      reg4476 <= ({((8'hb7) + (&reg4371))} ?
                          $unsigned(reg4389) : wire2);
                      reg4477 <= (($unsigned({forvar4459}) ?
                          $signed(reg4332[(1'h1):(1'h1)]) : (forvar4417 ?
                              (reg4394 << (8'ha5)) : $unsigned(reg4367))) + ($unsigned(reg4338) ?
                          reg4378 : $signed((reg4393 <<< reg4381))));
                    end
                  else
                    begin
                      reg4476 <= reg4333;
                      reg4477 <= $unsigned($unsigned($unsigned({reg4351})));
                    end
                  if (reg4371)
                    begin
                      reg4478 <= ((((~reg4463) >>> $signed(reg4435)) ?
                              reg4399[(4'hc):(3'h7)] : (reg4362 ?
                                  $unsigned(reg4365) : $signed(reg4362))) ?
                          {((reg4322 >= (8'haf)) >> reg4373)} : $signed($signed((~&wire2))));
                    end
                  else
                    begin
                      reg4478 <= $unsigned($unsigned($signed(reg4473)));
                      reg4479 <= reg4476[(3'h7):(2'h3)];
                    end
                end
              reg4483 <= forvar4461[(2'h3):(2'h3)];
            end
          else
            begin
              reg4461 <= (~&reg4431);
              for (forvar4462 = (1'h0); (forvar4462 < (2'h2)); forvar4462 = (forvar4462 + (1'h1)))
                begin
                  reg4463 <= reg4371;
                  if ((~^({reg4407[(3'h4):(1'h1)]} ?
                      {$unsigned(forvar4396)} : (reg4340[(1'h1):(1'h1)] ?
                          reg4369[(3'h4):(2'h2)] : {reg4387}))))
                    begin
                      reg4464 <= ($unsigned(reg4357) ?
                          ($unsigned({reg4480}) < reg4482) : {({reg4434} != (forvar4374 > reg4330))});
                    end
                  else
                    begin
                      reg4464 <= $signed((+(reg4483 >>> reg4358)));
                    end
                  if ($unsigned((~reg4332[(3'h4):(3'h4)])))
                    begin
                      reg4465 <= reg4342;
                      reg4466 <= $unsigned(forvar4467);
                      reg4467 <= $signed((reg4335 != $unsigned({(8'ha5)})));
                      reg4468 <= (($signed((reg4376 ~^ forvar4402)) == reg4349) ?
                          ($signed(reg4480[(2'h2):(1'h0)]) ?
                              reg4400[(1'h1):(1'h1)] : ($signed(forvar4428) ?
                                  (~reg4322) : wire4319)) : reg4451);
                    end
                  else
                    begin
                      reg4465 <= (((^~reg4324) < forvar4375[(1'h1):(1'h0)]) != $unsigned((~^(wire3 & reg4371))));
                      reg4466 <= forvar4416;
                    end
                end
            end
        end
      else
        begin
          if ((reg4367 ? reg4439[(1'h0):(1'h0)] : {(8'h9d)}))
            begin
              for (forvar4461 = (1'h0); (forvar4461 < (2'h2)); forvar4461 = (forvar4461 + (1'h1)))
                begin
                  reg4462 <= {reg4466};
                  reg4463 <= reg4388;
                  for (forvar4464 = (1'h0); (forvar4464 < (1'h1)); forvar4464 = (forvar4464 + (1'h1)))
                    begin
                      reg4465 <= (8'hb7);
                      reg4466 <= {wire3[(4'ha):(3'h4)]};
                      reg4467 <= reg4353;
                      reg4468 <= (~&reg4432[(1'h1):(1'h1)]);
                    end
                  reg4469 <= $unsigned(((~{reg4338}) ?
                      reg4387[(3'h5):(1'h1)] : {reg4328}));
                end
              for (forvar4470 = (1'h0); (forvar4470 < (1'h1)); forvar4470 = (forvar4470 + (1'h1)))
                begin
                  reg4471 <= reg4355;
                  reg4472 <= wire1;
                end
              for (forvar4473 = (1'h0); (forvar4473 < (1'h1)); forvar4473 = (forvar4473 + (1'h1)))
                begin
                  for (forvar4474 = (1'h0); (forvar4474 < (1'h0)); forvar4474 = (forvar4474 + (1'h1)))
                    begin
                      reg4475 <= $unsigned({$unsigned({reg4412})});
                      reg4476 <= reg4332;
                      reg4477 <= reg4381[(3'h6):(2'h2)];
                    end
                end
            end
          else
            begin
              if ((reg4401 <= (-(^$unsigned(forvar4467)))))
                begin
                  reg4461 <= {((-((8'had) ? reg4388 : reg4358)) ?
                          reg4480[(1'h1):(1'h0)] : {$unsigned(reg4418)})};
                end
              else
                begin
                  if (reg4460[(1'h0):(1'h0)])
                    begin
                      reg4461 <= $unsigned(($unsigned(forvar4448[(2'h3):(2'h2)]) || $signed((reg4347 ?
                          (8'hb1) : reg4359))));
                      reg4462 <= {($unsigned(reg4466[(4'ha):(4'h9)]) ?
                              (!(reg4434 == reg4465)) : {reg4364[(1'h0):(1'h0)]})};
                      reg4463 <= (|$signed($unsigned(((8'ha7) >> reg4351))));
                      reg4464 <= forvar4392;
                    end
                  else
                    begin
                      reg4461 <= reg4430[(3'h4):(2'h2)];
                      reg4462 <= $signed((reg4460 + reg4447[(3'h4):(1'h0)]));
                      reg4463 <= reg4357;
                    end
                  for (forvar4465 = (1'h0); (forvar4465 < (1'h0)); forvar4465 = (forvar4465 + (1'h1)))
                    begin
                      reg4466 <= $signed((~&($signed(forvar4448) + (reg4445 ?
                          reg4407 : (8'haf)))));
                    end
                end
            end
          for (forvar4478 = (1'h0); (forvar4478 < (1'h0)); forvar4478 = (forvar4478 + (1'h1)))
            begin
              if ($unsigned($signed($unsigned({forvar4376}))))
                begin
                  if (((+((reg4444 ? reg4423 : reg4336) ?
                      (forvar4464 >> (8'ha5)) : reg4351[(2'h3):(2'h2)])) != $unsigned($signed($signed((8'ha2))))))
                    begin
                      reg4479 <= forvar4392;
                      reg4480 <= reg4400;
                      reg4481 <= ($unsigned($signed(reg4386)) ?
                          {(+(8'hb2))} : reg4419[(3'h6):(2'h3)]);
                      reg4482 <= ({($unsigned(reg4476) ?
                                  {forvar4416} : $signed(reg4390))} ?
                          {(-reg4449[(1'h1):(1'h0)])} : (reg4391[(4'h9):(3'h5)] ?
                              reg4354[(3'h5):(1'h0)] : ((8'ha0) ?
                                  $signed(reg4364) : (~&reg4375))));
                    end
                  else
                    begin
                      reg4479 <= $unsigned(($signed((|reg4338)) ?
                          $unsigned(reg4345[(3'h7):(3'h5)]) : (~&reg4359[(3'h4):(1'h0)])));
                      reg4480 <= ((~&(((8'ha8) | reg4479) < $signed(reg4414))) ?
                          $unsigned($signed(forvar4396)) : $unsigned((&$signed(forvar4464))));
                      reg4481 <= ((^~(8'hb4)) + ((wire3 ?
                          reg4431 : (reg4424 << reg4433)) || reg4368[(2'h3):(2'h3)]));
                    end
                  if (reg4457[(4'hc):(4'h9)])
                    begin
                      reg4483 <= ({($signed((8'h9e)) || {(8'hb2)})} ?
                          reg4397[(4'ha):(2'h2)] : ((reg4385[(3'h4):(1'h1)] < reg4327) ?
                              wire2[(2'h2):(1'h0)] : reg4418));
                    end
                  else
                    begin
                      reg4483 <= (reg4408[(3'h4):(1'h1)] ?
                          forvar4403 : $unsigned({(forvar4417 && reg4385)}));
                      reg4484 <= (8'ha1);
                    end
                  if (reg4451)
                    begin
                      reg4485 <= ($signed($unsigned($signed(reg4467))) <= reg4395);
                      reg4486 <= {$unsigned((reg4369[(3'h4):(1'h0)] ^~ (~&forvar4478)))};
                    end
                  else
                    begin
                      reg4485 <= (($unsigned(reg4327) * reg4476) ?
                          $signed($signed(reg4447[(3'h5):(2'h2)])) : (forvar4448 ?
                              (-wire4318) : (~|{(8'hab)})));
                    end
                end
              else
                begin
                  for (forvar4479 = (1'h0); (forvar4479 < (2'h2)); forvar4479 = (forvar4479 + (1'h1)))
                    begin
                      reg4480 <= $unsigned(((reg4474[(3'h5):(2'h2)] ?
                              $unsigned(reg4444) : reg4476[(4'h8):(4'h8)]) ?
                          $unsigned((!forvar4467)) : ($signed(reg4456) ?
                              $unsigned((8'hb5)) : ((8'ha6) ?
                                  reg4383 : forvar4479))));
                    end
                  if ((((|(forvar4438 ? reg4387 : reg4445)) ?
                          (reg4331[(2'h3):(1'h0)] + (^reg4387)) : {(reg4335 ?
                                  reg4477 : (8'h9f))}) ?
                      $signed((reg4338 ?
                          (reg4473 ?
                              reg4358 : reg4400) : (~^(8'hb1)))) : $unsigned(((reg4404 ?
                          reg4342 : wire1) >= $unsigned(reg4362)))))
                    begin
                      reg4481 <= $unsigned((reg4414[(2'h3):(1'h1)] & reg4445[(1'h0):(1'h0)]));
                      reg4482 <= reg4445[(1'h0):(1'h0)];
                      reg4483 <= $unsigned(reg4376);
                    end
                  else
                    begin
                      reg4481 <= reg4476[(2'h3):(2'h2)];
                    end
                  for (forvar4484 = (1'h0); (forvar4484 < (1'h1)); forvar4484 = (forvar4484 + (1'h1)))
                    begin
                      reg4485 <= forvar4376[(2'h3):(2'h3)];
                      reg4486 <= (~reg4411);
                    end
                  reg4487 <= forvar4448[(4'hc):(3'h4)];
                end
              for (forvar4488 = (1'h0); (forvar4488 < (1'h0)); forvar4488 = (forvar4488 + (1'h1)))
                begin
                  reg4489 <= $unsigned((((8'h9e) >>> $signed(forvar4461)) ?
                      $unsigned((reg4389 << (8'hb2))) : reg4395));
                end
              for (forvar4490 = (1'h0); (forvar4490 < (2'h2)); forvar4490 = (forvar4490 + (1'h1)))
                begin
                  if ((&({reg4427} ~^ reg4362[(3'h5):(1'h0)])))
                    begin
                      reg4491 <= $signed({$unsigned((reg4356 & wire1))});
                      reg4492 <= (reg4363[(3'h4):(2'h3)] || (($unsigned(reg4337) | (reg4480 ?
                          reg4393 : forvar4442)) && $signed((reg4419 ?
                          (8'hb3) : (8'ha3)))));
                      reg4493 <= (forvar4405 ? {(8'ha1)} : (~&forvar4374));
                    end
                  else
                    begin
                      reg4491 <= reg4372[(2'h2):(1'h0)];
                      reg4492 <= (((reg4483[(3'h4):(3'h4)] ?
                                  (reg4465 >= forvar4374) : (~^(8'h9e))) ?
                              reg4436[(3'h5):(2'h2)] : (reg4341[(3'h5):(3'h4)] ^ (+forvar4448))) ?
                          (&reg4351[(3'h5):(1'h1)]) : (forvar4411[(1'h1):(1'h1)] ?
                              $signed(reg4397) : (|wire4316[(4'hc):(4'h9)])));
                    end
                end
              reg4494 <= (8'hb1);
            end
          if (reg4340)
            begin
              for (forvar4495 = (1'h0); (forvar4495 < (1'h1)); forvar4495 = (forvar4495 + (1'h1)))
                begin
                  reg4496 <= reg4339;
                  reg4497 <= $unsigned((&((reg4393 >>> forvar4473) ?
                      $signed(reg4476) : $signed(reg4333))));
                end
              for (forvar4498 = (1'h0); (forvar4498 < (1'h1)); forvar4498 = (forvar4498 + (1'h1)))
                begin
                  if (reg4336)
                    begin
                      reg4499 <= ((&reg4384[(1'h0):(1'h0)]) ?
                          ($unsigned((&reg4353)) ?
                              $signed(forvar4448[(2'h3):(2'h2)]) : (reg4375 ?
                                  reg4348 : (~reg4381))) : (reg4384 | {$signed(forvar4498)}));
                      reg4500 <= ((((reg4451 ?
                                  forvar4498 : reg4387) >>> $unsigned(forvar4429)) ?
                              {$unsigned(forvar4488)} : (reg4345[(4'hb):(2'h3)] ?
                                  $unsigned(reg4347) : (reg4441 ?
                                      reg4418 : forvar4438))) ?
                          forvar4383[(2'h2):(1'h1)] : ($signed($unsigned((8'haa))) >> $signed($unsigned((8'ha1)))));
                      reg4501 <= reg4334;
                    end
                  else
                    begin
                      reg4499 <= forvar4498[(1'h1):(1'h0)];
                      reg4500 <= reg4462[(2'h3):(2'h3)];
                      reg4501 <= (({forvar4405} ?
                              ((forvar4403 ? reg4352 : forvar4392) ~^ (reg4471 ?
                                  reg4370 : reg4475)) : (forvar4392 ?
                                  (reg4451 && reg4491) : (reg4424 ^ reg4355))) ?
                          $signed(reg4411[(1'h0):(1'h0)]) : wire4316[(3'h6):(2'h2)]);
                    end
                  reg4502 <= {(((reg4460 ? reg4355 : forvar4383) ?
                          forvar4429 : $unsigned(wire4316)) * (&$unsigned(reg4435)))};
                  for (forvar4503 = (1'h0); (forvar4503 < (2'h3)); forvar4503 = (forvar4503 + (1'h1)))
                    begin
                      reg4504 <= $signed($signed($signed(((8'ha6) ?
                          (8'hb2) : forvar4479))));
                      reg4505 <= $signed((|($unsigned(reg4354) ?
                          (forvar4442 ? reg4411 : reg4334) : reg4331)));
                      reg4506 <= (($unsigned((8'hb2)) ?
                          (&(-reg4349)) : {$signed(reg4451)}) >> {(^~$unsigned(reg4376))});
                      reg4507 <= ({reg4327} ?
                          (reg4432[(1'h1):(1'h0)] ?
                              (~forvar4461[(4'h8):(2'h3)]) : $unsigned((reg4358 ?
                                  reg4483 : reg4486))) : reg4465);
                    end
                end
              for (forvar4508 = (1'h0); (forvar4508 < (2'h2)); forvar4508 = (forvar4508 + (1'h1)))
                begin
                  if (reg4327[(2'h2):(2'h2)])
                    begin
                      reg4509 <= reg4393;
                    end
                  else
                    begin
                      reg4509 <= (reg4418[(2'h3):(2'h2)] != $unsigned((-forvar4479[(2'h3):(1'h1)])));
                    end
                  if ($signed($signed(reg4501)))
                    begin
                      reg4510 <= (8'ha3);
                      reg4511 <= (~$unsigned($signed($unsigned(reg4355))));
                      reg4512 <= (^(~|$signed((~^reg4476))));
                      reg4513 <= reg4509;
                    end
                  else
                    begin
                      reg4510 <= (^~(reg4431 ?
                          (forvar4383 == reg4451) : reg4427[(3'h4):(3'h4)]));
                      reg4511 <= ((({reg4486} > reg4370) >>> reg4359[(2'h2):(1'h1)]) >= reg4365);
                      reg4512 <= reg4466[(4'h9):(1'h1)];
                    end
                  if ((8'h9c))
                    begin
                      reg4514 <= reg4422;
                      reg4515 <= ($signed(((reg4475 * forvar4429) <= (reg4393 >> reg4355))) ?
                          {reg4467} : (reg4372 >= (^~reg4358)));
                      reg4516 <= reg4381[(3'h5):(1'h1)];
                      reg4517 <= ($signed((reg4363 ?
                              (reg4357 | reg4476) : $signed(reg4397))) ?
                          (~^$signed($signed((8'hb6)))) : reg4369[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg4514 <= {reg4413};
                    end
                end
            end
          else
            begin
              reg4495 <= $unsigned(({$unsigned(reg4414)} ?
                  (reg4372 << (reg4436 ?
                      reg4411 : (8'h9c))) : (^reg4358[(1'h0):(1'h0)])));
            end
        end
    end
  assign wire4518 = $unsigned(reg4370[(2'h3):(2'h2)]);
  always
    @(posedge clk) begin
      for (forvar4519 = (1'h0); (forvar4519 < (1'h1)); forvar4519 = (forvar4519 + (1'h1)))
        begin
          for (forvar4520 = (1'h0); (forvar4520 < (2'h3)); forvar4520 = (forvar4520 + (1'h1)))
            begin
              if ((~|{($signed(reg4506) ? (reg4386 + reg4437) : reg4340)}))
                begin
                  for (forvar4521 = (1'h0); (forvar4521 < (2'h3)); forvar4521 = (forvar4521 + (1'h1)))
                    begin
                      reg4522 <= $signed($signed($signed(reg4352[(1'h1):(1'h1)])));
                      reg4523 <= wire2;
                    end
                  if ((-$unsigned(reg4463)))
                    begin
                      reg4524 <= $unsigned((($signed(reg4371) && $unsigned(reg4477)) >> ({reg4511} ?
                          reg4475[(3'h4):(2'h3)] : (-reg4479))));
                    end
                  else
                    begin
                      reg4524 <= (reg4446 ?
                          (+$unsigned(reg4411)) : {(-(reg4449 ?
                                  reg4500 : reg4423))});
                      reg4525 <= reg4343[(4'hb):(4'h8)];
                    end
                  for (forvar4526 = (1'h0); (forvar4526 < (2'h2)); forvar4526 = (forvar4526 + (1'h1)))
                    begin
                      reg4527 <= $signed(reg4450);
                    end
                end
              else
                begin
                  reg4521 <= reg4486;
                  if ($unsigned(reg4523))
                    begin
                      reg4522 <= reg4430[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg4522 <= reg4406[(3'h5):(2'h2)];
                    end
                end
            end
          if (reg4460[(3'h4):(2'h3)])
            begin
              if ($signed((~reg4328)))
                begin
                  if ($signed((($unsigned(reg4358) ?
                          $unsigned(reg4475) : (|reg4475)) ?
                      (8'ha6) : (^reg4354))))
                    begin
                      reg4528 <= reg4406[(3'h4):(3'h4)];
                      reg4529 <= reg4412[(2'h3):(1'h1)];
                      reg4530 <= $unsigned(reg4493[(3'h7):(3'h5)]);
                    end
                  else
                    begin
                      reg4528 <= (~^{$signed((reg4360 ? (8'ha3) : reg4457))});
                      reg4529 <= ((~(8'ha7)) >= ($signed($signed(reg4489)) ?
                          ((^~reg4510) ?
                              (~|reg4433) : reg4407) : {$unsigned(reg4460)}));
                      reg4530 <= reg4451[(1'h0):(1'h0)];
                      reg4531 <= ((+reg4386) - (reg4445[(3'h6):(3'h5)] ^~ reg4387));
                    end
                end
              else
                begin
                  for (forvar4528 = (1'h0); (forvar4528 < (2'h3)); forvar4528 = (forvar4528 + (1'h1)))
                    begin
                      reg4529 <= (((~|reg4389) ?
                              $signed({reg4360}) : ($signed(reg4394) ?
                                  reg4332 : $signed(wire3))) ?
                          forvar4519 : ($signed((reg4489 * reg4341)) ?
                              (~^{reg4446}) : reg4405));
                    end
                end
              for (forvar4532 = (1'h0); (forvar4532 < (1'h0)); forvar4532 = (forvar4532 + (1'h1)))
                begin
                  reg4533 <= ($signed(($signed(forvar4528) ~^ (reg4322 || reg4484))) >= (({reg4427} ?
                          {(8'hb9)} : reg4343) ?
                      $signed((^reg4460)) : {((8'hb0) ^ reg4365)}));
                  for (forvar4534 = (1'h0); (forvar4534 < (1'h1)); forvar4534 = (forvar4534 + (1'h1)))
                    begin
                      reg4535 <= (reg4363 ?
                          $unsigned(({(8'ha4)} ?
                              {reg4430} : forvar4532)) : $signed(reg4331));
                      reg4536 <= forvar4534[(3'h5):(2'h2)];
                      reg4537 <= reg4528;
                      reg4538 <= (~reg4336);
                    end
                  for (forvar4539 = (1'h0); (forvar4539 < (2'h3)); forvar4539 = (forvar4539 + (1'h1)))
                    begin
                      reg4540 <= $signed((reg4351 ?
                          ((reg4360 ? reg4385 : reg4354) ?
                              reg4477[(4'he):(4'hd)] : $signed((8'h9e))) : (!(reg4372 | reg4341))));
                      reg4541 <= (-$signed(reg4427[(2'h3):(1'h0)]));
                    end
                end
              reg4542 <= (^~$signed(((-reg4351) ~^ reg4345[(4'hf):(4'hb)])));
            end
          else
            begin
              for (forvar4528 = (1'h0); (forvar4528 < (1'h0)); forvar4528 = (forvar4528 + (1'h1)))
                begin
                  for (forvar4529 = (1'h0); (forvar4529 < (2'h3)); forvar4529 = (forvar4529 + (1'h1)))
                    begin
                      reg4530 <= reg4529[(4'hb):(4'hb)];
                    end
                end
              reg4531 <= (($signed(reg4530) ?
                  reg4331[(1'h1):(1'h0)] : reg4529) || {$unsigned(reg4433[(2'h3):(2'h2)])});
              if (({((wire3 && reg4452) != $unsigned(reg4505))} ?
                  $signed(($signed(reg4502) ?
                      (reg4517 ?
                          reg4484 : reg4464) : (-(8'ha3)))) : $unsigned($signed(reg4407[(1'h0):(1'h0)]))))
                begin
                  if (reg4407)
                    begin
                      reg4532 <= (reg4482[(1'h1):(1'h1)] ?
                          reg4509[(1'h1):(1'h0)] : (8'hb3));
                    end
                  else
                    begin
                      reg4532 <= (~^reg4351);
                      reg4533 <= (^~(!((reg4385 ? reg4362 : reg4500) ?
                          (8'haa) : reg4510)));
                      reg4534 <= reg4504[(4'h9):(2'h2)];
                    end
                  reg4535 <= $signed($unsigned((!(reg4501 != (8'ha4)))));
                end
              else
                begin
                  for (forvar4532 = (1'h0); (forvar4532 < (1'h0)); forvar4532 = (forvar4532 + (1'h1)))
                    begin
                      reg4533 <= (($unsigned(reg4379[(4'hf):(4'ha)]) > (reg4424[(1'h0):(1'h0)] || (reg4447 ?
                          reg4453 : reg4352))) | $signed($unsigned($signed(wire0))));
                      reg4534 <= $unsigned($unsigned($unsigned((forvar4519 ?
                          (8'ha2) : (8'haf)))));
                      reg4535 <= (reg4353[(4'ha):(2'h2)] << {(reg4380 != reg4356)});
                    end
                  reg4536 <= $unsigned($unsigned($signed(reg4390)));
                  for (forvar4537 = (1'h0); (forvar4537 < (2'h2)); forvar4537 = (forvar4537 + (1'h1)))
                    begin
                      reg4538 <= ($unsigned(reg4468[(2'h2):(1'h0)]) ?
                          reg4439 : (8'hac));
                      reg4539 <= {reg4373};
                    end
                  if (wire4318[(4'hc):(4'h8)])
                    begin
                      reg4540 <= $signed($unsigned({((8'hb0) ^~ reg4356)}));
                      reg4541 <= {(reg4357[(4'he):(4'hb)] && ($unsigned(reg4394) ?
                              wire3 : $signed(reg4399)))};
                      reg4542 <= (~|$unsigned(reg4385[(3'h4):(1'h0)]));
                      reg4543 <= reg4373[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg4540 <= ((reg4464[(1'h0):(1'h0)] > $signed((8'hb2))) >> (~|(8'had)));
                      reg4541 <= wire3;
                      reg4542 <= (^~$unsigned((wire1 ?
                          {reg4496} : (reg4335 ^ reg4346))));
                      reg4543 <= (~&(8'haa));
                    end
                end
              if ($signed((-(reg4343 ? reg4332[(3'h4):(2'h3)] : reg4501))))
                begin
                  reg4544 <= reg4471[(2'h2):(1'h1)];
                  for (forvar4545 = (1'h0); (forvar4545 < (1'h0)); forvar4545 = (forvar4545 + (1'h1)))
                    begin
                      reg4546 <= $unsigned(($signed($unsigned(reg4353)) << reg4370));
                    end
                  if ($unsigned($signed($signed({reg4530}))))
                    begin
                      reg4547 <= {(reg4493 - {reg4436})};
                    end
                  else
                    begin
                      reg4547 <= wire4319[(2'h2):(1'h0)];
                      reg4548 <= $unsigned(($signed(((8'ha5) ?
                              reg4492 : reg4440)) ?
                          reg4362 : ((8'ha4) ~^ $unsigned(reg4468))));
                      reg4549 <= (~(^$unsigned(reg4348[(2'h2):(2'h2)])));
                    end
                end
              else
                begin
                  for (forvar4544 = (1'h0); (forvar4544 < (2'h2)); forvar4544 = (forvar4544 + (1'h1)))
                    begin
                      reg4545 <= $unsigned((((^wire0) << $signed(reg4538)) < $signed($signed(reg4476))));
                      reg4546 <= $signed(((!(^reg4479)) ?
                          (reg4339 <= (reg4502 >> reg4415)) : $signed((wire4518 ?
                              reg4390 : reg4515))));
                    end
                  for (forvar4547 = (1'h0); (forvar4547 < (2'h3)); forvar4547 = (forvar4547 + (1'h1)))
                    begin
                      reg4548 <= ((reg4434[(1'h0):(1'h0)] != ((reg4435 ^~ reg4358) ~^ reg4502[(4'hb):(3'h5)])) >= (($unsigned(reg4509) ?
                          $unsigned(reg4450) : {reg4477}) == reg4356));
                      reg4549 <= reg4384;
                    end
                end
            end
          for (forvar4550 = (1'h0); (forvar4550 < (2'h3)); forvar4550 = (forvar4550 + (1'h1)))
            begin
              if ((reg4322[(1'h0):(1'h0)] | ($signed(reg4423[(3'h7):(2'h3)]) ?
                  $unsigned((reg4482 ? (8'ha7) : (8'hb8))) : (+{reg4476}))))
                begin
                  for (forvar4551 = (1'h0); (forvar4551 < (1'h1)); forvar4551 = (forvar4551 + (1'h1)))
                    begin
                      reg4552 <= {($signed((~^reg4504)) ?
                              $unsigned(((8'hb9) >>> reg4445)) : (~|(reg4469 == reg4433)))};
                      reg4553 <= {$signed({wire0})};
                    end
                end
              else
                begin
                  reg4551 <= reg4539[(1'h0):(1'h0)];
                end
            end
        end
      if (((((reg4415 ? reg4468 : reg4432) ?
              reg4342 : $signed(reg4517)) ^~ {(8'hb5)}) ?
          $signed(reg4331) : $unsigned(((reg4344 >>> reg4334) == (reg4462 ?
              reg4330 : reg4377)))))
        begin
          reg4554 <= $unsigned($signed({reg4494[(3'h5):(2'h3)]}));
          for (forvar4555 = (1'h0); (forvar4555 < (1'h0)); forvar4555 = (forvar4555 + (1'h1)))
            begin
              for (forvar4556 = (1'h0); (forvar4556 < (2'h2)); forvar4556 = (forvar4556 + (1'h1)))
                begin
                  if ($signed($signed((!(^~(8'h9e))))))
                    begin
                      reg4557 <= $signed((~|(reg4553 ?
                          (8'ha7) : (reg4430 <<< reg4507))));
                      reg4558 <= $unsigned(reg4421[(3'h5):(2'h3)]);
                      reg4559 <= $signed($signed(reg4502[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg4557 <= $unsigned((~(reg4356 ?
                          $unsigned(reg4544) : reg4341)));
                    end
                  if ($unsigned(((^reg4401[(2'h2):(1'h0)]) ~^ ((!reg4424) > (reg4461 ?
                      reg4387 : reg4495)))))
                    begin
                      reg4560 <= ($unsigned(reg4450) ?
                          {$signed((~^(8'hae)))} : $signed({$signed(reg4544)}));
                    end
                  else
                    begin
                      reg4560 <= (+$unsigned(($unsigned(reg4535) ?
                          $unsigned(reg4450) : reg4449[(3'h4):(3'h4)])));
                    end
                  reg4561 <= (~|forvar4520);
                  reg4562 <= $signed($unsigned(wire1[(4'hd):(4'hb)]));
                end
              for (forvar4563 = (1'h0); (forvar4563 < (1'h1)); forvar4563 = (forvar4563 + (1'h1)))
                begin
                  if (((reg4480 ?
                      $unsigned(forvar4556) : (~$signed(reg4441))) & $signed({(^(8'ha0))})))
                    begin
                      reg4564 <= $unsigned({((reg4506 ?
                              reg4502 : reg4349) > (^~reg4525))});
                      reg4565 <= (reg4531[(4'hb):(2'h3)] ?
                          wire3[(4'hd):(4'hc)] : $signed((8'ha3)));
                    end
                  else
                    begin
                      reg4564 <= reg4344[(3'h6):(3'h6)];
                      reg4565 <= (|reg4561[(3'h6):(3'h6)]);
                      reg4566 <= ($unsigned(reg4482[(3'h4):(3'h4)]) ?
                          {reg4539} : $signed((reg4538[(3'h4):(1'h1)] << $unsigned(reg4440))));
                    end
                  if ($unsigned((8'hba)))
                    begin
                      reg4567 <= reg4451;
                      reg4568 <= (8'haa);
                      reg4569 <= {reg4530[(3'h6):(1'h0)]};
                    end
                  else
                    begin
                      reg4567 <= $signed(((reg4464 ?
                              $signed((8'haa)) : $signed(reg4423)) ?
                          $signed(reg4473) : $signed(reg4554[(3'h5):(2'h2)])));
                      reg4568 <= (8'hb0);
                    end
                  for (forvar4570 = (1'h0); (forvar4570 < (1'h0)); forvar4570 = (forvar4570 + (1'h1)))
                    begin
                      reg4571 <= (~&{(+{forvar4537})});
                      reg4572 <= (reg4557 ?
                          (reg4560[(3'h6):(1'h1)] ?
                              (reg4467[(2'h2):(2'h2)] ?
                                  ((8'ha8) <= (8'ha6)) : (reg4427 + reg4537)) : ($unsigned((8'hb6)) > reg4375[(4'hf):(3'h4)])) : $signed(wire2[(3'h5):(1'h0)]));
                      reg4573 <= (~$signed($unsigned(reg4564[(1'h1):(1'h0)])));
                    end
                  reg4574 <= reg4344;
                end
              if ($unsigned((~|(~&$unsigned(reg4507)))))
                begin
                  for (forvar4575 = (1'h0); (forvar4575 < (1'h0)); forvar4575 = (forvar4575 + (1'h1)))
                    begin
                      reg4576 <= reg4386[(1'h1):(1'h0)];
                      reg4577 <= ({(reg4446 ?
                              reg4337[(4'ha):(3'h7)] : (!reg4412))} ~^ $unsigned({(&reg4379)}));
                    end
                  reg4578 <= ((~^$unsigned(reg4391[(4'h9):(3'h6)])) ?
                      (((+reg4375) ?
                          (~reg4436) : (|(8'haf))) - ($signed((8'ha3)) ?
                          (reg4355 ?
                              reg4461 : reg4369) : {reg4338})) : $signed($unsigned(reg4571)));
                end
              else
                begin
                  for (forvar4575 = (1'h0); (forvar4575 < (2'h2)); forvar4575 = (forvar4575 + (1'h1)))
                    begin
                      reg4576 <= ($unsigned($unsigned((reg4578 ?
                              reg4560 : reg4354))) ?
                          $unsigned(reg4529[(4'hb):(3'h6)]) : {(&$signed((8'h9c)))});
                      reg4577 <= ($unsigned(reg4436[(4'h8):(3'h4)]) <<< (!(8'had)));
                      reg4578 <= (~^(($unsigned(reg4494) < (reg4465 * reg4527)) | ($unsigned(reg4573) ?
                          reg4578 : reg4473)));
                      reg4579 <= $signed((-{{(8'ha1)}}));
                    end
                  reg4580 <= (reg4363[(2'h3):(1'h1)] ?
                      reg4460 : (($unsigned(reg4349) ?
                          reg4424[(1'h1):(1'h1)] : ((8'h9d) ?
                              forvar4544 : reg4457)) != reg4357));
                end
            end
        end
      else
        begin
          for (forvar4554 = (1'h0); (forvar4554 < (2'h3)); forvar4554 = (forvar4554 + (1'h1)))
            begin
              for (forvar4555 = (1'h0); (forvar4555 < (2'h2)); forvar4555 = (forvar4555 + (1'h1)))
                begin
                  for (forvar4556 = (1'h0); (forvar4556 < (1'h1)); forvar4556 = (forvar4556 + (1'h1)))
                    begin
                      reg4557 <= $unsigned(reg4521);
                      reg4558 <= reg4371;
                    end
                end
              reg4559 <= $unsigned(reg4486[(4'hb):(3'h4)]);
            end
          if ($signed($unsigned($unsigned((+reg4547)))))
            begin
              for (forvar4560 = (1'h0); (forvar4560 < (1'h0)); forvar4560 = (forvar4560 + (1'h1)))
                begin
                  reg4561 <= $signed($unsigned($signed($signed(reg4440))));
                end
            end
          else
            begin
              for (forvar4560 = (1'h0); (forvar4560 < (2'h3)); forvar4560 = (forvar4560 + (1'h1)))
                begin
                  for (forvar4561 = (1'h0); (forvar4561 < (2'h2)); forvar4561 = (forvar4561 + (1'h1)))
                    begin
                      reg4562 <= ($signed($signed(reg4453)) >= ((+(forvar4537 ?
                              reg4538 : reg4380)) ?
                          $signed((reg4493 ?
                              reg4409 : reg4573)) : reg4469[(4'h9):(4'h9)]));
                      reg4563 <= ((^($signed(reg4393) ?
                          $unsigned(reg4375) : (reg4451 ?
                              reg4348 : reg4560))) << reg4387);
                    end
                end
              for (forvar4564 = (1'h0); (forvar4564 < (2'h3)); forvar4564 = (forvar4564 + (1'h1)))
                begin
                  reg4565 <= (^(((8'hba) ?
                      $unsigned((8'ha4)) : reg4435[(1'h0):(1'h0)]) - $signed($unsigned(reg4468))));
                  reg4566 <= $signed((($unsigned(reg4366) ?
                      $signed(reg4481) : $signed(reg4496)) != reg4397));
                  for (forvar4567 = (1'h0); (forvar4567 < (1'h1)); forvar4567 = (forvar4567 + (1'h1)))
                    begin
                      reg4568 <= $unsigned((reg4399 ?
                          ((|reg4487) | $signed(reg4337)) : $unsigned($unsigned(reg4495))));
                      reg4569 <= $signed($unsigned($signed($signed(wire4319))));
                      reg4570 <= $unsigned(((^~(|reg4343)) ?
                          reg4460 : reg4431));
                      reg4571 <= ($signed(((8'hb3) ?
                          {reg4499} : $unsigned(reg4541))) ^ reg4346);
                    end
                end
              for (forvar4572 = (1'h0); (forvar4572 < (2'h3)); forvar4572 = (forvar4572 + (1'h1)))
                begin
                  for (forvar4573 = (1'h0); (forvar4573 < (1'h1)); forvar4573 = (forvar4573 + (1'h1)))
                    begin
                      reg4574 <= reg4332;
                      reg4575 <= reg4507[(3'h6):(2'h2)];
                      reg4576 <= reg4390[(2'h3):(1'h1)];
                      reg4577 <= reg4439[(1'h1):(1'h0)];
                    end
                  if ({$signed(({reg4577} ? (reg4452 & reg4536) : {reg4541}))})
                    begin
                      reg4578 <= $unsigned(($signed({reg4553}) - ((reg4500 ?
                              reg4453 : reg4331) ?
                          reg4379[(2'h2):(2'h2)] : (&(8'hba)))));
                      reg4579 <= {((8'ha7) >= forvar4567)};
                      reg4580 <= ((^~{(reg4540 && reg4413)}) ?
                          $signed((reg4491 ?
                              $signed((8'hb7)) : $unsigned(reg4363))) : (({reg4366} != (reg4465 | reg4352)) >= ($unsigned(reg4479) ?
                              $unsigned(reg4362) : (~|(8'ha7)))));
                      reg4581 <= (reg4543 <= ((reg4431[(2'h2):(1'h0)] ?
                              $unsigned((8'hba)) : reg4552) ?
                          reg4478 : (+reg4339)));
                    end
                  else
                    begin
                      reg4578 <= {((^~(8'hac)) == (^~(8'hb1)))};
                      reg4579 <= (((forvar4532[(2'h3):(2'h2)] ?
                              $signed(reg4398) : (!reg4497)) ^~ ((wire1 & reg4560) && $unsigned(forvar4572))) ?
                          {$signed(((8'hab) << reg4408))} : {({reg4512} ?
                                  ((8'hae) ?
                                      reg4399 : reg4399) : $signed(reg4364))});
                      reg4580 <= ($signed($signed((reg4492 + reg4405))) | {((8'ha5) < {reg4497})});
                    end
                  for (forvar4582 = (1'h0); (forvar4582 < (2'h3)); forvar4582 = (forvar4582 + (1'h1)))
                    begin
                      reg4583 <= (^~{((^reg4516) << $signed(reg4382))});
                    end
                end
            end
        end
      for (forvar4584 = (1'h0); (forvar4584 < (2'h2)); forvar4584 = (forvar4584 + (1'h1)))
        begin
          if (($signed((^reg4355[(4'hc):(1'h0)])) ~^ (~|reg4344)))
            begin
              if (reg4338[(2'h3):(2'h3)])
                begin
                  for (forvar4585 = (1'h0); (forvar4585 < (1'h0)); forvar4585 = (forvar4585 + (1'h1)))
                    begin
                      reg4586 <= (((8'ha5) || (reg4338[(1'h0):(1'h0)] ?
                          (reg4468 ?
                              wire0 : reg4387) : (reg4514 <<< wire3))) == (~forvar4532[(4'h9):(2'h3)]));
                      reg4587 <= (({(reg4477 != reg4393)} ?
                              reg4531 : ((reg4510 << reg4349) ?
                                  reg4497[(2'h3):(2'h2)] : (reg4525 >> (8'hb2)))) ?
                          reg4517[(4'h9):(3'h7)] : $signed((~&(reg4444 ?
                              reg4512 : reg4384))));
                      reg4588 <= $unsigned(($unsigned($unsigned(reg4377)) ?
                          $unsigned(reg4348) : reg4400));
                      reg4589 <= $unsigned((~reg4570));
                    end
                  if (({reg4467[(2'h2):(2'h2)]} + {{$unsigned(reg4483)}}))
                    begin
                      reg4590 <= reg4579[(3'h7):(3'h4)];
                      reg4591 <= reg4464[(1'h0):(1'h0)];
                      reg4592 <= $unsigned((8'h9d));
                    end
                  else
                    begin
                      reg4590 <= reg4573[(1'h1):(1'h1)];
                      reg4591 <= $signed(($unsigned($signed(reg4348)) * (((8'hac) ?
                              forvar4575 : wire4319) ?
                          $signed(reg4500) : $unsigned(reg4527))));
                    end
                  if ($signed(((|(reg4380 ? reg4436 : forvar4575)) ?
                      (|(!reg4506)) : $signed($unsigned(reg4484)))))
                    begin
                      reg4593 <= reg4552[(3'h4):(1'h0)];
                      reg4594 <= reg4504[(4'h8):(3'h6)];
                      reg4595 <= ($signed(($signed(reg4575) ?
                          (forvar4584 ^ reg4440) : {reg4394})) * reg4495);
                    end
                  else
                    begin
                      reg4593 <= reg4533;
                      reg4594 <= ((((~^reg4445) ^ (|reg4571)) <<< (^~$unsigned(reg4464))) ?
                          (-forvar4567[(2'h3):(2'h2)]) : ($signed(forvar4550[(2'h2):(1'h0)]) ?
                              (+reg4455[(3'h5):(1'h0)]) : forvar4564[(1'h0):(1'h0)]));
                      reg4595 <= forvar4520;
                      reg4596 <= $signed($unsigned($unsigned($signed(reg4421))));
                    end
                end
              else
                begin
                  if (($signed((reg4593[(3'h7):(1'h1)] ?
                      forvar4550[(1'h1):(1'h0)] : reg4574[(2'h2):(2'h2)])) >> (~|(~|$unsigned((8'ha8))))))
                    begin
                      reg4585 <= {$unsigned(reg4586[(1'h1):(1'h1)])};
                    end
                  else
                    begin
                      reg4585 <= ((reg4578[(4'hc):(4'h9)] ?
                          reg4514 : reg4449[(3'h5):(1'h0)]) != $signed(forvar4561[(2'h3):(2'h3)]));
                      reg4586 <= (^(($unsigned(reg4571) ?
                              (forvar4519 & reg4383) : forvar4539) ?
                          ((~^(8'ha1)) && (8'hb1)) : reg4540));
                      reg4587 <= (reg4577 << reg4344);
                      reg4588 <= {($unsigned({reg4546}) > $signed($signed(reg4376)))};
                    end
                  for (forvar4589 = (1'h0); (forvar4589 < (2'h3)); forvar4589 = (forvar4589 + (1'h1)))
                    begin
                      reg4590 <= {forvar4545[(1'h1):(1'h1)]};
                      reg4591 <= reg4476[(1'h1):(1'h1)];
                      reg4592 <= ($unsigned(reg4407) ?
                          $unsigned(reg4352[(1'h1):(1'h1)]) : reg4386);
                    end
                end
              if ($signed((!reg4338)))
                begin
                  for (forvar4597 = (1'h0); (forvar4597 < (2'h3)); forvar4597 = (forvar4597 + (1'h1)))
                    begin
                      reg4598 <= $signed((~^({forvar4521} == $signed(reg4432))));
                      reg4599 <= (reg4351 ? reg4360 : reg4548);
                      reg4600 <= (((forvar4537 ? reg4546 : {forvar4547}) ?
                              (^~{(8'hab)}) : ((^~reg4368) ?
                                  $unsigned(reg4376) : (reg4590 ?
                                      reg4548 : reg4327))) ?
                          (8'hae) : (($unsigned(reg4376) == (reg4450 ?
                              reg4509 : reg4380)) << (reg4450[(3'h4):(2'h3)] > reg4524[(4'hc):(3'h7)])));
                    end
                  for (forvar4601 = (1'h0); (forvar4601 < (1'h1)); forvar4601 = (forvar4601 + (1'h1)))
                    begin
                      reg4602 <= {$signed(reg4328)};
                    end
                  for (forvar4603 = (1'h0); (forvar4603 < (2'h2)); forvar4603 = (forvar4603 + (1'h1)))
                    begin
                      reg4604 <= (({forvar4589[(1'h1):(1'h1)]} ?
                              ({reg4368} ?
                                  {(8'ha6)} : (reg4336 >= reg4600)) : reg4592) ?
                          reg4500[(3'h4):(2'h2)] : $signed($unsigned((~&reg4338))));
                    end
                  for (forvar4605 = (1'h0); (forvar4605 < (2'h2)); forvar4605 = (forvar4605 + (1'h1)))
                    begin
                      reg4606 <= {reg4585[(3'h4):(3'h4)]};
                      reg4607 <= reg4409;
                    end
                end
              else
                begin
                  for (forvar4597 = (1'h0); (forvar4597 < (1'h0)); forvar4597 = (forvar4597 + (1'h1)))
                    begin
                      reg4598 <= $unsigned((^~$unsigned($unsigned(reg4522))));
                      reg4599 <= (+(8'hb5));
                      reg4600 <= $signed($signed($signed(reg4390[(1'h0):(1'h0)])));
                    end
                  if (reg4398)
                    begin
                      reg4601 <= (&reg4537[(3'h5):(3'h5)]);
                      reg4602 <= {reg4385[(1'h1):(1'h1)]};
                    end
                  else
                    begin
                      reg4601 <= {$signed(($unsigned(reg4413) * (reg4523 || reg4332)))};
                      reg4602 <= (reg4346 >> $signed({$unsigned(reg4359)}));
                      reg4603 <= {((reg4529[(3'h6):(3'h6)] ?
                              reg4565[(2'h3):(2'h3)] : $signed(reg4351)) == reg4351[(2'h2):(1'h0)])};
                    end
                end
              for (forvar4608 = (1'h0); (forvar4608 < (2'h2)); forvar4608 = (forvar4608 + (1'h1)))
                begin
                  for (forvar4609 = (1'h0); (forvar4609 < (1'h0)); forvar4609 = (forvar4609 + (1'h1)))
                    begin
                      reg4610 <= $unsigned(reg4457);
                      reg4611 <= (&$signed((+$signed(forvar4521))));
                      reg4612 <= (!(~&reg4444));
                    end
                  for (forvar4613 = (1'h0); (forvar4613 < (1'h1)); forvar4613 = (forvar4613 + (1'h1)))
                    begin
                      reg4614 <= (~&$unsigned(((reg4539 << forvar4554) ?
                          $signed(reg4478) : (8'hb2))));
                      reg4615 <= {reg4489};
                      reg4616 <= $unsigned({$unsigned(reg4548[(1'h1):(1'h0)])});
                    end
                end
              for (forvar4617 = (1'h0); (forvar4617 < (1'h1)); forvar4617 = (forvar4617 + (1'h1)))
                begin
                  reg4618 <= (^$unsigned((~|(forvar4584 || forvar4534))));
                end
            end
          else
            begin
              reg4585 <= reg4415[(4'ha):(3'h6)];
              if ($signed((+reg4351[(3'h4):(1'h1)])))
                begin
                  reg4586 <= reg4445;
                  if (reg4372[(3'h5):(2'h3)])
                    begin
                      reg4587 <= ($signed((8'hb0)) ?
                          $unsigned(((+(8'hb6)) & $unsigned(reg4522))) : {$unsigned((reg4547 < reg4422))});
                      reg4588 <= forvar4609;
                      reg4589 <= (((+(reg4387 != reg4338)) ?
                              forvar4563[(3'h5):(3'h4)] : reg4353[(3'h4):(2'h2)]) ?
                          {reg4547} : wire4319);
                    end
                  else
                    begin
                      reg4587 <= (($unsigned($unsigned(reg4449)) ?
                          ((~&reg4398) ?
                              (reg4579 <<< reg4612) : forvar4605) : reg4379) - reg4576);
                      reg4588 <= (+(~^{$unsigned((8'h9d))}));
                      reg4589 <= {reg4387[(1'h0):(1'h0)]};
                      reg4590 <= $unsigned((~&reg4380[(4'h8):(2'h3)]));
                    end
                  if ((~^$signed((!(forvar4585 ? reg4523 : reg4601)))))
                    begin
                      reg4591 <= reg4424;
                      reg4592 <= ($unsigned(((reg4551 >= (8'hb0)) ?
                              (wire1 >= (8'haf)) : wire4320[(4'h8):(2'h2)])) ?
                          reg4492[(3'h4):(1'h0)] : ($signed($signed(forvar4601)) * (~|$signed(reg4370))));
                    end
                  else
                    begin
                      reg4591 <= $signed($signed($unsigned(((8'haf) == reg4445))));
                      reg4592 <= reg4433;
                      reg4593 <= (!$unsigned((&(|reg4483))));
                      reg4594 <= $unsigned({((reg4592 || forvar4555) ?
                              (reg4355 ~^ wire0) : (~(8'ha2)))});
                    end
                  if ((8'ha8))
                    begin
                      reg4595 <= $unsigned($unsigned((((8'hb0) << reg4333) ^~ (reg4474 >= reg4433))));
                      reg4596 <= forvar4601[(4'h8):(3'h6)];
                      reg4597 <= (~&wire4518);
                      reg4598 <= reg4444[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg4595 <= (|$signed($unsigned((reg4562 ?
                          reg4513 : (8'ha1)))));
                      reg4596 <= ((forvar4520[(3'h7):(3'h7)] ?
                              $signed($signed(reg4339)) : (-(|reg4509))) ?
                          (!reg4499[(2'h2):(1'h0)]) : reg4357[(4'hf):(2'h3)]);
                      reg4597 <= (reg4381[(3'h5):(1'h1)] ?
                          reg4601 : $unsigned(((8'hb9) << $signed(wire4316))));
                      reg4598 <= $unsigned((forvar4534[(3'h7):(3'h6)] || ($unsigned(forvar4544) ?
                          (reg4574 | forvar4572) : $signed(reg4377))));
                    end
                end
              else
                begin
                  if ($unsigned(reg4548[(4'hf):(2'h3)]))
                    begin
                      reg4586 <= (reg4533[(1'h1):(1'h0)] ?
                          reg4327[(2'h2):(2'h2)] : $unsigned(reg4588));
                      reg4587 <= reg4542[(1'h0):(1'h0)];
                      reg4588 <= (((^$unsigned(reg4587)) ?
                          $signed(((8'hb1) <<< reg4340)) : ($unsigned(reg4372) || {reg4338})) <<< $signed($unsigned(reg4445[(1'h1):(1'h0)])));
                      reg4589 <= $unsigned($signed((+$signed(forvar4570))));
                    end
                  else
                    begin
                      reg4586 <= (8'hba);
                      reg4587 <= $signed(((|(reg4532 ? (8'ha3) : (8'ha9))) ?
                          ($unsigned(reg4383) ?
                              $unsigned(reg4510) : (&forvar4572)) : (reg4603[(3'h7):(2'h3)] < reg4597[(1'h1):(1'h1)])));
                      reg4588 <= (-({$unsigned(reg4562)} - reg4599));
                    end
                end
              for (forvar4599 = (1'h0); (forvar4599 < (2'h2)); forvar4599 = (forvar4599 + (1'h1)))
                begin
                  if ($unsigned((($signed(reg4553) ?
                          $signed(reg4334) : (+(8'hba))) ?
                      reg4561[(4'hd):(4'hc)] : reg4524[(4'hd):(3'h7)])))
                    begin
                      reg4600 <= (!forvar4551[(3'h6):(3'h6)]);
                    end
                  else
                    begin
                      reg4600 <= ((reg4430 ^ $signed({reg4348})) ?
                          $signed(reg4585) : reg4360[(3'h5):(2'h3)]);
                      reg4601 <= ($unsigned(($signed(reg4540) ^~ reg4408[(2'h2):(2'h2)])) < $signed(reg4534[(2'h3):(1'h0)]));
                      reg4602 <= $signed({(reg4464 - forvar4545[(1'h1):(1'h1)])});
                    end
                  if ((|(((~^(8'hb8)) ~^ (+reg4612)) - reg4527)))
                    begin
                      reg4603 <= $signed($unsigned((&reg4411)));
                    end
                  else
                    begin
                      reg4603 <= ((^~($signed(reg4592) ?
                              $signed(reg4581) : $signed(reg4340))) ?
                          (|$unsigned((~^forvar4561))) : forvar4573[(1'h0):(1'h0)]);
                    end
                  for (forvar4604 = (1'h0); (forvar4604 < (1'h0)); forvar4604 = (forvar4604 + (1'h1)))
                    begin
                      reg4605 <= reg4377;
                      reg4606 <= ({$unsigned(forvar4575[(2'h2):(1'h1)])} >>> (8'ha3));
                      reg4607 <= reg4419[(2'h3):(2'h3)];
                      reg4608 <= $unsigned(reg4441[(1'h0):(1'h0)]);
                    end
                  for (forvar4609 = (1'h0); (forvar4609 < (2'h3)); forvar4609 = (forvar4609 + (1'h1)))
                    begin
                      reg4610 <= {{(^~(wire2 ? forvar4561 : (8'h9c)))}};
                      reg4611 <= $unsigned(reg4385[(3'h4):(2'h2)]);
                      reg4612 <= (~^(({wire3} * $signed(wire3)) & ((^~reg4474) ?
                          forvar4519[(3'h7):(1'h0)] : (reg4541 ?
                              (8'h9f) : reg4463))));
                      reg4613 <= reg4327[(1'h0):(1'h0)];
                    end
                end
              reg4614 <= (forvar4613 ~^ {$unsigned((reg4493 ?
                      reg4603 : reg4365))});
            end
        end
      for (forvar4619 = (1'h0); (forvar4619 < (1'h0)); forvar4619 = (forvar4619 + (1'h1)))
        begin
          if ($signed((reg4364 ?
              ((reg4346 ? (8'haa) : reg4604) ?
                  $signed(reg4430) : (reg4446 >= reg4493)) : ($signed(reg4363) ?
                  reg4462 : reg4563))))
            begin
              if (reg4327)
                begin
                  if (forvar4532)
                    begin
                      reg4620 <= {((+(!reg4344)) ?
                              reg4497[(2'h3):(2'h2)] : (reg4566[(1'h0):(1'h0)] ?
                                  reg4598 : {reg4345}))};
                      reg4621 <= (~(((reg4331 && reg4533) || reg4615[(2'h3):(2'h2)]) >> {{reg4489}}));
                    end
                  else
                    begin
                      reg4620 <= reg4501;
                      reg4621 <= (reg4507[(1'h0):(1'h0)] ^~ $signed(((reg4349 ^~ reg4553) < $unsigned(reg4347))));
                      reg4622 <= $unsigned({(reg4393 ?
                              (reg4354 ?
                                  reg4521 : reg4494) : (reg4355 * forvar4589))});
                    end
                  for (forvar4623 = (1'h0); (forvar4623 < (2'h2)); forvar4623 = (forvar4623 + (1'h1)))
                    begin
                      reg4624 <= ($unsigned($unsigned((~&(8'hb5)))) * reg4586);
                      reg4625 <= forvar4604[(4'hb):(1'h1)];
                    end
                  for (forvar4626 = (1'h0); (forvar4626 < (1'h0)); forvar4626 = (forvar4626 + (1'h1)))
                    begin
                      reg4627 <= ((($unsigned(reg4333) ?
                          (forvar4526 ?
                              reg4341 : reg4389) : $signed(forvar4551)) << {$unsigned(reg4615)}) >>> {reg4624[(2'h2):(1'h0)]});
                      reg4628 <= $signed($unsigned((~^(|reg4563))));
                      reg4629 <= {{(~^((8'ha3) ? reg4380 : forvar4534))}};
                      reg4630 <= reg4338[(4'ha):(4'ha)];
                    end
                end
              else
                begin
                  for (forvar4620 = (1'h0); (forvar4620 < (1'h0)); forvar4620 = (forvar4620 + (1'h1)))
                    begin
                      reg4621 <= $signed(((reg4439 + $unsigned(reg4567)) >>> reg4601));
                      reg4622 <= (-{$unsigned(forvar4599)});
                      reg4623 <= (|(8'h9e));
                      reg4624 <= forvar4564;
                    end
                  for (forvar4625 = (1'h0); (forvar4625 < (1'h1)); forvar4625 = (forvar4625 + (1'h1)))
                    begin
                      reg4626 <= reg4468[(1'h0):(1'h0)];
                      reg4627 <= (-reg4397);
                      reg4628 <= reg4512[(2'h3):(1'h0)];
                      reg4629 <= reg4328[(2'h2):(1'h0)];
                    end
                  for (forvar4630 = (1'h0); (forvar4630 < (1'h1)); forvar4630 = (forvar4630 + (1'h1)))
                    begin
                      reg4631 <= ({$unsigned(reg4449)} >> (reg4585 << (8'hba)));
                    end
                  for (forvar4632 = (1'h0); (forvar4632 < (2'h2)); forvar4632 = (forvar4632 + (1'h1)))
                    begin
                      reg4633 <= (^~$signed(reg4630[(3'h7):(3'h7)]));
                      reg4634 <= $signed((~|reg4620));
                      reg4635 <= ((~$unsigned($signed(reg4613))) ?
                          (~^{reg4580[(2'h3):(2'h2)]}) : (^~((reg4339 <= reg4620) ?
                              {reg4344} : (^(8'hb8)))));
                    end
                end
              for (forvar4636 = (1'h0); (forvar4636 < (2'h3)); forvar4636 = (forvar4636 + (1'h1)))
                begin
                  reg4637 <= reg4601;
                  reg4638 <= reg4354;
                end
            end
          else
            begin
              for (forvar4620 = (1'h0); (forvar4620 < (2'h2)); forvar4620 = (forvar4620 + (1'h1)))
                begin
                  for (forvar4621 = (1'h0); (forvar4621 < (1'h1)); forvar4621 = (forvar4621 + (1'h1)))
                    begin
                      reg4622 <= forvar4609[(3'h7):(2'h2)];
                      reg4623 <= reg4408[(1'h1):(1'h0)];
                      reg4624 <= ((reg4616 ?
                              (^(reg4487 ?
                                  reg4525 : reg4585)) : $unsigned(reg4347[(4'h8):(1'h1)])) ?
                          $signed($unsigned($signed(forvar4605))) : $unsigned((+{reg4381})));
                    end
                  reg4625 <= reg4469;
                end
              for (forvar4626 = (1'h0); (forvar4626 < (2'h3)); forvar4626 = (forvar4626 + (1'h1)))
                begin
                  reg4627 <= $unsigned((~^(|$unsigned(reg4446))));
                  if ({(~((8'h9e) << (forvar4589 ? reg4535 : forvar4617)))})
                    begin
                      reg4628 <= ({((-reg4589) << $signed(reg4445))} ?
                          $unsigned($signed(reg4533[(3'h4):(2'h3)])) : ((^$unsigned(forvar4556)) ?
                              $unsigned(reg4596[(2'h2):(1'h0)]) : $unsigned($signed(forvar4551))));
                      reg4629 <= reg4404[(3'h4):(3'h4)];
                      reg4630 <= {{(^~(forvar4609 ? reg4570 : (8'hae)))}};
                      reg4631 <= reg4440[(3'h5):(1'h0)];
                    end
                  else
                    begin
                      reg4628 <= (^~$signed(reg4566[(1'h1):(1'h0)]));
                      reg4629 <= ({forvar4603[(3'h7):(3'h4)]} ?
                          (|($unsigned(reg4552) << reg4494)) : $unsigned($unsigned((reg4504 ?
                              reg4338 : (8'hb4)))));
                      reg4630 <= $unsigned((~((~reg4350) ?
                          (reg4565 ? forvar4534 : reg4565) : forvar4534)));
                      reg4631 <= forvar4601;
                    end
                  for (forvar4632 = (1'h0); (forvar4632 < (1'h0)); forvar4632 = (forvar4632 + (1'h1)))
                    begin
                      reg4633 <= (~&(~^(+reg4375[(2'h3):(2'h3)])));
                    end
                end
              reg4634 <= (^$signed({(reg4394 * reg4346)}));
            end
          for (forvar4639 = (1'h0); (forvar4639 < (1'h1)); forvar4639 = (forvar4639 + (1'h1)))
            begin
              reg4640 <= $signed($signed(reg4505));
              for (forvar4641 = (1'h0); (forvar4641 < (2'h3)); forvar4641 = (forvar4641 + (1'h1)))
                begin
                  for (forvar4642 = (1'h0); (forvar4642 < (2'h3)); forvar4642 = (forvar4642 + (1'h1)))
                    begin
                      reg4643 <= reg4616[(4'hc):(4'hc)];
                      reg4644 <= (~|reg4485[(4'hc):(3'h4)]);
                      reg4645 <= (($unsigned($signed((8'h9c))) >> (8'hb8)) < {$signed((~|reg4504))});
                    end
                  for (forvar4646 = (1'h0); (forvar4646 < (2'h2)); forvar4646 = (forvar4646 + (1'h1)))
                    begin
                      reg4647 <= (reg4604 << $signed(((|(8'hb3)) >>> $signed(forvar4646))));
                      reg4648 <= ($signed(reg4335[(4'ha):(3'h4)]) ?
                          reg4586 : $signed((forvar4636[(4'h9):(3'h7)] ?
                              ((8'ha5) == reg4638) : (reg4453 | reg4331))));
                      reg4649 <= reg4378[(3'h4):(1'h1)];
                    end
                  if ((((^((8'h9d) ?
                      reg4514 : reg4435)) >= (reg4351[(1'h1):(1'h1)] ?
                      reg4434[(2'h3):(2'h2)] : {reg4638})) - ((!(8'ha2)) & $signed($unsigned(reg4623)))))
                    begin
                      reg4650 <= {(^((reg4430 ^~ forvar4589) == $signed(reg4586)))};
                      reg4651 <= (forvar4601 ?
                          (($unsigned(forvar4550) ?
                                  reg4542[(2'h3):(1'h1)] : (forvar4575 == (8'hb9))) ?
                              $signed(reg4635[(2'h3):(1'h1)]) : ($signed(reg4511) > (~&(8'hb7)))) : $unsigned((!(reg4468 ?
                              reg4497 : reg4465))));
                      reg4652 <= {$signed($signed($unsigned(reg4524)))};
                    end
                  else
                    begin
                      reg4650 <= forvar4550[(2'h3):(1'h0)];
                      reg4651 <= ($signed(reg4651) == {((~reg4610) >> (~|reg4552))});
                    end
                  for (forvar4653 = (1'h0); (forvar4653 < (1'h0)); forvar4653 = (forvar4653 + (1'h1)))
                    begin
                      reg4654 <= (8'ha3);
                      reg4655 <= ($unsigned({(reg4445 ?
                              reg4472 : reg4407)}) ~^ reg4631);
                      reg4656 <= $unsigned((~^$unsigned($signed(reg4568))));
                      reg4657 <= reg4597[(1'h0):(1'h0)];
                    end
                end
              for (forvar4658 = (1'h0); (forvar4658 < (1'h0)); forvar4658 = (forvar4658 + (1'h1)))
                begin
                  reg4659 <= (reg4378 ^~ ((|{reg4649}) & (-reg4607)));
                end
            end
        end
    end
  assign wire4660 = ($signed(reg4574[(2'h3):(2'h3)]) ?
                        reg4537 : {((reg4409 ? reg4656 : reg4515) ?
                                reg4450[(1'h1):(1'h1)] : (reg4365 ?
                                    reg4340 : reg4423))});
  assign wire4661 = reg4592[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      if ((reg4593 ? reg4338[(1'h0):(1'h0)] : (8'ha6)))
        begin
          for (forvar4662 = (1'h0); (forvar4662 < (2'h3)); forvar4662 = (forvar4662 + (1'h1)))
            begin
              if (((reg4399 ?
                  ((^reg4581) ?
                      reg4598 : (reg4450 != reg4624)) : reg4647) <<< $signed($unsigned((wire4316 >>> reg4422)))))
                begin
                  for (forvar4663 = (1'h0); (forvar4663 < (1'h1)); forvar4663 = (forvar4663 + (1'h1)))
                    begin
                      reg4664 <= $signed($unsigned($unsigned((reg4492 - reg4342))));
                    end
                  reg4665 <= {reg4542};
                  if (((~|$unsigned($signed(reg4363))) << {(!$unsigned(reg4625))}))
                    begin
                      reg4666 <= reg4551[(1'h0):(1'h0)];
                      reg4667 <= $unsigned((~|(&$unsigned(reg4612))));
                    end
                  else
                    begin
                      reg4666 <= $unsigned(($unsigned($signed(reg4335)) ?
                          (8'ha1) : reg4337));
                      reg4667 <= {((&(reg4375 ?
                              reg4388 : reg4513)) > (&(wire0 < reg4552)))};
                      reg4668 <= reg4616[(3'h7):(3'h7)];
                    end
                end
              else
                begin
                  for (forvar4663 = (1'h0); (forvar4663 < (1'h0)); forvar4663 = (forvar4663 + (1'h1)))
                    begin
                      reg4664 <= $signed(reg4388);
                      reg4665 <= ($signed(reg4538) + (~|reg4574[(1'h0):(1'h0)]));
                    end
                  reg4666 <= (^~$signed({(8'hb9)}));
                end
            end
          reg4669 <= ($unsigned(reg4605) << (^~(8'hb1)));
          for (forvar4670 = (1'h0); (forvar4670 < (2'h2)); forvar4670 = (forvar4670 + (1'h1)))
            begin
              for (forvar4671 = (1'h0); (forvar4671 < (2'h3)); forvar4671 = (forvar4671 + (1'h1)))
                begin
                  reg4672 <= reg4543;
                  reg4673 <= reg4327;
                  reg4674 <= $signed({($signed(reg4457) && reg4547[(4'hb):(3'h6)])});
                end
              for (forvar4675 = (1'h0); (forvar4675 < (1'h1)); forvar4675 = (forvar4675 + (1'h1)))
                begin
                  for (forvar4676 = (1'h0); (forvar4676 < (2'h3)); forvar4676 = (forvar4676 + (1'h1)))
                    begin
                      reg4677 <= reg4596;
                    end
                end
            end
        end
      else
        begin
          if ((reg4471 ? reg4348 : reg4432))
            begin
              reg4662 <= reg4626[(3'h4):(1'h1)];
              if ($signed($unsigned(reg4398)))
                begin
                  reg4663 <= (+reg4534[(1'h1):(1'h0)]);
                  for (forvar4664 = (1'h0); (forvar4664 < (2'h2)); forvar4664 = (forvar4664 + (1'h1)))
                    begin
                      reg4665 <= $signed((^(8'ha5)));
                      reg4666 <= reg4493[(1'h0):(1'h0)];
                      reg4667 <= $unsigned((reg4469[(3'h6):(1'h0)] ?
                          (reg4343 ~^ (8'ha2)) : (8'haa)));
                    end
                  reg4668 <= ((reg4363 < reg4651[(3'h5):(2'h3)]) ?
                      ((~&(reg4348 & reg4344)) <<< (+reg4463)) : $unsigned(reg4495[(3'h6):(1'h0)]));
                  if (($signed(((reg4543 ^ (8'hac)) ?
                          (-reg4497) : ((8'ha4) ? reg4551 : reg4529))) ?
                      (~|$signed((reg4450 <= reg4563))) : reg4614))
                    begin
                      reg4669 <= (((-(-reg4340)) ?
                              reg4471 : ((reg4349 ^ reg4667) ?
                                  (reg4623 ?
                                      reg4414 : reg4475) : (~|reg4375))) ?
                          $signed((^~(|reg4604))) : reg4615[(3'h4):(2'h3)]);
                      reg4670 <= (reg4407 == reg4489[(3'h6):(3'h4)]);
                      reg4671 <= ({$signed(((8'hb7) ? reg4607 : reg4662))} ?
                          (8'ha1) : ((~&reg4378) & reg4674[(1'h1):(1'h1)]));
                      reg4672 <= $signed((reg4379[(4'h8):(2'h3)] ?
                          $unsigned($signed(reg4469)) : reg4486));
                    end
                  else
                    begin
                      reg4669 <= $unsigned($unsigned((reg4369 ?
                          {forvar4662} : ((8'hb9) ? (8'hba) : (8'ha1)))));
                      reg4670 <= reg4557;
                      reg4671 <= $unsigned($signed(((reg4677 ?
                              reg4674 : reg4628) ?
                          {(8'hb1)} : (reg4427 ? reg4514 : (8'hb3)))));
                    end
                end
              else
                begin
                  if ({reg4527[(2'h3):(1'h1)]})
                    begin
                      reg4663 <= $unsigned($unsigned(((8'hb8) ?
                          (&reg4387) : (^wire1))));
                      reg4664 <= ({reg4541} + {(reg4537[(4'h8):(2'h2)] ?
                              $signed(reg4562) : $unsigned(reg4522))});
                    end
                  else
                    begin
                      reg4663 <= ($signed($signed((reg4451 ?
                              reg4381 : (8'ha2)))) ?
                          (-((reg4356 != reg4517) ?
                              (~^(8'hae)) : reg4599)) : (8'hab));
                    end
                  if (reg4393[(4'hd):(3'h7)])
                    begin
                      reg4665 <= (reg4355[(3'h4):(1'h0)] << reg4517);
                      reg4666 <= $unsigned($unsigned(reg4333[(2'h2):(1'h1)]));
                      reg4667 <= (reg4324[(3'h4):(3'h4)] << {(reg4626 ?
                              $unsigned(reg4435) : (reg4384 ?
                                  wire4316 : reg4607))});
                      reg4668 <= reg4474[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg4665 <= (~|reg4347[(4'hc):(3'h5)]);
                      reg4666 <= $signed(reg4409);
                      reg4667 <= $signed({(+(reg4341 ? reg4631 : reg4380))});
                      reg4668 <= {reg4482[(1'h1):(1'h0)]};
                    end
                  if ($signed({(reg4545 ~^ $signed(reg4553))}))
                    begin
                      reg4669 <= {({reg4509[(3'h4):(1'h0)]} & ((reg4559 >> reg4638) * $unsigned(reg4350)))};
                      reg4670 <= reg4605;
                      reg4671 <= reg4357;
                      reg4672 <= (reg4401 ?
                          $signed(reg4336) : reg4407[(4'hc):(4'ha)]);
                    end
                  else
                    begin
                      reg4669 <= reg4668;
                      reg4670 <= ((((reg4506 ? reg4628 : reg4387) ?
                              $signed(reg4599) : (reg4525 << reg4669)) >>> (reg4322[(3'h5):(1'h1)] ?
                              reg4648 : (reg4341 ? (8'hb9) : (8'hb8)))) ?
                          (-$signed(reg4597[(1'h1):(1'h0)])) : reg4324[(1'h0):(1'h0)]);
                    end
                end
              for (forvar4673 = (1'h0); (forvar4673 < (2'h2)); forvar4673 = (forvar4673 + (1'h1)))
                begin
                  if (($unsigned(((reg4366 >> reg4605) ?
                      reg4522[(1'h0):(1'h0)] : $unsigned(reg4449))) * reg4606))
                    begin
                      reg4674 <= $unsigned(({$unsigned(reg4572)} << reg4462[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg4674 <= ($signed(reg4350[(1'h0):(1'h0)]) == reg4563[(2'h3):(1'h0)]);
                    end
                end
              if ($signed($unsigned(((reg4607 | reg4506) - (reg4328 ?
                  reg4589 : reg4474)))))
                begin
                  for (forvar4675 = (1'h0); (forvar4675 < (2'h3)); forvar4675 = (forvar4675 + (1'h1)))
                    begin
                      reg4676 <= ((reg4635 + reg4421[(2'h3):(1'h0)]) < (reg4541[(4'hd):(4'hd)] != reg4340));
                      reg4677 <= ({(reg4455[(1'h0):(1'h0)] ~^ (-reg4480))} >> reg4568[(3'h7):(2'h3)]);
                      reg4678 <= ((+$unsigned((reg4426 >= reg4398))) ?
                          ((~&(reg4461 >= reg4379)) ?
                              $unsigned(reg4437) : reg4651[(4'h9):(1'h1)]) : (!((~^(8'ha8)) ?
                              $unsigned(reg4400) : reg4559[(1'h0):(1'h0)])));
                      reg4679 <= wire4318;
                    end
                  for (forvar4680 = (1'h0); (forvar4680 < (1'h1)); forvar4680 = (forvar4680 + (1'h1)))
                    begin
                      reg4681 <= (~|$signed(((reg4372 ? (8'hb2) : (8'hb9)) ?
                          $unsigned(reg4533) : $signed(reg4467))));
                      reg4682 <= ($signed($signed((8'had))) ?
                          (~|$unsigned($signed(reg4357))) : (({(8'hb3)} >= $unsigned(reg4439)) ?
                              (8'ha2) : $unsigned(reg4391)));
                      reg4683 <= ($signed(reg4512[(2'h3):(1'h0)]) > ($unsigned(reg4626) ?
                          reg4338[(3'h7):(1'h1)] : ($unsigned(reg4585) == reg4679[(3'h6):(3'h6)])));
                      reg4684 <= ((($unsigned((8'hba)) >> reg4395) ^ $signed({reg4422})) ?
                          reg4517 : (^$unsigned(reg4579)));
                    end
                  if ((reg4571[(4'ha):(3'h5)] ?
                      $unsigned(((~|reg4598) ?
                          reg4408[(1'h1):(1'h1)] : $unsigned(reg4506))) : reg4606))
                    begin
                      reg4685 <= ((($unsigned(reg4580) << (reg4430 == reg4468)) ?
                          (-wire4320) : $unsigned($unsigned(reg4387))) >= (~|(^~$unsigned(reg4395))));
                      reg4686 <= (reg4578 >= reg4369[(1'h1):(1'h0)]);
                      reg4687 <= (($signed($unsigned((8'had))) ?
                          $signed((reg4430 ?
                              reg4599 : reg4657)) : reg4554[(3'h5):(2'h2)]) - $unsigned(reg4457[(3'h4):(3'h4)]));
                    end
                  else
                    begin
                      reg4685 <= reg4523[(2'h2):(2'h2)];
                      reg4686 <= (reg4338[(4'ha):(3'h5)] | ($signed(reg4447[(3'h4):(2'h3)]) > {reg4566}));
                      reg4687 <= reg4500[(1'h0):(1'h0)];
                    end
                  for (forvar4688 = (1'h0); (forvar4688 < (1'h0)); forvar4688 = (forvar4688 + (1'h1)))
                    begin
                      reg4689 <= (~(reg4487 ?
                          ($signed(reg4628) ?
                              reg4343[(1'h0):(1'h0)] : $signed(reg4561)) : (-reg4553)));
                      reg4690 <= reg4621;
                      reg4691 <= $unsigned(reg4643);
                    end
                end
              else
                begin
                  for (forvar4675 = (1'h0); (forvar4675 < (1'h1)); forvar4675 = (forvar4675 + (1'h1)))
                    begin
                      reg4676 <= reg4373;
                    end
                  if (((reg4494 ?
                          $signed(reg4624[(4'hd):(4'h8)]) : $signed({reg4571})) ?
                      (8'ha2) : $unsigned((8'hab))))
                    begin
                      reg4677 <= $unsigned((^~({forvar4662} == (reg4473 * reg4585))));
                      reg4678 <= (reg4506[(2'h3):(2'h2)] ?
                          ($unsigned(reg4455[(2'h2):(2'h2)]) ?
                              {(reg4603 ?
                                      reg4546 : reg4334)} : ({reg4497} * (~|reg4407))) : ($signed((8'ha4)) - (~|(reg4354 - (8'hb0)))));
                      reg4679 <= $unsigned((((~&reg4596) | reg4673[(2'h2):(1'h1)]) != (+(~&reg4626))));
                      reg4680 <= (reg4349 ?
                          ($unsigned($unsigned((8'hb3))) ?
                              $signed((reg4346 ?
                                  reg4506 : reg4650)) : $unsigned($unsigned(reg4444))) : ((~reg4371) != (reg4624[(4'ha):(4'h8)] * (reg4371 ?
                              (8'hba) : reg4441))));
                    end
                  else
                    begin
                      reg4677 <= reg4322[(1'h1):(1'h0)];
                      reg4678 <= $signed((reg4463 | $signed((reg4640 > reg4601))));
                      reg4679 <= reg4384;
                    end
                  if (((reg4667[(2'h2):(1'h1)] != reg4685) >>> $unsigned(reg4687)))
                    begin
                      reg4681 <= reg4506[(3'h4):(1'h0)];
                      reg4682 <= $signed(reg4379);
                    end
                  else
                    begin
                      reg4681 <= $unsigned($signed(reg4559));
                      reg4682 <= $unsigned((reg4491[(2'h2):(2'h2)] ?
                          (~reg4475[(3'h4):(3'h4)]) : ((8'ha3) ?
                              ((8'ha3) ? (8'ha4) : reg4354) : (~reg4548))));
                    end
                end
            end
          else
            begin
              for (forvar4662 = (1'h0); (forvar4662 < (1'h0)); forvar4662 = (forvar4662 + (1'h1)))
                begin
                  reg4663 <= ($signed((!wire4319)) ^ $signed(({(8'ha6)} ?
                      (reg4522 | reg4531) : reg4336)));
                  for (forvar4664 = (1'h0); (forvar4664 < (1'h1)); forvar4664 = (forvar4664 + (1'h1)))
                    begin
                      reg4665 <= (({reg4473} >> (^reg4638)) & (((~&reg4501) ?
                          reg4676 : $unsigned((8'haf))) || ($signed(reg4665) ^ reg4348[(4'h8):(3'h5)])));
                      reg4666 <= reg4327[(1'h0):(1'h0)];
                      reg4667 <= (reg4411 || {((reg4670 ^~ reg4682) || $unsigned(reg4523))});
                    end
                  if ((-((~&$signed(reg4689)) ?
                      ((reg4324 >= reg4536) ?
                          wire4661 : ((8'h9d) ^~ reg4481)) : reg4531[(4'h8):(3'h6)])))
                    begin
                      reg4668 <= {reg4415[(4'hb):(4'h9)]};
                      reg4669 <= $signed(reg4500);
                      reg4670 <= {(+($unsigned(reg4383) ?
                              $unsigned(reg4336) : reg4387))};
                      reg4671 <= reg4478[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg4668 <= (8'hac);
                    end
                end
              for (forvar4672 = (1'h0); (forvar4672 < (2'h3)); forvar4672 = (forvar4672 + (1'h1)))
                begin
                  for (forvar4673 = (1'h0); (forvar4673 < (2'h2)); forvar4673 = (forvar4673 + (1'h1)))
                    begin
                      reg4674 <= (&(~^reg4383[(2'h2):(2'h2)]));
                      reg4675 <= (8'ha8);
                      reg4676 <= (~(($signed(reg4453) * $signed(reg4515)) ?
                          reg4497[(2'h3):(2'h2)] : {(~&(8'had))}));
                      reg4677 <= ((reg4656 ?
                              (^$signed(reg4537)) : {reg4669[(3'h5):(1'h1)]}) ?
                          (~^$signed(((8'hb0) ?
                              reg4574 : reg4663))) : reg4592[(1'h0):(1'h0)]);
                    end
                  reg4678 <= $signed((^~forvar4675[(2'h3):(2'h2)]));
                end
              if (reg4578)
                begin
                  if ($unsigned($unsigned(reg4562[(3'h4):(1'h0)])))
                    begin
                      reg4679 <= $signed(($unsigned(reg4605) ^ (reg4592 ?
                          reg4564 : (8'ha2))));
                      reg4680 <= $signed(reg4397);
                      reg4681 <= wire2[(4'h9):(4'h9)];
                    end
                  else
                    begin
                      reg4679 <= $signed({reg4681});
                      reg4680 <= ((-reg4560[(3'h4):(3'h4)]) | (8'hb8));
                      reg4681 <= reg4386;
                    end
                  reg4682 <= $signed(reg4373[(3'h4):(2'h3)]);
                  for (forvar4683 = (1'h0); (forvar4683 < (2'h3)); forvar4683 = (forvar4683 + (1'h1)))
                    begin
                      reg4684 <= reg4464;
                      reg4685 <= $signed({($unsigned(reg4499) ?
                              (^~reg4355) : $signed(reg4534))});
                    end
                  for (forvar4686 = (1'h0); (forvar4686 < (1'h0)); forvar4686 = (forvar4686 + (1'h1)))
                    begin
                      reg4687 <= ((~|$signed(((8'h9c) < reg4439))) >>> (~&reg4481));
                      reg4688 <= reg4610;
                      reg4689 <= {forvar4673[(2'h3):(1'h1)]};
                    end
                end
              else
                begin
                  for (forvar4679 = (1'h0); (forvar4679 < (2'h3)); forvar4679 = (forvar4679 + (1'h1)))
                    begin
                      reg4680 <= reg4474;
                      reg4681 <= (~&reg4553);
                    end
                end
              if ((|{$unsigned($signed(reg4444))}))
                begin
                  for (forvar4690 = (1'h0); (forvar4690 < (2'h3)); forvar4690 = (forvar4690 + (1'h1)))
                    begin
                      reg4691 <= {($signed($unsigned(reg4685)) * (^~reg4570))};
                      reg4692 <= (-(~|forvar4680));
                    end
                  reg4693 <= ((^~reg4668) ?
                      $unsigned(reg4415[(3'h7):(3'h6)]) : reg4495);
                end
              else
                begin
                  for (forvar4690 = (1'h0); (forvar4690 < (2'h2)); forvar4690 = (forvar4690 + (1'h1)))
                    begin
                      reg4691 <= $signed((~reg4412[(3'h4):(1'h0)]));
                      reg4692 <= (reg4324 >>> (&$unsigned({reg4365})));
                    end
                  if (reg4543[(2'h3):(1'h0)])
                    begin
                      reg4693 <= (reg4445[(1'h0):(1'h0)] ~^ reg4589[(1'h0):(1'h0)]);
                      reg4694 <= reg4657[(1'h1):(1'h0)];
                      reg4695 <= ($signed($signed(reg4379)) >= reg4484[(2'h2):(1'h1)]);
                      reg4696 <= (^~($unsigned(reg4577) == (reg4424[(1'h0):(1'h0)] ?
                          $signed(reg4386) : $signed(reg4577))));
                    end
                  else
                    begin
                      reg4693 <= (|$unsigned((-(reg4612 ? reg4593 : reg4439))));
                      reg4694 <= ($signed(({reg4513} >= (8'hb6))) < (((8'ha1) ^~ (reg4644 ?
                              reg4651 : reg4532)) ?
                          $signed($unsigned(reg4675)) : reg4691));
                    end
                  for (forvar4697 = (1'h0); (forvar4697 < (2'h2)); forvar4697 = (forvar4697 + (1'h1)))
                    begin
                      reg4698 <= (forvar4690[(1'h1):(1'h0)] >= (8'ha7));
                    end
                  for (forvar4699 = (1'h0); (forvar4699 < (2'h2)); forvar4699 = (forvar4699 + (1'h1)))
                    begin
                      reg4700 <= reg4601;
                      reg4701 <= (&(reg4466 ?
                          ({reg4523} ?
                              reg4378 : reg4477[(3'h6):(1'h0)]) : (!$signed(reg4506))));
                    end
                end
            end
        end
      if ((reg4560[(4'h9):(3'h6)] > (-reg4408)))
        begin
          reg4702 <= {(reg4691 ? reg4544 : (^$unsigned(wire2)))};
          for (forvar4703 = (1'h0); (forvar4703 < (2'h3)); forvar4703 = (forvar4703 + (1'h1)))
            begin
              for (forvar4704 = (1'h0); (forvar4704 < (1'h0)); forvar4704 = (forvar4704 + (1'h1)))
                begin
                  for (forvar4705 = (1'h0); (forvar4705 < (2'h2)); forvar4705 = (forvar4705 + (1'h1)))
                    begin
                      reg4706 <= $signed(($unsigned((-(8'hb5))) ?
                          ((reg4635 <<< reg4413) ?
                              reg4667[(2'h2):(1'h0)] : $unsigned(forvar4676)) : {(reg4493 ?
                                  reg4335 : forvar4664)}));
                      reg4707 <= (8'hb0);
                    end
                  for (forvar4708 = (1'h0); (forvar4708 < (2'h3)); forvar4708 = (forvar4708 + (1'h1)))
                    begin
                      reg4709 <= (reg4373[(3'h5):(2'h2)] ?
                          $unsigned($unsigned(forvar4675)) : (((reg4379 == (8'hb1)) ?
                                  $unsigned((8'hba)) : $signed(reg4606)) ?
                              reg4482 : reg4378[(3'h4):(2'h3)]));
                    end
                  if (reg4380)
                    begin
                      reg4710 <= $signed(wire4316);
                    end
                  else
                    begin
                      reg4710 <= ((((reg4407 & reg4382) ?
                          (reg4684 ?
                              reg4530 : reg4560) : reg4456) ~^ $unsigned($unsigned(reg4695))) > (~&$signed((reg4493 ?
                          reg4695 : forvar4673))));
                      reg4711 <= (!reg4637[(3'h4):(1'h1)]);
                    end
                  for (forvar4712 = (1'h0); (forvar4712 < (2'h3)); forvar4712 = (forvar4712 + (1'h1)))
                    begin
                      reg4713 <= (($signed(((8'ha1) >= reg4376)) - $signed(((8'ha5) ?
                          forvar4671 : reg4622))) != (reg4348[(2'h3):(2'h2)] ^~ ($unsigned(reg4411) ?
                          (reg4471 << (8'h9d)) : {reg4510})));
                      reg4714 <= ({reg4422} ?
                          ((!$signed(reg4453)) ?
                              $signed($signed(reg4536)) : {(^~reg4395)}) : ($unsigned((~^reg4349)) ?
                              reg4479 : $signed(reg4696)));
                      reg4715 <= {$unsigned($signed({reg4648}))};
                    end
                end
              for (forvar4716 = (1'h0); (forvar4716 < (2'h3)); forvar4716 = (forvar4716 + (1'h1)))
                begin
                  if ($signed(reg4715))
                    begin
                      reg4717 <= {wire4661};
                      reg4718 <= $unsigned(reg4449);
                      reg4719 <= ($signed({(8'ha2)}) ^~ (reg4421 ~^ $unsigned((reg4688 | (8'h9f)))));
                    end
                  else
                    begin
                      reg4717 <= reg4589[(2'h3):(2'h3)];
                      reg4718 <= reg4557;
                      reg4719 <= reg4431[(3'h7):(3'h4)];
                    end
                  for (forvar4720 = (1'h0); (forvar4720 < (2'h3)); forvar4720 = (forvar4720 + (1'h1)))
                    begin
                      reg4721 <= reg4548[(5'h10):(2'h3)];
                      reg4722 <= reg4499[(3'h6):(1'h1)];
                      reg4723 <= reg4322[(3'h4):(3'h4)];
                    end
                end
            end
        end
      else
        begin
          reg4702 <= $signed(forvar4683[(2'h3):(2'h3)]);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4  (y, clk, wire5, wire6, wire7, wire8);
  output wire [(32'h1e80):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire5;
  input wire [(4'hc):(1'h0)] wire6;
  input wire [(4'h8):(1'h0)] wire7;
  input wire [(3'h7):(1'h0)] wire8;
  wire signed [(2'h3):(1'h0)] wire4100;
  wire [(3'h7):(1'h0)] wire4099;
  wire [(3'h5):(1'h0)] wire4098;
  wire [(3'h6):(1'h0)] wire4097;
  wire [(3'h5):(1'h0)] wire4096;
  wire signed [(3'h4):(1'h0)] wire3919;
  wire signed [(4'hf):(1'h0)] wire3721;
  wire signed [(4'h9):(1'h0)] wire3720;
  wire [(3'h7):(1'h0)] wire3636;
  wire [(3'h4):(1'h0)] wire3634;
  wire [(4'h9):(1'h0)] wire85;
  wire [(4'h9):(1'h0)] wire3632;
  reg [(4'hb):(1'h0)] reg4315 = (1'h0);
  reg [(4'he):(1'h0)] reg4314 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4313 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4312 = (1'h0);
  reg [(4'h8):(1'h0)] reg4310 = (1'h0);
  reg [(2'h3):(1'h0)] reg4309 = (1'h0);
  reg [(4'h8):(1'h0)] reg4307 = (1'h0);
  reg [(4'ha):(1'h0)] reg4306 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4305 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4304 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4302 = (1'h0);
  reg [(4'h8):(1'h0)] reg4301 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4300 = (1'h0);
  reg [(4'h9):(1'h0)] reg4299 = (1'h0);
  reg [(3'h5):(1'h0)] reg4298 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4296 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4295 = (1'h0);
  reg [(3'h7):(1'h0)] reg4294 = (1'h0);
  reg [(4'hb):(1'h0)] reg4293 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4291 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4290 = (1'h0);
  reg [(5'h10):(1'h0)] reg4286 = (1'h0);
  reg [(4'h8):(1'h0)] reg4283 = (1'h0);
  reg [(3'h7):(1'h0)] reg4289 = (1'h0);
  reg [(3'h4):(1'h0)] reg4288 = (1'h0);
  reg [(4'hb):(1'h0)] reg4287 = (1'h0);
  reg [(4'h9):(1'h0)] reg4285 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4284 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4281 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4280 = (1'h0);
  reg [(4'hd):(1'h0)] reg4279 = (1'h0);
  reg [(4'h8):(1'h0)] reg4278 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4277 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4275 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4274 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4273 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4272 = (1'h0);
  reg [(2'h3):(1'h0)] reg4271 = (1'h0);
  reg [(4'hb):(1'h0)] reg4270 = (1'h0);
  reg [(3'h5):(1'h0)] reg4268 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4265 = (1'h0);
  reg [(3'h6):(1'h0)] reg4261 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4260 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4259 = (1'h0);
  reg [(4'hc):(1'h0)] reg4258 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4249 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4248 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4239 = (1'h0);
  reg [(2'h3):(1'h0)] reg4257 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4256 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4255 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4254 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4253 = (1'h0);
  reg [(3'h7):(1'h0)] reg4251 = (1'h0);
  reg [(3'h7):(1'h0)] reg4250 = (1'h0);
  reg [(2'h2):(1'h0)] reg4247 = (1'h0);
  reg [(4'hc):(1'h0)] reg4246 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4245 = (1'h0);
  reg [(3'h5):(1'h0)] reg4244 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4243 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4242 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4241 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4240 = (1'h0);
  reg [(4'hc):(1'h0)] reg4238 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4236 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4234 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4233 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4232 = (1'h0);
  reg [(4'ha):(1'h0)] reg4231 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4230 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4229 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4228 = (1'h0);
  reg [(2'h2):(1'h0)] reg4225 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4222 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4227 = (1'h0);
  reg [(4'he):(1'h0)] reg4226 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4224 = (1'h0);
  reg [(4'hd):(1'h0)] reg4223 = (1'h0);
  reg [(5'h10):(1'h0)] reg4221 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4220 = (1'h0);
  reg [(5'h10):(1'h0)] reg4218 = (1'h0);
  reg [(4'he):(1'h0)] reg4217 = (1'h0);
  reg [(4'hc):(1'h0)] reg4215 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4212 = (1'h0);
  reg [(4'he):(1'h0)] reg4214 = (1'h0);
  reg [(4'h8):(1'h0)] reg4207 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4213 = (1'h0);
  reg [(3'h5):(1'h0)] reg4211 = (1'h0);
  reg [(4'hc):(1'h0)] reg4210 = (1'h0);
  reg [(3'h7):(1'h0)] reg4209 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4208 = (1'h0);
  reg [(3'h5):(1'h0)] reg4206 = (1'h0);
  reg [(4'hd):(1'h0)] reg4205 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4204 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4203 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4202 = (1'h0);
  reg [(5'h10):(1'h0)] reg4201 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4200 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4198 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4197 = (1'h0);
  reg [(4'ha):(1'h0)] reg4196 = (1'h0);
  reg [(4'hd):(1'h0)] reg4195 = (1'h0);
  reg [(5'h10):(1'h0)] reg4193 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4194 = (1'h0);
  reg [(4'h9):(1'h0)] reg4192 = (1'h0);
  reg [(4'he):(1'h0)] reg4191 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4190 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4189 = (1'h0);
  reg [(4'hb):(1'h0)] reg4178 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4187 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4186 = (1'h0);
  reg [(5'h10):(1'h0)] reg4185 = (1'h0);
  reg [(2'h3):(1'h0)] reg4184 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4183 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4182 = (1'h0);
  reg [(3'h6):(1'h0)] reg4181 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4180 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4179 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4175 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4174 = (1'h0);
  reg [(5'h10):(1'h0)] reg4173 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4172 = (1'h0);
  reg [(5'h10):(1'h0)] reg4171 = (1'h0);
  reg [(3'h6):(1'h0)] reg4170 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4169 = (1'h0);
  reg [(4'he):(1'h0)] reg4160 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4167 = (1'h0);
  reg [(3'h6):(1'h0)] reg4166 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4165 = (1'h0);
  reg [(4'hd):(1'h0)] reg4164 = (1'h0);
  reg [(3'h6):(1'h0)] reg4163 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4162 = (1'h0);
  reg [(4'hf):(1'h0)] reg4161 = (1'h0);
  reg [(2'h3):(1'h0)] reg4159 = (1'h0);
  reg [(4'hc):(1'h0)] reg4158 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4157 = (1'h0);
  reg [(4'hb):(1'h0)] reg4156 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4153 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4152 = (1'h0);
  reg [(2'h2):(1'h0)] reg4151 = (1'h0);
  reg [(4'ha):(1'h0)] reg4150 = (1'h0);
  reg [(4'hc):(1'h0)] reg4148 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4146 = (1'h0);
  reg [(5'h10):(1'h0)] reg4145 = (1'h0);
  reg [(4'h8):(1'h0)] reg4142 = (1'h0);
  reg [(3'h7):(1'h0)] reg4141 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4140 = (1'h0);
  reg [(3'h5):(1'h0)] reg4139 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4137 = (1'h0);
  reg [(5'h10):(1'h0)] reg4136 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4135 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4134 = (1'h0);
  reg [(3'h7):(1'h0)] reg4133 = (1'h0);
  reg [(2'h2):(1'h0)] reg4130 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4129 = (1'h0);
  reg [(4'hd):(1'h0)] reg4126 = (1'h0);
  reg [(4'hf):(1'h0)] reg4128 = (1'h0);
  reg [(3'h7):(1'h0)] reg4127 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4125 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4124 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4122 = (1'h0);
  reg [(5'h10):(1'h0)] reg4121 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4118 = (1'h0);
  reg [(3'h6):(1'h0)] reg4117 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4116 = (1'h0);
  reg [(3'h4):(1'h0)] reg4114 = (1'h0);
  reg [(4'h8):(1'h0)] reg4108 = (1'h0);
  reg [(5'h10):(1'h0)] reg4103 = (1'h0);
  reg [(4'h9):(1'h0)] reg4113 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4112 = (1'h0);
  reg [(4'h8):(1'h0)] reg4111 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4110 = (1'h0);
  reg [(3'h5):(1'h0)] reg4109 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4107 = (1'h0);
  reg [(3'h6):(1'h0)] reg4106 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4105 = (1'h0);
  reg [(4'hd):(1'h0)] reg4104 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4102 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4101 = (1'h0);
  reg [(5'h10):(1'h0)] reg4095 = (1'h0);
  reg [(2'h2):(1'h0)] reg4094 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4093 = (1'h0);
  reg [(3'h7):(1'h0)] reg4092 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4089 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4088 = (1'h0);
  reg [(3'h5):(1'h0)] reg4087 = (1'h0);
  reg [(2'h3):(1'h0)] reg4086 = (1'h0);
  reg [(4'ha):(1'h0)] reg4084 = (1'h0);
  reg [(5'h10):(1'h0)] reg4083 = (1'h0);
  reg [(4'h9):(1'h0)] reg4082 = (1'h0);
  reg [(3'h6):(1'h0)] reg4080 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4079 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4078 = (1'h0);
  reg [(3'h7):(1'h0)] reg4077 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4076 = (1'h0);
  reg [(5'h10):(1'h0)] reg4075 = (1'h0);
  reg [(4'h9):(1'h0)] reg4074 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4069 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4072 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4071 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4070 = (1'h0);
  reg [(3'h6):(1'h0)] reg4068 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4067 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4065 = (1'h0);
  reg [(3'h5):(1'h0)] reg4064 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4063 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4059 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4058 = (1'h0);
  reg [(4'h9):(1'h0)] reg4057 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4056 = (1'h0);
  reg [(4'hb):(1'h0)] reg4055 = (1'h0);
  reg [(4'h8):(1'h0)] reg4054 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4053 = (1'h0);
  reg [(3'h4):(1'h0)] reg4052 = (1'h0);
  reg [(4'he):(1'h0)] reg4051 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4050 = (1'h0);
  reg [(4'hb):(1'h0)] reg4049 = (1'h0);
  reg [(2'h2):(1'h0)] reg4047 = (1'h0);
  reg [(3'h5):(1'h0)] reg4046 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4045 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4043 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4042 = (1'h0);
  reg [(4'hf):(1'h0)] reg4040 = (1'h0);
  reg [(5'h10):(1'h0)] reg4039 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4038 = (1'h0);
  reg [(3'h4):(1'h0)] reg4037 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4036 = (1'h0);
  reg [(3'h6):(1'h0)] reg4034 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4033 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4032 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4031 = (1'h0);
  reg [(3'h7):(1'h0)] reg4030 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4028 = (1'h0);
  reg [(3'h4):(1'h0)] reg4027 = (1'h0);
  reg [(4'hc):(1'h0)] reg4026 = (1'h0);
  reg [(3'h5):(1'h0)] reg4025 = (1'h0);
  reg [(3'h6):(1'h0)] reg4022 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4021 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4020 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4019 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4017 = (1'h0);
  reg [(2'h2):(1'h0)] reg4016 = (1'h0);
  reg [(5'h10):(1'h0)] reg4015 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4014 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4013 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4012 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3999 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4011 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4010 = (1'h0);
  reg [(3'h4):(1'h0)] reg4009 = (1'h0);
  reg [(4'hd):(1'h0)] reg4008 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4007 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4006 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4005 = (1'h0);
  reg [(4'he):(1'h0)] reg4004 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4002 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4001 = (1'h0);
  reg [(4'hc):(1'h0)] reg4000 = (1'h0);
  reg [(4'ha):(1'h0)] reg3998 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3997 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3980 = (1'h0);
  reg [(2'h3):(1'h0)] reg3974 = (1'h0);
  reg [(4'hf):(1'h0)] reg3989 = (1'h0);
  reg [(4'ha):(1'h0)] reg3996 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3995 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3994 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3993 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3992 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3991 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3990 = (1'h0);
  reg [(3'h6):(1'h0)] reg3988 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3987 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3986 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3985 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3984 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3983 = (1'h0);
  reg [(4'h9):(1'h0)] reg3982 = (1'h0);
  reg [(3'h4):(1'h0)] reg3981 = (1'h0);
  reg [(4'hd):(1'h0)] reg3979 = (1'h0);
  reg [(4'hb):(1'h0)] reg3978 = (1'h0);
  reg [(3'h5):(1'h0)] reg3977 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3976 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3959 = (1'h0);
  reg [(4'hd):(1'h0)] reg3954 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3950 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3949 = (1'h0);
  reg [(2'h2):(1'h0)] reg3973 = (1'h0);
  reg [(5'h10):(1'h0)] reg3972 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3971 = (1'h0);
  reg [(3'h7):(1'h0)] reg3970 = (1'h0);
  reg [(4'hb):(1'h0)] reg3969 = (1'h0);
  reg [(4'hf):(1'h0)] reg3968 = (1'h0);
  reg [(4'hb):(1'h0)] reg3967 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3966 = (1'h0);
  reg [(4'hd):(1'h0)] reg3965 = (1'h0);
  reg [(3'h5):(1'h0)] reg3964 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3962 = (1'h0);
  reg [(3'h7):(1'h0)] reg3961 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3960 = (1'h0);
  reg [(4'hc):(1'h0)] reg3958 = (1'h0);
  reg [(4'h8):(1'h0)] reg3957 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3956 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3955 = (1'h0);
  reg [(4'ha):(1'h0)] reg3953 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3952 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3951 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3948 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3947 = (1'h0);
  reg [(3'h6):(1'h0)] reg3946 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3945 = (1'h0);
  reg [(2'h2):(1'h0)] reg3944 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3943 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3942 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3941 = (1'h0);
  reg [(4'hb):(1'h0)] reg3940 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3939 = (1'h0);
  reg [(3'h5):(1'h0)] reg3938 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3937 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3936 = (1'h0);
  reg [(3'h5):(1'h0)] reg3935 = (1'h0);
  reg [(4'ha):(1'h0)] reg3934 = (1'h0);
  reg [(3'h6):(1'h0)] reg3933 = (1'h0);
  reg [(4'ha):(1'h0)] reg3932 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3931 = (1'h0);
  reg [(2'h2):(1'h0)] reg3927 = (1'h0);
  reg [(4'hc):(1'h0)] reg3925 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3924 = (1'h0);
  reg [(5'h10):(1'h0)] reg3923 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3918 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3917 = (1'h0);
  reg [(3'h6):(1'h0)] reg3911 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3916 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3915 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3914 = (1'h0);
  reg [(3'h7):(1'h0)] reg3913 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3912 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3909 = (1'h0);
  reg [(3'h7):(1'h0)] reg3908 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3907 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3906 = (1'h0);
  reg [(3'h6):(1'h0)] reg3905 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3903 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3902 = (1'h0);
  reg [(4'hc):(1'h0)] reg3899 = (1'h0);
  reg [(3'h7):(1'h0)] reg3898 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3897 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3896 = (1'h0);
  reg [(4'h8):(1'h0)] reg3895 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3894 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3892 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3891 = (1'h0);
  reg [(4'ha):(1'h0)] reg3886 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3884 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3883 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3882 = (1'h0);
  reg [(4'hb):(1'h0)] reg3880 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3879 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3878 = (1'h0);
  reg [(3'h6):(1'h0)] reg3877 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3876 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3875 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3874 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3873 = (1'h0);
  reg [(5'h10):(1'h0)] reg3872 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3871 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3869 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3868 = (1'h0);
  reg [(4'h9):(1'h0)] reg3859 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3867 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3866 = (1'h0);
  reg [(4'h8):(1'h0)] reg3865 = (1'h0);
  reg [(2'h3):(1'h0)] reg3864 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3863 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3861 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3860 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3858 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3857 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3855 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3854 = (1'h0);
  reg [(3'h4):(1'h0)] reg3853 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3852 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3850 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3849 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3848 = (1'h0);
  reg [(4'hd):(1'h0)] reg3847 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3843 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3846 = (1'h0);
  reg [(4'ha):(1'h0)] reg3845 = (1'h0);
  reg [(5'h10):(1'h0)] reg3844 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3842 = (1'h0);
  reg [(5'h10):(1'h0)] reg3841 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3840 = (1'h0);
  reg [(4'hd):(1'h0)] reg3839 = (1'h0);
  reg [(4'h8):(1'h0)] reg3837 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3836 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3835 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3834 = (1'h0);
  reg [(5'h10):(1'h0)] reg3833 = (1'h0);
  reg [(5'h10):(1'h0)] reg3832 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3830 = (1'h0);
  reg [(4'h8):(1'h0)] reg3829 = (1'h0);
  reg [(2'h3):(1'h0)] reg3828 = (1'h0);
  reg [(5'h10):(1'h0)] reg3827 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3826 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3825 = (1'h0);
  reg [(2'h2):(1'h0)] reg3824 = (1'h0);
  reg [(4'he):(1'h0)] reg3823 = (1'h0);
  reg [(3'h5):(1'h0)] reg3822 = (1'h0);
  reg [(2'h2):(1'h0)] reg3810 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3802 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3801 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3799 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3797 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3818 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3817 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3816 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3815 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3814 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3813 = (1'h0);
  reg [(4'hf):(1'h0)] reg3812 = (1'h0);
  reg [(5'h10):(1'h0)] reg3811 = (1'h0);
  reg [(5'h10):(1'h0)] reg3809 = (1'h0);
  reg [(4'h8):(1'h0)] reg3808 = (1'h0);
  reg [(4'hf):(1'h0)] reg3807 = (1'h0);
  reg [(3'h7):(1'h0)] reg3806 = (1'h0);
  reg [(5'h10):(1'h0)] reg3805 = (1'h0);
  reg [(4'he):(1'h0)] reg3804 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3803 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3800 = (1'h0);
  reg [(4'hb):(1'h0)] reg3798 = (1'h0);
  reg [(4'hb):(1'h0)] reg3796 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3795 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3794 = (1'h0);
  reg [(4'ha):(1'h0)] reg3791 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3790 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3788 = (1'h0);
  reg [(3'h5):(1'h0)] reg3787 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3786 = (1'h0);
  reg [(2'h3):(1'h0)] reg3785 = (1'h0);
  reg [(4'hf):(1'h0)] reg3784 = (1'h0);
  reg [(4'hc):(1'h0)] reg3781 = (1'h0);
  reg [(3'h5):(1'h0)] reg3779 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3778 = (1'h0);
  reg [(3'h6):(1'h0)] reg3777 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3776 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3775 = (1'h0);
  reg [(2'h3):(1'h0)] reg3773 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3772 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3771 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3769 = (1'h0);
  reg [(2'h2):(1'h0)] reg3768 = (1'h0);
  reg [(3'h4):(1'h0)] reg3767 = (1'h0);
  reg [(3'h7):(1'h0)] reg3766 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3764 = (1'h0);
  reg [(4'ha):(1'h0)] reg3763 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3761 = (1'h0);
  reg [(4'hd):(1'h0)] reg3758 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3757 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3756 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3755 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3753 = (1'h0);
  reg [(3'h5):(1'h0)] reg3752 = (1'h0);
  reg [(4'hf):(1'h0)] reg3751 = (1'h0);
  reg [(3'h7):(1'h0)] reg3750 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3749 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3748 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3747 = (1'h0);
  reg [(4'h8):(1'h0)] reg3746 = (1'h0);
  reg [(4'h8):(1'h0)] reg3745 = (1'h0);
  reg [(2'h2):(1'h0)] reg3743 = (1'h0);
  reg [(2'h3):(1'h0)] reg3742 = (1'h0);
  reg [(4'hd):(1'h0)] reg3725 = (1'h0);
  reg [(4'hf):(1'h0)] reg3739 = (1'h0);
  reg [(4'ha):(1'h0)] reg3738 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3737 = (1'h0);
  reg [(4'h9):(1'h0)] reg3736 = (1'h0);
  reg [(3'h6):(1'h0)] reg3735 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3734 = (1'h0);
  reg [(3'h7):(1'h0)] reg3731 = (1'h0);
  reg [(4'he):(1'h0)] reg3733 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3732 = (1'h0);
  reg [(4'hb):(1'h0)] reg3730 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3729 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3728 = (1'h0);
  reg [(4'h9):(1'h0)] reg3727 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3726 = (1'h0);
  reg [(3'h4):(1'h0)] reg3724 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3723 = (1'h0);
  reg [(3'h4):(1'h0)] reg3722 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3691 = (1'h0);
  reg [(3'h4):(1'h0)] reg3719 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3718 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3717 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3716 = (1'h0);
  reg [(4'hf):(1'h0)] reg3715 = (1'h0);
  reg [(2'h2):(1'h0)] reg3714 = (1'h0);
  reg [(4'hb):(1'h0)] reg3713 = (1'h0);
  reg [(4'he):(1'h0)] reg3712 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3710 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3709 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3706 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3705 = (1'h0);
  reg [(4'hc):(1'h0)] reg3704 = (1'h0);
  reg [(4'hc):(1'h0)] reg3703 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3702 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3701 = (1'h0);
  reg [(4'hb):(1'h0)] reg3700 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3699 = (1'h0);
  reg [(4'ha):(1'h0)] reg3698 = (1'h0);
  reg [(4'h8):(1'h0)] reg3697 = (1'h0);
  reg [(5'h10):(1'h0)] reg3696 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3695 = (1'h0);
  reg [(3'h5):(1'h0)] reg3694 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3693 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3692 = (1'h0);
  reg [(2'h3):(1'h0)] reg3686 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3684 = (1'h0);
  reg [(3'h4):(1'h0)] reg3690 = (1'h0);
  reg [(3'h5):(1'h0)] reg3689 = (1'h0);
  reg [(4'h8):(1'h0)] reg3688 = (1'h0);
  reg [(4'he):(1'h0)] reg3687 = (1'h0);
  reg [(4'hd):(1'h0)] reg3685 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3683 = (1'h0);
  reg [(2'h2):(1'h0)] reg3682 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3681 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3679 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3678 = (1'h0);
  reg [(4'ha):(1'h0)] reg3677 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3675 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3674 = (1'h0);
  reg [(3'h5):(1'h0)] reg3673 = (1'h0);
  reg [(3'h4):(1'h0)] reg3672 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3670 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3669 = (1'h0);
  reg [(2'h2):(1'h0)] reg3668 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3667 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3666 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3665 = (1'h0);
  reg [(3'h7):(1'h0)] reg3656 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3648 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3662 = (1'h0);
  reg [(4'hb):(1'h0)] reg3661 = (1'h0);
  reg [(4'ha):(1'h0)] reg3660 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3659 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3658 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3657 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3655 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3654 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3649 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3653 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3652 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3651 = (1'h0);
  reg [(3'h6):(1'h0)] reg3650 = (1'h0);
  reg [(3'h6):(1'h0)] reg3647 = (1'h0);
  reg [(5'h10):(1'h0)] reg3646 = (1'h0);
  reg [(4'h9):(1'h0)] reg3645 = (1'h0);
  reg [(2'h2):(1'h0)] reg3644 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3643 = (1'h0);
  reg [(3'h6):(1'h0)] reg3642 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3641 = (1'h0);
  reg [(3'h7):(1'h0)] reg3639 = (1'h0);
  reg [(2'h2):(1'h0)] reg3640 = (1'h0);
  reg [(4'h8):(1'h0)] reg3637 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg10 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg12 = (1'h0);
  reg [(4'hb):(1'h0)] reg13 = (1'h0);
  reg [(4'hd):(1'h0)] reg15 = (1'h0);
  reg [(3'h6):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg17 = (1'h0);
  reg [(4'ha):(1'h0)] reg18 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg20 = (1'h0);
  reg [(4'hb):(1'h0)] reg21 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg22 = (1'h0);
  reg [(3'h5):(1'h0)] reg14 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg24 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg25 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg26 = (1'h0);
  reg [(4'hc):(1'h0)] reg27 = (1'h0);
  reg [(4'hc):(1'h0)] reg28 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg31 = (1'h0);
  reg [(5'h10):(1'h0)] reg32 = (1'h0);
  reg [(4'hc):(1'h0)] reg33 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg34 = (1'h0);
  reg [(2'h3):(1'h0)] reg36 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg37 = (1'h0);
  reg [(4'h9):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg43 = (1'h0);
  reg [(2'h3):(1'h0)] reg44 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg45 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg47 = (1'h0);
  reg [(4'he):(1'h0)] reg48 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg49 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg50 = (1'h0);
  reg [(4'h9):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg52 = (1'h0);
  reg [(4'h8):(1'h0)] reg53 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg54 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg57 = (1'h0);
  reg [(4'hd):(1'h0)] reg59 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg60 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg61 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg63 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg64 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg67 = (1'h0);
  reg [(3'h7):(1'h0)] reg68 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg69 = (1'h0);
  reg [(4'h9):(1'h0)] reg70 = (1'h0);
  reg [(4'he):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg72 = (1'h0);
  reg [(3'h6):(1'h0)] reg73 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg74 = (1'h0);
  reg [(4'hc):(1'h0)] reg75 = (1'h0);
  reg [(3'h4):(1'h0)] reg76 = (1'h0);
  reg [(4'hd):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg79 = (1'h0);
  reg [(3'h4):(1'h0)] reg80 = (1'h0);
  reg [(4'ha):(1'h0)] reg81 = (1'h0);
  reg [(4'hc):(1'h0)] reg83 = (1'h0);
  reg [(4'h9):(1'h0)] reg84 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4311 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4308 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4303 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4298 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4297 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4292 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4286 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4283 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4282 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4276 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4269 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4267 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4266 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4264 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4263 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4262 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4253 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4241 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4252 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4249 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4248 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4239 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4237 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4235 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4225 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4222 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4219 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4216 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4213 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4208 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4196 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4212 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4207 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4199 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4191 = (1'h0);
  reg [(4'he):(1'h0)] forvar4193 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4188 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4179 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4178 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4177 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4176 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4168 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4163 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4160 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4155 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4154 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4149 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4147 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4144 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4143 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4138 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4132 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4131 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4126 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4123 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4120 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4119 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4115 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4113 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4111 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4107 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4104 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4102 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4105 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4108 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4103 = (1'h0);
  reg [(4'he):(1'h0)] forvar4101 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4091 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4090 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4085 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4081 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4073 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4069 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4066 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4062 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4061 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4060 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4055 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4048 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4042 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4044 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4041 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4035 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4029 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4024 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4023 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4018 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4012 = (1'h0);
  reg [(4'he):(1'h0)] forvar4003 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3999 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3994 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3991 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3987 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3986 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3981 = (1'h0);
  reg [(4'he):(1'h0)] forvar3976 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3989 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3980 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3975 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3974 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3962 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3957 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3953 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3951 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3963 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3959 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3954 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3950 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3949 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3930 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3929 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3928 = (1'h0);
  reg [(4'he):(1'h0)] forvar3926 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3922 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3921 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3920 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3911 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3910 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3904 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3901 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3900 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3893 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3890 = (1'h0);
  reg [(4'he):(1'h0)] forvar3889 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3888 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3887 = (1'h0);
  reg [(4'he):(1'h0)] forvar3885 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3881 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3874 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3870 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3865 = (1'h0);
  reg [(4'he):(1'h0)] forvar3862 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3859 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3856 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3851 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3846 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3842 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3839 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3843 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3838 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3833 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3831 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3821 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3820 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3819 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3806 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3794 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3810 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3802 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3801 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3799 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3797 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3793 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3792 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3730 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3727 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3722 = (1'h0);
  reg [(4'he):(1'h0)] forvar3789 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3783 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3782 = (1'h0);
  reg [(4'he):(1'h0)] forvar3780 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3774 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3770 = (1'h0);
  reg [(4'he):(1'h0)] forvar3765 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3762 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3760 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3759 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3754 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3744 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3741 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3740 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3735 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3733 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3728 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3724 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3723 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3732 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3729 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3731 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3725 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3693 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3685 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3711 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3708 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3707 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3699 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3694 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3691 = (1'h0);
  reg [(4'he):(1'h0)] forvar3683 = (1'h0);
  reg [(4'he):(1'h0)] forvar3686 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3684 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3680 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3676 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3671 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3664 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3663 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3655 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3651 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3656 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3649 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3648 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3639 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3638 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar75 = (1'h0);
  reg [(3'h5):(1'h0)] forvar71 = (1'h0);
  reg [(4'hc):(1'h0)] forvar82 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar78 = (1'h0);
  reg [(2'h2):(1'h0)] forvar66 = (1'h0);
  reg [(5'h10):(1'h0)] forvar65 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar62 = (1'h0);
  reg [(4'hc):(1'h0)] forvar58 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar55 = (1'h0);
  reg [(2'h2):(1'h0)] forvar42 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar41 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar39 = (1'h0);
  reg [(4'hb):(1'h0)] forvar38 = (1'h0);
  reg [(3'h5):(1'h0)] forvar35 = (1'h0);
  reg [(3'h5):(1'h0)] forvar30 = (1'h0);
  reg [(2'h2):(1'h0)] forvar29 = (1'h0);
  reg [(4'h8):(1'h0)] forvar23 = (1'h0);
  reg [(3'h4):(1'h0)] forvar22 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar19 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar16 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar17 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar14 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar11 = (1'h0);
  reg [(4'hc):(1'h0)] forvar9 = (1'h0);
  assign y = {wire4100,
                 wire4099,
                 wire4098,
                 wire4097,
                 wire4096,
                 wire3919,
                 wire3721,
                 wire3720,
                 wire3636,
                 wire3634,
                 wire85,
                 wire3632,
                 reg4315,
                 reg4314,
                 reg4313,
                 reg4312,
                 reg4310,
                 reg4309,
                 reg4307,
                 reg4306,
                 reg4305,
                 reg4304,
                 reg4302,
                 reg4301,
                 reg4300,
                 reg4299,
                 reg4298,
                 reg4296,
                 reg4295,
                 reg4294,
                 reg4293,
                 reg4291,
                 reg4290,
                 reg4286,
                 reg4283,
                 reg4289,
                 reg4288,
                 reg4287,
                 reg4285,
                 reg4284,
                 reg4281,
                 reg4280,
                 reg4279,
                 reg4278,
                 reg4277,
                 reg4275,
                 reg4274,
                 reg4273,
                 reg4272,
                 reg4271,
                 reg4270,
                 reg4268,
                 reg4265,
                 reg4261,
                 reg4260,
                 reg4259,
                 reg4258,
                 reg4249,
                 reg4248,
                 reg4239,
                 reg4257,
                 reg4256,
                 reg4255,
                 reg4254,
                 reg4253,
                 reg4251,
                 reg4250,
                 reg4247,
                 reg4246,
                 reg4245,
                 reg4244,
                 reg4243,
                 reg4242,
                 reg4241,
                 reg4240,
                 reg4238,
                 reg4236,
                 reg4234,
                 reg4233,
                 reg4232,
                 reg4231,
                 reg4230,
                 reg4229,
                 reg4228,
                 reg4225,
                 reg4222,
                 reg4227,
                 reg4226,
                 reg4224,
                 reg4223,
                 reg4221,
                 reg4220,
                 reg4218,
                 reg4217,
                 reg4215,
                 reg4212,
                 reg4214,
                 reg4207,
                 reg4213,
                 reg4211,
                 reg4210,
                 reg4209,
                 reg4208,
                 reg4206,
                 reg4205,
                 reg4204,
                 reg4203,
                 reg4202,
                 reg4201,
                 reg4200,
                 reg4198,
                 reg4197,
                 reg4196,
                 reg4195,
                 reg4193,
                 reg4194,
                 reg4192,
                 reg4191,
                 reg4190,
                 reg4189,
                 reg4178,
                 reg4187,
                 reg4186,
                 reg4185,
                 reg4184,
                 reg4183,
                 reg4182,
                 reg4181,
                 reg4180,
                 reg4179,
                 reg4175,
                 reg4174,
                 reg4173,
                 reg4172,
                 reg4171,
                 reg4170,
                 reg4169,
                 reg4160,
                 reg4167,
                 reg4166,
                 reg4165,
                 reg4164,
                 reg4163,
                 reg4162,
                 reg4161,
                 reg4159,
                 reg4158,
                 reg4157,
                 reg4156,
                 reg4153,
                 reg4152,
                 reg4151,
                 reg4150,
                 reg4148,
                 reg4146,
                 reg4145,
                 reg4142,
                 reg4141,
                 reg4140,
                 reg4139,
                 reg4137,
                 reg4136,
                 reg4135,
                 reg4134,
                 reg4133,
                 reg4130,
                 reg4129,
                 reg4126,
                 reg4128,
                 reg4127,
                 reg4125,
                 reg4124,
                 reg4122,
                 reg4121,
                 reg4118,
                 reg4117,
                 reg4116,
                 reg4114,
                 reg4108,
                 reg4103,
                 reg4113,
                 reg4112,
                 reg4111,
                 reg4110,
                 reg4109,
                 reg4107,
                 reg4106,
                 reg4105,
                 reg4104,
                 reg4102,
                 reg4101,
                 reg4095,
                 reg4094,
                 reg4093,
                 reg4092,
                 reg4089,
                 reg4088,
                 reg4087,
                 reg4086,
                 reg4084,
                 reg4083,
                 reg4082,
                 reg4080,
                 reg4079,
                 reg4078,
                 reg4077,
                 reg4076,
                 reg4075,
                 reg4074,
                 reg4069,
                 reg4072,
                 reg4071,
                 reg4070,
                 reg4068,
                 reg4067,
                 reg4065,
                 reg4064,
                 reg4063,
                 reg4059,
                 reg4058,
                 reg4057,
                 reg4056,
                 reg4055,
                 reg4054,
                 reg4053,
                 reg4052,
                 reg4051,
                 reg4050,
                 reg4049,
                 reg4047,
                 reg4046,
                 reg4045,
                 reg4043,
                 reg4042,
                 reg4040,
                 reg4039,
                 reg4038,
                 reg4037,
                 reg4036,
                 reg4034,
                 reg4033,
                 reg4032,
                 reg4031,
                 reg4030,
                 reg4028,
                 reg4027,
                 reg4026,
                 reg4025,
                 reg4022,
                 reg4021,
                 reg4020,
                 reg4019,
                 reg4017,
                 reg4016,
                 reg4015,
                 reg4014,
                 reg4013,
                 reg4012,
                 reg3999,
                 reg4011,
                 reg4010,
                 reg4009,
                 reg4008,
                 reg4007,
                 reg4006,
                 reg4005,
                 reg4004,
                 reg4002,
                 reg4001,
                 reg4000,
                 reg3998,
                 reg3997,
                 reg3980,
                 reg3974,
                 reg3989,
                 reg3996,
                 reg3995,
                 reg3994,
                 reg3993,
                 reg3992,
                 reg3991,
                 reg3990,
                 reg3988,
                 reg3987,
                 reg3986,
                 reg3985,
                 reg3984,
                 reg3983,
                 reg3982,
                 reg3981,
                 reg3979,
                 reg3978,
                 reg3977,
                 reg3976,
                 reg3959,
                 reg3954,
                 reg3950,
                 reg3949,
                 reg3973,
                 reg3972,
                 reg3971,
                 reg3970,
                 reg3969,
                 reg3968,
                 reg3967,
                 reg3966,
                 reg3965,
                 reg3964,
                 reg3962,
                 reg3961,
                 reg3960,
                 reg3958,
                 reg3957,
                 reg3956,
                 reg3955,
                 reg3953,
                 reg3952,
                 reg3951,
                 reg3948,
                 reg3947,
                 reg3946,
                 reg3945,
                 reg3944,
                 reg3943,
                 reg3942,
                 reg3941,
                 reg3940,
                 reg3939,
                 reg3938,
                 reg3937,
                 reg3936,
                 reg3935,
                 reg3934,
                 reg3933,
                 reg3932,
                 reg3931,
                 reg3927,
                 reg3925,
                 reg3924,
                 reg3923,
                 reg3918,
                 reg3917,
                 reg3911,
                 reg3916,
                 reg3915,
                 reg3914,
                 reg3913,
                 reg3912,
                 reg3909,
                 reg3908,
                 reg3907,
                 reg3906,
                 reg3905,
                 reg3903,
                 reg3902,
                 reg3899,
                 reg3898,
                 reg3897,
                 reg3896,
                 reg3895,
                 reg3894,
                 reg3892,
                 reg3891,
                 reg3886,
                 reg3884,
                 reg3883,
                 reg3882,
                 reg3880,
                 reg3879,
                 reg3878,
                 reg3877,
                 reg3876,
                 reg3875,
                 reg3874,
                 reg3873,
                 reg3872,
                 reg3871,
                 reg3869,
                 reg3868,
                 reg3859,
                 reg3867,
                 reg3866,
                 reg3865,
                 reg3864,
                 reg3863,
                 reg3861,
                 reg3860,
                 reg3858,
                 reg3857,
                 reg3855,
                 reg3854,
                 reg3853,
                 reg3852,
                 reg3850,
                 reg3849,
                 reg3848,
                 reg3847,
                 reg3843,
                 reg3846,
                 reg3845,
                 reg3844,
                 reg3842,
                 reg3841,
                 reg3840,
                 reg3839,
                 reg3837,
                 reg3836,
                 reg3835,
                 reg3834,
                 reg3833,
                 reg3832,
                 reg3830,
                 reg3829,
                 reg3828,
                 reg3827,
                 reg3826,
                 reg3825,
                 reg3824,
                 reg3823,
                 reg3822,
                 reg3810,
                 reg3802,
                 reg3801,
                 reg3799,
                 reg3797,
                 reg3818,
                 reg3817,
                 reg3816,
                 reg3815,
                 reg3814,
                 reg3813,
                 reg3812,
                 reg3811,
                 reg3809,
                 reg3808,
                 reg3807,
                 reg3806,
                 reg3805,
                 reg3804,
                 reg3803,
                 reg3800,
                 reg3798,
                 reg3796,
                 reg3795,
                 reg3794,
                 reg3791,
                 reg3790,
                 reg3788,
                 reg3787,
                 reg3786,
                 reg3785,
                 reg3784,
                 reg3781,
                 reg3779,
                 reg3778,
                 reg3777,
                 reg3776,
                 reg3775,
                 reg3773,
                 reg3772,
                 reg3771,
                 reg3769,
                 reg3768,
                 reg3767,
                 reg3766,
                 reg3764,
                 reg3763,
                 reg3761,
                 reg3758,
                 reg3757,
                 reg3756,
                 reg3755,
                 reg3753,
                 reg3752,
                 reg3751,
                 reg3750,
                 reg3749,
                 reg3748,
                 reg3747,
                 reg3746,
                 reg3745,
                 reg3743,
                 reg3742,
                 reg3725,
                 reg3739,
                 reg3738,
                 reg3737,
                 reg3736,
                 reg3735,
                 reg3734,
                 reg3731,
                 reg3733,
                 reg3732,
                 reg3730,
                 reg3729,
                 reg3728,
                 reg3727,
                 reg3726,
                 reg3724,
                 reg3723,
                 reg3722,
                 reg3691,
                 reg3719,
                 reg3718,
                 reg3717,
                 reg3716,
                 reg3715,
                 reg3714,
                 reg3713,
                 reg3712,
                 reg3710,
                 reg3709,
                 reg3706,
                 reg3705,
                 reg3704,
                 reg3703,
                 reg3702,
                 reg3701,
                 reg3700,
                 reg3699,
                 reg3698,
                 reg3697,
                 reg3696,
                 reg3695,
                 reg3694,
                 reg3693,
                 reg3692,
                 reg3686,
                 reg3684,
                 reg3690,
                 reg3689,
                 reg3688,
                 reg3687,
                 reg3685,
                 reg3683,
                 reg3682,
                 reg3681,
                 reg3679,
                 reg3678,
                 reg3677,
                 reg3675,
                 reg3674,
                 reg3673,
                 reg3672,
                 reg3670,
                 reg3669,
                 reg3668,
                 reg3667,
                 reg3666,
                 reg3665,
                 reg3656,
                 reg3648,
                 reg3662,
                 reg3661,
                 reg3660,
                 reg3659,
                 reg3658,
                 reg3657,
                 reg3655,
                 reg3654,
                 reg3649,
                 reg3653,
                 reg3652,
                 reg3651,
                 reg3650,
                 reg3647,
                 reg3646,
                 reg3645,
                 reg3644,
                 reg3643,
                 reg3642,
                 reg3641,
                 reg3639,
                 reg3640,
                 reg3637,
                 reg10,
                 reg12,
                 reg13,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg14,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 reg28,
                 reg31,
                 reg32,
                 reg33,
                 reg34,
                 reg36,
                 reg37,
                 reg40,
                 reg43,
                 reg44,
                 reg45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 reg51,
                 reg52,
                 reg53,
                 reg54,
                 reg56,
                 reg57,
                 reg59,
                 reg60,
                 reg61,
                 reg63,
                 reg64,
                 reg67,
                 reg68,
                 reg69,
                 reg70,
                 reg71,
                 reg72,
                 reg73,
                 reg74,
                 reg75,
                 reg76,
                 reg77,
                 reg79,
                 reg80,
                 reg81,
                 reg83,
                 reg84,
                 forvar4311,
                 forvar4308,
                 forvar4303,
                 forvar4298,
                 forvar4297,
                 forvar4292,
                 forvar4286,
                 forvar4283,
                 forvar4282,
                 forvar4276,
                 forvar4269,
                 forvar4267,
                 forvar4266,
                 forvar4264,
                 forvar4263,
                 forvar4262,
                 forvar4253,
                 forvar4241,
                 forvar4252,
                 forvar4249,
                 forvar4248,
                 forvar4239,
                 forvar4237,
                 forvar4235,
                 forvar4225,
                 forvar4222,
                 forvar4219,
                 forvar4216,
                 forvar4213,
                 forvar4208,
                 forvar4196,
                 forvar4212,
                 forvar4207,
                 forvar4199,
                 forvar4191,
                 forvar4193,
                 forvar4188,
                 forvar4179,
                 forvar4178,
                 forvar4177,
                 forvar4176,
                 forvar4168,
                 forvar4163,
                 forvar4160,
                 forvar4155,
                 forvar4154,
                 forvar4149,
                 forvar4147,
                 forvar4144,
                 forvar4143,
                 forvar4138,
                 forvar4132,
                 forvar4131,
                 forvar4126,
                 forvar4123,
                 forvar4120,
                 forvar4119,
                 forvar4115,
                 forvar4113,
                 forvar4111,
                 forvar4107,
                 forvar4104,
                 forvar4102,
                 forvar4105,
                 forvar4108,
                 forvar4103,
                 forvar4101,
                 forvar4091,
                 forvar4090,
                 forvar4085,
                 forvar4081,
                 forvar4073,
                 forvar4069,
                 forvar4066,
                 forvar4062,
                 forvar4061,
                 forvar4060,
                 forvar4055,
                 forvar4048,
                 forvar4042,
                 forvar4044,
                 forvar4041,
                 forvar4035,
                 forvar4029,
                 forvar4024,
                 forvar4023,
                 forvar4018,
                 forvar4012,
                 forvar4003,
                 forvar3999,
                 forvar3994,
                 forvar3991,
                 forvar3987,
                 forvar3986,
                 forvar3981,
                 forvar3976,
                 forvar3989,
                 forvar3980,
                 forvar3975,
                 forvar3974,
                 forvar3962,
                 forvar3957,
                 forvar3953,
                 forvar3951,
                 forvar3963,
                 forvar3959,
                 forvar3954,
                 forvar3950,
                 forvar3949,
                 forvar3930,
                 forvar3929,
                 forvar3928,
                 forvar3926,
                 forvar3922,
                 forvar3921,
                 forvar3920,
                 forvar3911,
                 forvar3910,
                 forvar3904,
                 forvar3901,
                 forvar3900,
                 forvar3893,
                 forvar3890,
                 forvar3889,
                 forvar3888,
                 forvar3887,
                 forvar3885,
                 forvar3881,
                 forvar3874,
                 forvar3870,
                 forvar3865,
                 forvar3862,
                 forvar3859,
                 forvar3856,
                 forvar3851,
                 forvar3846,
                 forvar3842,
                 forvar3839,
                 forvar3843,
                 forvar3838,
                 forvar3833,
                 forvar3831,
                 forvar3821,
                 forvar3820,
                 forvar3819,
                 forvar3806,
                 forvar3794,
                 forvar3810,
                 forvar3802,
                 forvar3801,
                 forvar3799,
                 forvar3797,
                 forvar3793,
                 forvar3792,
                 forvar3730,
                 forvar3727,
                 forvar3722,
                 forvar3789,
                 forvar3783,
                 forvar3782,
                 forvar3780,
                 forvar3774,
                 forvar3770,
                 forvar3765,
                 forvar3762,
                 forvar3760,
                 forvar3759,
                 forvar3754,
                 forvar3744,
                 forvar3741,
                 forvar3740,
                 forvar3735,
                 forvar3733,
                 forvar3728,
                 forvar3724,
                 forvar3723,
                 forvar3732,
                 forvar3729,
                 forvar3731,
                 forvar3725,
                 forvar3693,
                 forvar3685,
                 forvar3711,
                 forvar3708,
                 forvar3707,
                 forvar3699,
                 forvar3694,
                 forvar3691,
                 forvar3683,
                 forvar3686,
                 forvar3684,
                 forvar3680,
                 forvar3676,
                 forvar3671,
                 forvar3664,
                 forvar3663,
                 forvar3655,
                 forvar3651,
                 forvar3656,
                 forvar3649,
                 forvar3648,
                 forvar3639,
                 forvar3638,
                 forvar75,
                 forvar71,
                 forvar82,
                 forvar78,
                 forvar66,
                 forvar65,
                 forvar62,
                 forvar58,
                 forvar55,
                 forvar42,
                 forvar41,
                 forvar39,
                 forvar38,
                 forvar35,
                 forvar30,
                 forvar29,
                 forvar23,
                 forvar22,
                 forvar19,
                 forvar16,
                 forvar17,
                 forvar14,
                 forvar11,
                 forvar9,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar9 = (1'h0); (forvar9 < (1'h0)); forvar9 = (forvar9 + (1'h1)))
        begin
          reg10 <= $unsigned({$signed((^~forvar9))});
          if ((!$unsigned((forvar9[(3'h5):(3'h4)] ?
              (reg10 && wire7) : (8'ha9)))))
            begin
              for (forvar11 = (1'h0); (forvar11 < (1'h0)); forvar11 = (forvar11 + (1'h1)))
                begin
                  if ({($signed($unsigned(reg10)) ^~ (8'hba))})
                    begin
                      reg12 <= ($signed(forvar11[(2'h3):(2'h2)]) != $unsigned(($signed(wire6) ?
                          (wire8 ? (8'ha7) : wire5) : $signed(wire5))));
                      reg13 <= {((reg12 || wire5[(1'h1):(1'h0)]) ?
                              ((reg12 ? wire7 : (8'h9d)) ?
                                  ((8'hb3) + (8'hb6)) : {forvar9}) : ((wire5 ?
                                      wire8 : forvar11) ?
                                  forvar9[(4'h9):(3'h7)] : forvar11))};
                    end
                  else
                    begin
                      reg12 <= ((($unsigned(wire6) ^ wire7) ?
                          $signed((^forvar9)) : $unsigned((wire7 ?
                              wire7 : wire5))) ^ (((+(8'h9f)) - $signed(reg13)) <<< forvar9[(4'h8):(1'h0)]));
                    end
                end
              if (forvar9[(4'hb):(4'h8)])
                begin
                  for (forvar14 = (1'h0); (forvar14 < (2'h2)); forvar14 = (forvar14 + (1'h1)))
                    begin
                      reg15 <= (forvar14 > reg13);
                      reg16 <= $signed(reg13[(3'h6):(2'h2)]);
                      reg17 <= reg16[(3'h5):(3'h5)];
                    end
                  if ($unsigned(wire8[(3'h5):(1'h0)]))
                    begin
                      reg18 <= ($unsigned(((forvar11 ? (8'ha0) : forvar11) ?
                          wire5[(2'h3):(1'h1)] : forvar14)) || {({reg16} * $signed(forvar9))});
                    end
                  else
                    begin
                      reg18 <= (reg18 ^ {reg10[(4'hd):(4'hb)]});
                      reg19 <= (wire7[(2'h3):(1'h0)] > reg10[(4'h8):(4'h8)]);
                    end
                  if (($unsigned((wire5[(1'h1):(1'h1)] ?
                      (reg12 ^~ reg15) : reg16)) - $signed(((reg10 ?
                          wire6 : forvar11) ?
                      reg17 : (!reg16)))))
                    begin
                      reg20 <= $unsigned($unsigned($signed((reg18 ?
                          wire8 : reg10))));
                    end
                  else
                    begin
                      reg20 <= {($signed({wire7}) ?
                              (forvar11[(4'h8):(3'h5)] <= wire5) : ($signed(wire5) ?
                                  {reg15} : (+wire7)))};
                      reg21 <= (reg10 ? {(~|(~&forvar9))} : wire5);
                      reg22 <= $signed({($signed(reg12) || (reg16 ?
                              (8'haa) : reg18))});
                    end
                end
              else
                begin
                  reg14 <= reg12[(1'h1):(1'h0)];
                  if (reg16)
                    begin
                      reg15 <= $unsigned((wire8 <<< (((8'hb5) >> reg18) | (&forvar9))));
                    end
                  else
                    begin
                      reg15 <= reg21[(4'h9):(4'h9)];
                      reg16 <= {($signed(reg18) ? forvar14 : (~^{(8'h9d)}))};
                    end
                  for (forvar17 = (1'h0); (forvar17 < (1'h1)); forvar17 = (forvar17 + (1'h1)))
                    begin
                      reg18 <= reg12;
                      reg19 <= (^((~forvar11) * $signed(reg21[(4'h9):(3'h5)])));
                      reg20 <= wire7[(4'h8):(2'h2)];
                    end
                end
            end
          else
            begin
              for (forvar11 = (1'h0); (forvar11 < (1'h1)); forvar11 = (forvar11 + (1'h1)))
                begin
                  if ({$signed((^$signed(reg14)))})
                    begin
                      reg12 <= {(wire5 ?
                              (forvar11[(1'h1):(1'h1)] != reg12[(2'h2):(2'h2)]) : reg15)};
                    end
                  else
                    begin
                      reg12 <= reg14[(1'h0):(1'h0)];
                      reg13 <= ((($signed(forvar11) != (forvar17 ?
                                  forvar11 : forvar17)) ?
                              reg22[(2'h3):(2'h2)] : ($signed(forvar11) <<< $unsigned(wire7))) ?
                          ({forvar17} || ((wire6 ?
                              reg12 : (8'ha7)) && (reg16 & reg10))) : {forvar9});
                      reg14 <= $unsigned(reg22);
                      reg15 <= {{{$unsigned(wire5)}}};
                    end
                end
              for (forvar16 = (1'h0); (forvar16 < (1'h1)); forvar16 = (forvar16 + (1'h1)))
                begin
                  if ($signed($signed(reg22)))
                    begin
                      reg17 <= $unsigned((reg15 ?
                          $signed(((8'ha0) ?
                              (8'ha7) : wire5)) : {$unsigned(wire7)}));
                      reg18 <= $unsigned(reg21[(4'ha):(3'h4)]);
                    end
                  else
                    begin
                      reg17 <= (^~$unsigned(reg20[(3'h4):(2'h3)]));
                    end
                  for (forvar19 = (1'h0); (forvar19 < (2'h2)); forvar19 = (forvar19 + (1'h1)))
                    begin
                      reg20 <= $signed({reg12});
                      reg21 <= ($unsigned({reg15[(4'hd):(4'hc)]}) ?
                          reg19 : $signed($unsigned((reg12 ^~ reg18))));
                    end
                end
              for (forvar22 = (1'h0); (forvar22 < (1'h1)); forvar22 = (forvar22 + (1'h1)))
                begin
                  for (forvar23 = (1'h0); (forvar23 < (2'h2)); forvar23 = (forvar23 + (1'h1)))
                    begin
                      reg24 <= ((((-reg21) <= wire8) ?
                              (!$signed(forvar11)) : (~{reg16})) ?
                          forvar23 : $signed(((reg19 > reg16) <<< wire6[(3'h7):(3'h4)])));
                      reg25 <= {(!($unsigned((8'hb3)) ?
                              (forvar14 ?
                                  (8'hb2) : reg22) : forvar19[(3'h7):(1'h0)]))};
                      reg26 <= reg20[(3'h4):(1'h1)];
                      reg27 <= {(~(8'ha3))};
                    end
                  reg28 <= reg20;
                end
            end
          for (forvar29 = (1'h0); (forvar29 < (1'h0)); forvar29 = (forvar29 + (1'h1)))
            begin
              for (forvar30 = (1'h0); (forvar30 < (2'h2)); forvar30 = (forvar30 + (1'h1)))
                begin
                  if ($signed(wire7))
                    begin
                      reg31 <= $unsigned($signed((8'h9e)));
                    end
                  else
                    begin
                      reg31 <= forvar30[(2'h3):(2'h3)];
                      reg32 <= ((^$signed((&reg12))) ?
                          $signed(reg22[(1'h1):(1'h1)]) : (~^((8'ha5) >> (forvar16 ?
                              forvar22 : wire6))));
                      reg33 <= reg12[(2'h3):(2'h2)];
                      reg34 <= $unsigned(reg28[(1'h0):(1'h0)]);
                    end
                  for (forvar35 = (1'h0); (forvar35 < (2'h2)); forvar35 = (forvar35 + (1'h1)))
                    begin
                      reg36 <= (((+$unsigned((8'ha3))) || reg16[(3'h6):(1'h0)]) + (~&reg19));
                      reg37 <= reg20;
                    end
                end
              for (forvar38 = (1'h0); (forvar38 < (2'h3)); forvar38 = (forvar38 + (1'h1)))
                begin
                  for (forvar39 = (1'h0); (forvar39 < (1'h0)); forvar39 = (forvar39 + (1'h1)))
                    begin
                      reg40 <= $unsigned(forvar17);
                    end
                end
              for (forvar41 = (1'h0); (forvar41 < (1'h1)); forvar41 = (forvar41 + (1'h1)))
                begin
                  for (forvar42 = (1'h0); (forvar42 < (2'h2)); forvar42 = (forvar42 + (1'h1)))
                    begin
                      reg43 <= forvar16;
                      reg44 <= $signed($signed(wire8));
                      reg45 <= (forvar17[(1'h1):(1'h1)] * $unsigned(reg14[(3'h4):(1'h0)]));
                      reg46 <= ($unsigned((wire5[(1'h1):(1'h1)] ?
                          $unsigned((8'ha1)) : {wire7})) ^~ (!($signed(reg26) ?
                          (reg13 ? reg21 : reg27) : forvar41[(4'hc):(1'h0)])));
                    end
                  if (reg28)
                    begin
                      reg47 <= (!(((&forvar41) | $signed(reg21)) ?
                          forvar35[(2'h2):(1'h1)] : ((~^reg13) ?
                              {reg46} : reg13[(2'h3):(2'h3)])));
                    end
                  else
                    begin
                      reg47 <= reg44[(2'h2):(1'h0)];
                      reg48 <= ((reg27 | reg10[(3'h5):(2'h2)]) ?
                          reg34[(1'h1):(1'h0)] : (8'hb6));
                      reg49 <= (($unsigned((reg44 <<< reg36)) <= ($unsigned((8'ha6)) ?
                          (+wire5) : (reg14 + reg24))) > (reg31[(2'h3):(1'h1)] ?
                          ($signed(reg15) ~^ $unsigned((8'ha0))) : (!(~|reg45))));
                      reg50 <= (($unsigned({reg36}) ?
                          reg40[(2'h3):(1'h0)] : $unsigned((reg13 ^~ reg17))) && ($signed((reg19 ?
                          wire6 : reg20)) ^~ $signed((reg48 ?
                          reg43 : (8'haf)))));
                    end
                  if (wire5[(1'h1):(1'h0)])
                    begin
                      reg51 <= {$signed(reg28)};
                      reg52 <= $unsigned(forvar19[(2'h2):(2'h2)]);
                      reg53 <= (forvar9[(2'h2):(1'h1)] ^ ($unsigned($signed((8'hab))) | (^~$signed(reg26))));
                      reg54 <= $signed($unsigned(reg46));
                    end
                  else
                    begin
                      reg51 <= {$unsigned($unsigned((8'hb0)))};
                      reg52 <= ($signed(wire5) > $signed(($unsigned(reg44) ?
                          $unsigned(reg18) : $unsigned(forvar23))));
                    end
                  for (forvar55 = (1'h0); (forvar55 < (1'h0)); forvar55 = (forvar55 + (1'h1)))
                    begin
                      reg56 <= $unsigned($unsigned({(|forvar39)}));
                      reg57 <= ($unsigned($unsigned($unsigned(reg19))) ?
                          (~^$signed((reg33 ?
                              reg52 : reg27))) : $signed(((reg31 > reg40) ?
                              ((8'hb8) >> reg22) : {reg21})));
                    end
                end
              for (forvar58 = (1'h0); (forvar58 < (1'h0)); forvar58 = (forvar58 + (1'h1)))
                begin
                  if (reg53[(1'h1):(1'h0)])
                    begin
                      reg59 <= $signed((({(8'hb9)} ?
                          (&reg13) : forvar11) && forvar22));
                      reg60 <= $signed((8'hb1));
                      reg61 <= (({$signed(forvar42)} ?
                              (~&wire6[(1'h1):(1'h1)]) : $unsigned($signed(wire8))) ?
                          reg14 : (^$signed(wire6)));
                    end
                  else
                    begin
                      reg59 <= ({reg24[(1'h1):(1'h1)]} | ((|(reg25 ?
                          reg13 : reg37)) >>> $signed((reg24 || reg49))));
                      reg60 <= ((forvar17 >= ($signed((8'ha4)) ?
                              $signed(wire8) : forvar58)) ?
                          reg25[(3'h7):(3'h6)] : $signed((!(reg12 ?
                              forvar17 : reg28))));
                    end
                  for (forvar62 = (1'h0); (forvar62 < (1'h1)); forvar62 = (forvar62 + (1'h1)))
                    begin
                      reg63 <= {forvar55[(1'h1):(1'h1)]};
                    end
                  reg64 <= (reg25[(2'h2):(1'h1)] ?
                      (8'hb9) : reg13[(2'h3):(1'h1)]);
                end
            end
          for (forvar65 = (1'h0); (forvar65 < (1'h0)); forvar65 = (forvar65 + (1'h1)))
            begin
              for (forvar66 = (1'h0); (forvar66 < (1'h1)); forvar66 = (forvar66 + (1'h1)))
                begin
                  if ({(wire7 < (+$unsigned(forvar58)))})
                    begin
                      reg67 <= ((~((reg63 ?
                          reg34 : reg16) << (reg14 ~^ forvar66))) ^~ wire7[(1'h1):(1'h0)]);
                      reg68 <= ({{forvar38[(3'h4):(2'h3)]}} ?
                          (8'h9f) : $signed((&{forvar39})));
                    end
                  else
                    begin
                      reg67 <= $unsigned(reg32);
                      reg68 <= (reg18 ? forvar42 : (|(~^$signed(reg28))));
                      reg69 <= (8'hae);
                    end
                  if ((^(-((+(8'h9d)) >>> (reg49 & forvar17)))))
                    begin
                      reg70 <= reg57;
                    end
                  else
                    begin
                      reg70 <= forvar17;
                    end
                end
              if ($signed(((reg44[(1'h1):(1'h1)] > $signed(reg25)) ^ $signed((8'ha8)))))
                begin
                  if (reg24)
                    begin
                      reg71 <= ({(wire8[(2'h3):(1'h0)] ?
                                  (~|reg57) : (reg18 ? reg28 : forvar9))} ?
                          (^(reg10[(4'h9):(4'h9)] - (forvar41 <<< reg22))) : $signed(reg37));
                      reg72 <= reg28;
                      reg73 <= ((($unsigned(reg72) ~^ reg49) & $signed((reg53 ?
                              reg68 : reg19))) ?
                          $signed(reg19[(2'h3):(2'h2)]) : forvar29);
                      reg74 <= ((-(reg47 ? (~^(8'ha5)) : $unsigned(reg16))) ?
                          $signed((+(reg15 | forvar22))) : (~&{(reg60 ?
                                  reg37 : reg56)}));
                    end
                  else
                    begin
                      reg71 <= $signed(forvar11);
                      reg72 <= ((^~reg72[(3'h5):(3'h4)]) || reg60[(3'h4):(2'h2)]);
                    end
                  if ((($signed($signed(wire6)) < (reg15[(3'h4):(2'h3)] != (forvar11 ?
                          reg45 : reg67))) ?
                      $signed(reg54) : ((+forvar65) ?
                          ((~^(8'h9d)) && (~^forvar14)) : (^(wire6 ?
                              reg18 : reg64)))))
                    begin
                      reg75 <= $unsigned(reg73);
                      reg76 <= $signed($unsigned(($unsigned(reg46) ?
                          (&reg12) : (reg14 << (8'hae)))));
                      reg77 <= (reg70[(3'h4):(1'h1)] & $unsigned(reg49));
                    end
                  else
                    begin
                      reg75 <= {($signed((^forvar38)) - $unsigned({forvar39}))};
                      reg76 <= ($unsigned(((forvar55 ? reg24 : forvar55) ?
                              $unsigned(reg77) : reg75[(2'h3):(2'h2)])) ?
                          ($signed($signed(forvar42)) ?
                              ($signed(reg34) <= $unsigned(reg13)) : $signed(reg25)) : reg12[(2'h3):(2'h2)]);
                      reg77 <= $unsigned({reg33});
                    end
                  for (forvar78 = (1'h0); (forvar78 < (2'h2)); forvar78 = (forvar78 + (1'h1)))
                    begin
                      reg79 <= (forvar16[(1'h1):(1'h0)] ?
                          (!$unsigned($unsigned(reg37))) : $signed((8'hba)));
                      reg80 <= $unsigned($signed(((forvar14 ? reg50 : (8'hb6)) ?
                          wire6[(3'h7):(1'h1)] : (|reg69))));
                      reg81 <= {{(~&(reg49 <= forvar78))}};
                    end
                  for (forvar82 = (1'h0); (forvar82 < (1'h1)); forvar82 = (forvar82 + (1'h1)))
                    begin
                      reg83 <= $unsigned($signed(forvar42[(1'h0):(1'h0)]));
                      reg84 <= reg37[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar71 = (1'h0); (forvar71 < (2'h2)); forvar71 = (forvar71 + (1'h1)))
                    begin
                      reg72 <= reg22[(4'h9):(4'h8)];
                    end
                  if (reg49)
                    begin
                      reg73 <= ({$unsigned($unsigned(forvar62))} ?
                          $unsigned((~(reg31 <= reg51))) : ($unsigned((-forvar65)) ?
                              {reg70} : wire5));
                      reg74 <= $unsigned((($signed((8'hb9)) ?
                          reg61 : $unsigned(wire7)) & (+reg40)));
                    end
                  else
                    begin
                      reg73 <= reg75[(2'h2):(1'h0)];
                      reg74 <= forvar35[(3'h5):(2'h2)];
                    end
                  for (forvar75 = (1'h0); (forvar75 < (2'h3)); forvar75 = (forvar75 + (1'h1)))
                    begin
                      reg76 <= ((8'ha4) ?
                          {(~|(forvar11 == forvar19))} : (!$unsigned((reg49 ^ forvar71))));
                    end
                end
            end
        end
    end
  assign wire85 = (&reg67);
  module86 #() modinst3633 (.clk(clk), .y(wire3632), .wire89(reg31), .wire90(reg40), .wire87(wire85), .wire88(reg77));
  module3045 #() modinst3635 (.wire3049(reg45), .clk(clk), .y(wire3634), .wire3048(reg18), .wire3047(reg27), .wire3046(reg68));
  assign wire3636 = $unsigned(wire3632[(3'h6):(1'h1)]);
  always
    @(posedge clk) begin
      reg3637 <= reg37;
      for (forvar3638 = (1'h0); (forvar3638 < (2'h3)); forvar3638 = (forvar3638 + (1'h1)))
        begin
          if (reg53[(1'h0):(1'h0)])
            begin
              if ($signed((|$unsigned((forvar3638 <= reg21)))))
                begin
                  for (forvar3639 = (1'h0); (forvar3639 < (2'h3)); forvar3639 = (forvar3639 + (1'h1)))
                    begin
                      reg3640 <= (|(wire5 < (((8'hb1) ? reg51 : (8'h9d)) ?
                          (reg59 ? reg75 : reg46) : $signed((8'hba)))));
                    end
                end
              else
                begin
                  reg3639 <= (reg13 <= ({reg84} ?
                      $unsigned($signed((8'ha6))) : (8'ha4)));
                end
            end
          else
            begin
              for (forvar3639 = (1'h0); (forvar3639 < (2'h3)); forvar3639 = (forvar3639 + (1'h1)))
                begin
                  if (((8'ha4) ?
                      (($signed((8'hac)) ?
                          (reg10 <= reg18) : (~&reg56)) <= ((reg50 ?
                          reg28 : reg31) >= $unsigned((8'hac)))) : ((reg45 ?
                          reg33[(2'h3):(2'h2)] : (wire3632 | reg33)) * reg84)))
                    begin
                      reg3640 <= ({{(~reg10)}} ?
                          ($signed($unsigned(wire7)) != {(|reg15)}) : reg61);
                      reg3641 <= reg75[(2'h2):(1'h0)];
                      reg3642 <= $signed(reg69);
                      reg3643 <= $unsigned((reg26 < (-(reg45 ?
                          reg25 : wire3634))));
                    end
                  else
                    begin
                      reg3640 <= (&(!$unsigned(((8'ha4) >= (8'h9c)))));
                      reg3641 <= {$signed(reg40)};
                      reg3642 <= {$signed($unsigned(reg26))};
                    end
                  if ($unsigned((reg3643[(2'h3):(2'h2)] ?
                      reg43[(3'h6):(1'h1)] : {(^reg32)})))
                    begin
                      reg3644 <= ($signed(reg21) ? (~&{{reg22}}) : reg68);
                      reg3645 <= reg37[(1'h1):(1'h0)];
                      reg3646 <= (($signed((&reg83)) ?
                              $unsigned(reg79[(3'h5):(3'h4)]) : $signed(reg47)) ?
                          $signed($signed((reg33 >> reg15))) : $signed($unsigned(reg3645[(1'h0):(1'h0)])));
                      reg3647 <= ((^~$signed((reg3642 || reg15))) ?
                          {{(^reg47)}} : (!{(reg75 && reg81)}));
                    end
                  else
                    begin
                      reg3644 <= ((($unsigned((8'hb1)) <= ((8'hb4) <<< wire85)) != ((^~reg83) ?
                          (reg72 ~^ reg22) : $unsigned(reg3640))) << $signed(reg31));
                      reg3645 <= wire3636;
                      reg3646 <= reg67;
                    end
                end
            end
          if ($unsigned($signed(reg60)))
            begin
              for (forvar3648 = (1'h0); (forvar3648 < (2'h3)); forvar3648 = (forvar3648 + (1'h1)))
                begin
                  for (forvar3649 = (1'h0); (forvar3649 < (2'h3)); forvar3649 = (forvar3649 + (1'h1)))
                    begin
                      reg3650 <= (|reg3646);
                      reg3651 <= (reg14 == reg56);
                      reg3652 <= ({(reg26[(2'h3):(2'h2)] >>> {reg28})} ?
                          reg53 : reg44[(1'h1):(1'h0)]);
                      reg3653 <= {(8'hb9)};
                    end
                end
            end
          else
            begin
              if (($signed(((forvar3639 == reg64) ^~ reg46)) + $unsigned(reg63[(1'h1):(1'h1)])))
                begin
                  for (forvar3648 = (1'h0); (forvar3648 < (2'h2)); forvar3648 = (forvar3648 + (1'h1)))
                    begin
                      reg3649 <= (^reg67);
                      reg3650 <= (reg59[(2'h3):(2'h2)] + {{(~&reg3639)}});
                      reg3651 <= (&(reg3641[(4'hb):(1'h1)] <<< {reg43[(1'h0):(1'h0)]}));
                      reg3652 <= (($signed((&reg47)) ?
                          reg77 : {{reg3649}}) * (~((+reg3644) < $signed(reg26))));
                    end
                  if ($unsigned($unsigned((8'hb9))))
                    begin
                      reg3653 <= (!(reg3642 <= ($signed(wire85) & {reg49})));
                      reg3654 <= ((8'haf) ? reg56[(3'h4):(1'h1)] : reg75);
                      reg3655 <= $signed(((reg76[(2'h3):(1'h0)] && reg83) ^ ((reg3654 ?
                          reg56 : reg3649) && $unsigned(reg46))));
                    end
                  else
                    begin
                      reg3653 <= reg73[(2'h2):(1'h0)];
                      reg3654 <= $signed($signed($unsigned((&reg16))));
                    end
                  for (forvar3656 = (1'h0); (forvar3656 < (1'h0)); forvar3656 = (forvar3656 + (1'h1)))
                    begin
                      reg3657 <= ($signed(reg63[(1'h0):(1'h0)]) ?
                          reg21[(2'h2):(2'h2)] : $unsigned((+$signed(wire3634))));
                      reg3658 <= reg20;
                      reg3659 <= (wire3636 || $unsigned($signed(reg3652[(1'h0):(1'h0)])));
                    end
                  if ((~&$signed($unsigned((8'hb9)))))
                    begin
                      reg3660 <= ($signed((^(reg37 ?
                          reg3659 : reg52))) != (+((reg71 != reg3637) > reg12)));
                    end
                  else
                    begin
                      reg3660 <= (reg33[(4'h8):(3'h4)] ?
                          $unsigned(((reg3659 ?
                              reg3653 : (8'ha0)) ^ ((8'hac) << reg59))) : $unsigned((reg3637[(3'h4):(3'h4)] <= $signed(reg32))));
                      reg3661 <= ($signed((+reg43[(4'hb):(3'h5)])) ?
                          (((reg21 ? reg22 : (8'ha3)) ?
                                  $unsigned(reg69) : $signed(reg13)) ?
                              reg37 : reg3643[(4'hb):(4'h9)]) : (($unsigned(reg21) + wire6) ?
                              (^~reg3660) : $signed($signed(wire3634))));
                      reg3662 <= ((~&reg79) ?
                          $signed(($signed(reg68) && (reg45 + reg64))) : $signed($signed(reg80[(2'h2):(2'h2)])));
                    end
                end
              else
                begin
                  if ($signed(($signed({reg17}) ?
                      ((8'ha0) & {wire5}) : (8'ha5))))
                    begin
                      reg3648 <= $signed((((+reg3646) ?
                          {reg83} : reg3641) & $unsigned((forvar3649 & reg34))));
                      reg3649 <= {reg76};
                      reg3650 <= (((reg3659 && reg73[(3'h6):(3'h6)]) ?
                              reg37[(2'h2):(1'h0)] : (reg76[(2'h3):(2'h2)] <= $signed(reg3662))) ?
                          ({{(8'hb4)}} && (reg64[(2'h2):(1'h1)] ?
                              (^~(8'ha1)) : reg3661[(4'h8):(4'h8)])) : ($signed(wire3632) != (~((8'hb1) ~^ (8'h9c)))));
                    end
                  else
                    begin
                      reg3648 <= ((reg69[(2'h2):(2'h2)] ?
                              ((+reg3651) >> (~^reg22)) : $signed(reg46)) ?
                          $signed((|$unsigned(reg63))) : $unsigned({$unsigned(forvar3649)}));
                      reg3649 <= $unsigned((($unsigned(reg12) ?
                          $unsigned(reg45) : reg3643[(4'h9):(3'h4)]) > reg75));
                      reg3650 <= (((reg3642 ?
                              {reg3648} : (~reg20)) || reg15[(2'h3):(1'h1)]) ?
                          reg3650[(1'h0):(1'h0)] : (((~&reg83) ?
                                  $signed(reg84) : reg72) ?
                              $signed($signed(reg28)) : reg74));
                    end
                  for (forvar3651 = (1'h0); (forvar3651 < (2'h2)); forvar3651 = (forvar3651 + (1'h1)))
                    begin
                      reg3652 <= $unsigned($unsigned((((8'had) != reg46) ?
                          (reg3655 ? reg15 : reg3639) : (|reg67))));
                      reg3653 <= {reg19};
                      reg3654 <= reg25;
                    end
                  for (forvar3655 = (1'h0); (forvar3655 < (2'h2)); forvar3655 = (forvar3655 + (1'h1)))
                    begin
                      reg3656 <= {{{(reg40 | reg3662)}}};
                      reg3657 <= ($signed($unsigned((8'ha2))) ?
                          ($unsigned($unsigned(reg17)) ?
                              (reg44 ?
                                  (&reg79) : wire3632) : reg24[(3'h5):(3'h5)]) : ($signed((reg15 << reg3643)) ?
                              {wire3634} : $signed($unsigned(reg53))));
                    end
                end
              for (forvar3663 = (1'h0); (forvar3663 < (2'h2)); forvar3663 = (forvar3663 + (1'h1)))
                begin
                  for (forvar3664 = (1'h0); (forvar3664 < (1'h1)); forvar3664 = (forvar3664 + (1'h1)))
                    begin
                      reg3665 <= (^(!$unsigned(reg25)));
                      reg3666 <= $unsigned(((reg40[(3'h6):(3'h6)] ?
                          (reg18 ? reg21 : wire6) : (&reg67)) & wire3636));
                      reg3667 <= {$unsigned((&((8'hb5) + (8'hb1))))};
                    end
                  if (reg64)
                    begin
                      reg3668 <= $unsigned($signed((^$unsigned(wire85))));
                      reg3669 <= $signed((8'h9c));
                      reg3670 <= $unsigned({((wire7 - (8'hba)) ?
                              (reg68 ? reg64 : reg3655) : (^~reg32))});
                    end
                  else
                    begin
                      reg3668 <= (((wire3634[(2'h2):(1'h1)] > $unsigned((8'haf))) || ((^~reg13) ?
                          (^~reg34) : $unsigned(reg3658))) != reg3659[(3'h4):(3'h4)]);
                      reg3669 <= {reg15};
                    end
                  for (forvar3671 = (1'h0); (forvar3671 < (2'h3)); forvar3671 = (forvar3671 + (1'h1)))
                    begin
                      reg3672 <= $signed((forvar3656 ?
                          $signed(reg67) : $unsigned((forvar3664 ?
                              forvar3648 : reg18))));
                      reg3673 <= (!(reg18 ^~ reg84[(2'h3):(2'h3)]));
                      reg3674 <= (&$unsigned((^(reg22 ^ reg40))));
                      reg3675 <= {$signed(reg10)};
                    end
                  for (forvar3676 = (1'h0); (forvar3676 < (1'h1)); forvar3676 = (forvar3676 + (1'h1)))
                    begin
                      reg3677 <= $unsigned((+forvar3671));
                    end
                end
            end
        end
      reg3678 <= reg52[(3'h6):(1'h0)];
      if (forvar3651)
        begin
          reg3679 <= $signed((8'ha9));
        end
      else
        begin
          reg3679 <= ({(+$signed(reg3641))} ?
              ($signed((reg75 ?
                  reg49 : wire5)) ^~ ((^~reg68) << $signed(reg14))) : forvar3655);
          if ((~(~&((8'had) ? reg50 : $signed(forvar3639)))))
            begin
              if ($signed(reg56))
                begin
                  for (forvar3680 = (1'h0); (forvar3680 < (2'h2)); forvar3680 = (forvar3680 + (1'h1)))
                    begin
                      reg3681 <= $signed(((&forvar3671[(1'h0):(1'h0)]) ?
                          (8'h9c) : forvar3649));
                      reg3682 <= (reg31 + {($signed(wire85) - $unsigned(reg34))});
                      reg3683 <= ($unsigned((~&$unsigned(reg22))) ?
                          $unsigned((&(reg3672 != reg3674))) : reg17);
                    end
                  for (forvar3684 = (1'h0); (forvar3684 < (2'h2)); forvar3684 = (forvar3684 + (1'h1)))
                    begin
                      reg3685 <= (&$unsigned(reg51));
                    end
                  for (forvar3686 = (1'h0); (forvar3686 < (2'h2)); forvar3686 = (forvar3686 + (1'h1)))
                    begin
                      reg3687 <= (reg76[(2'h3):(2'h2)] ?
                          $unsigned((reg67[(3'h6):(3'h5)] ?
                              $signed(reg3642) : reg3675[(1'h1):(1'h0)])) : (((reg74 ^~ reg3641) ?
                              (reg13 ? reg17 : reg3667) : (reg3678 ?
                                  reg3641 : reg3666)) - {(&forvar3648)}));
                      reg3688 <= $unsigned(((~|reg46[(3'h4):(2'h2)]) < $signed(wire3634[(1'h0):(1'h0)])));
                      reg3689 <= (reg80 ?
                          $unsigned($signed((reg3665 ?
                              (8'hb8) : reg83))) : reg3668[(1'h0):(1'h0)]);
                      reg3690 <= reg83[(4'h8):(4'h8)];
                    end
                end
              else
                begin
                  for (forvar3680 = (1'h0); (forvar3680 < (2'h3)); forvar3680 = (forvar3680 + (1'h1)))
                    begin
                      reg3681 <= (reg25[(2'h2):(1'h0)] ?
                          reg68 : $unsigned((~^(~reg3675))));
                    end
                  if ($signed((+({reg3687} ? forvar3684 : reg21))))
                    begin
                      reg3682 <= reg3658[(4'h9):(4'h9)];
                    end
                  else
                    begin
                      reg3682 <= (~&reg3675);
                    end
                  for (forvar3683 = (1'h0); (forvar3683 < (2'h2)); forvar3683 = (forvar3683 + (1'h1)))
                    begin
                      reg3684 <= forvar3656[(1'h1):(1'h0)];
                      reg3685 <= $signed((^reg10[(1'h0):(1'h0)]));
                      reg3686 <= reg57[(3'h5):(2'h3)];
                      reg3687 <= {$signed(reg63[(1'h1):(1'h1)])};
                    end
                end
              if ($unsigned(reg14[(3'h5):(1'h1)]))
                begin
                  for (forvar3691 = (1'h0); (forvar3691 < (1'h1)); forvar3691 = (forvar3691 + (1'h1)))
                    begin
                      reg3692 <= $unsigned(reg3678[(3'h4):(2'h2)]);
                      reg3693 <= $unsigned((&$unsigned(reg3675[(2'h3):(2'h2)])));
                    end
                  if ((~{reg67[(1'h0):(1'h0)]}))
                    begin
                      reg3694 <= ((reg83[(2'h3):(2'h3)] >>> $unsigned($unsigned(reg32))) <= (reg27 ?
                          (|$signed(reg3690)) : $unsigned(reg49)));
                      reg3695 <= (wire5 ?
                          $unsigned(reg28[(4'hb):(4'hb)]) : (^$signed(reg40)));
                      reg3696 <= ({(~^(reg17 ? wire3634 : (8'hb1)))} ?
                          (^~$unsigned(reg3672)) : {$signed((reg3650 ?
                                  reg63 : reg31))});
                      reg3697 <= ({(~(8'h9e))} ?
                          (!reg14) : ((^~(forvar3676 & reg16)) ?
                              (~$unsigned(forvar3664)) : ((reg13 ?
                                  reg77 : reg31) ^ reg76)));
                    end
                  else
                    begin
                      reg3694 <= {$signed($unsigned((|reg80)))};
                    end
                  if ($unsigned(((8'haf) ?
                      (wire8 ?
                          $signed((8'ha0)) : ((8'hb7) ?
                              reg70 : (8'ha8))) : $unsigned($unsigned(reg3655)))))
                    begin
                      reg3698 <= $signed($signed((~^(^reg24))));
                      reg3699 <= ((reg3665 ~^ forvar3655[(3'h7):(3'h6)]) ?
                          (8'ha7) : (!(!(~&wire85))));
                    end
                  else
                    begin
                      reg3698 <= ($unsigned(reg3656[(1'h1):(1'h1)]) | {((reg83 - wire85) ?
                              reg3669[(3'h5):(3'h5)] : reg77)});
                      reg3699 <= reg34;
                      reg3700 <= wire3636;
                      reg3701 <= reg3673;
                    end
                  if ({$unsigned(forvar3639)})
                    begin
                      reg3702 <= $signed((^(8'hb0)));
                      reg3703 <= reg70[(1'h1):(1'h1)];
                      reg3704 <= (8'ha7);
                      reg3705 <= reg43;
                    end
                  else
                    begin
                      reg3702 <= reg3673[(3'h5):(3'h4)];
                      reg3703 <= (~{reg84[(1'h0):(1'h0)]});
                      reg3704 <= $unsigned((reg3702[(4'h8):(4'h8)] >> ((^~reg33) <<< {(8'hab)})));
                    end
                end
              else
                begin
                  for (forvar3691 = (1'h0); (forvar3691 < (2'h2)); forvar3691 = (forvar3691 + (1'h1)))
                    begin
                      reg3692 <= reg37[(2'h2):(2'h2)];
                      reg3693 <= $unsigned(((~&(reg3683 >> reg3678)) != (^~$signed(reg3697))));
                    end
                  for (forvar3694 = (1'h0); (forvar3694 < (2'h3)); forvar3694 = (forvar3694 + (1'h1)))
                    begin
                      reg3695 <= reg74[(3'h4):(2'h2)];
                      reg3696 <= ((({(8'h9d)} ?
                              reg48 : (reg3652 ?
                                  forvar3663 : reg3645)) || ($signed(reg3679) | reg12)) ?
                          reg3660 : $signed({reg3659}));
                      reg3697 <= $signed(reg3649);
                    end
                  reg3698 <= (((8'ha8) ^~ ((reg3641 << reg3694) + reg54[(2'h2):(1'h1)])) ?
                      {((~&wire3634) << (reg3672 ^~ reg63))} : reg48);
                  for (forvar3699 = (1'h0); (forvar3699 < (1'h0)); forvar3699 = (forvar3699 + (1'h1)))
                    begin
                      reg3700 <= reg60;
                      reg3701 <= ((reg22 & {wire8[(1'h1):(1'h1)]}) < (((forvar3648 ^~ reg27) ?
                          $signed(reg48) : (reg3685 ?
                              reg61 : wire3634)) ^~ (~$unsigned(forvar3683))));
                      reg3702 <= ((~|$unsigned($signed(reg3699))) - $signed(((reg75 * reg36) << (~|wire3632))));
                    end
                end
              reg3706 <= reg79;
              for (forvar3707 = (1'h0); (forvar3707 < (1'h0)); forvar3707 = (forvar3707 + (1'h1)))
                begin
                  for (forvar3708 = (1'h0); (forvar3708 < (2'h2)); forvar3708 = (forvar3708 + (1'h1)))
                    begin
                      reg3709 <= ($signed(((~(8'ha7)) ?
                          reg31 : $signed(reg3666))) && reg3687);
                      reg3710 <= (!$unsigned($unsigned((-reg3692))));
                    end
                  for (forvar3711 = (1'h0); (forvar3711 < (1'h1)); forvar3711 = (forvar3711 + (1'h1)))
                    begin
                      reg3712 <= $signed({(reg3658 - (~^reg3702))});
                      reg3713 <= $unsigned(((|((8'ha8) | (8'ha2))) ?
                          forvar3638[(3'h4):(1'h0)] : ({reg56} <<< $unsigned(reg3642))));
                      reg3714 <= $unsigned($unsigned($unsigned(((8'ha6) ^~ reg3709))));
                    end
                  if ((|($signed((reg3700 ^~ (8'hb7))) != $unsigned((reg3667 & (8'h9d))))))
                    begin
                      reg3715 <= (^{(~(~(8'h9d)))});
                      reg3716 <= $signed((~|$signed(reg3702[(3'h4):(1'h1)])));
                      reg3717 <= forvar3708;
                      reg3718 <= (~&((~&(!(8'haf))) ?
                          $unsigned($signed(reg3653)) : reg19));
                    end
                  else
                    begin
                      reg3715 <= $signed(reg3714[(2'h2):(1'h0)]);
                      reg3716 <= ($unsigned((^((8'hba) ? reg3643 : reg3693))) ?
                          ((&reg3661) == ($signed(reg73) != {reg33})) : (+$signed((reg51 + reg67))));
                      reg3717 <= $unsigned(({$unsigned(reg3648)} ?
                          $signed($unsigned(reg18)) : (+reg32)));
                    end
                  reg3719 <= (8'ha1);
                end
            end
          else
            begin
              for (forvar3680 = (1'h0); (forvar3680 < (1'h1)); forvar3680 = (forvar3680 + (1'h1)))
                begin
                  if (reg3687)
                    begin
                      reg3681 <= (~{$signed(reg3687[(4'hd):(1'h1)])});
                      reg3682 <= reg3717[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg3681 <= forvar3676;
                    end
                end
              reg3683 <= ((forvar3694[(2'h2):(1'h0)] ~^ ($signed(reg16) ?
                  {forvar3663} : reg3688[(2'h2):(1'h0)])) | (^~{(~&reg3637)}));
              reg3684 <= ($signed(((&forvar3664) << (reg3675 ?
                      reg3697 : reg52))) ?
                  $unsigned({$unsigned(reg3675)}) : (|$unsigned($signed(wire8))));
              if ($unsigned(($signed($signed((8'hb9))) >> (8'ha6))))
                begin
                  for (forvar3685 = (1'h0); (forvar3685 < (1'h0)); forvar3685 = (forvar3685 + (1'h1)))
                    begin
                      reg3686 <= {(8'hb8)};
                      reg3687 <= $signed((reg73 <= (-$signed(reg19))));
                      reg3688 <= (^(reg54 & reg3693));
                      reg3689 <= (8'hae);
                    end
                  if (reg3698)
                    begin
                      reg3690 <= reg3666[(1'h1):(1'h0)];
                      reg3691 <= $unsigned(forvar3699[(1'h1):(1'h1)]);
                      reg3692 <= (~reg3674[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg3690 <= $unsigned(reg3710);
                      reg3691 <= reg3694[(2'h3):(1'h1)];
                    end
                  for (forvar3693 = (1'h0); (forvar3693 < (2'h2)); forvar3693 = (forvar3693 + (1'h1)))
                    begin
                      reg3694 <= reg21[(1'h0):(1'h0)];
                      reg3695 <= forvar3656;
                    end
                  if (($signed({{reg3656}}) << reg59))
                    begin
                      reg3696 <= ($unsigned(reg54) ? reg48 : $signed(wire8));
                      reg3697 <= (reg24 ?
                          (reg3689 <<< $unsigned((reg26 && reg43))) : reg32);
                    end
                  else
                    begin
                      reg3696 <= $unsigned(reg13);
                      reg3697 <= {{$signed((~|reg3679))}};
                      reg3698 <= ({(|(^~reg3712))} ?
                          $signed(wire3636) : reg3714);
                    end
                end
              else
                begin
                  if ((forvar3708 ^ $unsigned(($signed(reg3647) < {forvar3671}))))
                    begin
                      reg3685 <= (8'ha5);
                      reg3686 <= (forvar3651 || (((8'hb9) + $signed(forvar3638)) << (8'hb3)));
                      reg3687 <= (|(((reg24 && reg3683) ^ reg3682) ?
                          (^~(reg3695 ?
                              reg33 : reg3646)) : $signed(forvar3680)));
                      reg3688 <= $unsigned($unsigned($signed((~|reg57))));
                    end
                  else
                    begin
                      reg3685 <= $unsigned((|{forvar3649[(3'h6):(3'h5)]}));
                      reg3686 <= (((~|$unsigned(wire3632)) <<< (~$unsigned(reg76))) ?
                          $signed(((&reg3655) ?
                              (reg75 ?
                                  reg3698 : reg79) : reg3654)) : {(!$signed(reg3669))});
                      reg3687 <= (~&({((8'h9f) >>> reg3657)} ?
                          reg3650 : $unsigned(((8'hb0) < wire3636))));
                    end
                end
            end
        end
    end
  assign wire3720 = reg70[(1'h1):(1'h0)];
  assign wire3721 = $unsigned((reg3673 >> $signed($unsigned(wire3720))));
  always
    @(posedge clk) begin
      if ($unsigned(((reg3673[(2'h3):(1'h1)] >= (reg3701 ? (8'haf) : reg3694)) ?
          $signed(reg3640) : reg73[(1'h0):(1'h0)])))
        begin
          if ($signed(reg32))
            begin
              reg3722 <= reg3679;
              reg3723 <= ($unsigned(wire6[(4'h9):(1'h1)]) + $signed(reg54[(3'h7):(1'h1)]));
              reg3724 <= reg49;
              if (reg10[(3'h6):(3'h4)])
                begin
                  for (forvar3725 = (1'h0); (forvar3725 < (1'h1)); forvar3725 = (forvar3725 + (1'h1)))
                    begin
                      reg3726 <= (reg75 >> reg3656);
                      reg3727 <= (reg72 != $unsigned((-$unsigned((8'ha1)))));
                      reg3728 <= (reg3687 > (~&($signed(reg3690) ?
                          wire7 : {reg53})));
                      reg3729 <= ($unsigned($unsigned($signed(reg3696))) ?
                          reg3658 : (8'ha7));
                    end
                  reg3730 <= $unsigned($unsigned($unsigned($unsigned(reg51))));
                  for (forvar3731 = (1'h0); (forvar3731 < (1'h0)); forvar3731 = (forvar3731 + (1'h1)))
                    begin
                      reg3732 <= $signed($unsigned($unsigned((reg46 ?
                          reg54 : reg50))));
                      reg3733 <= (~&reg3649[(3'h4):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar3725 = (1'h0); (forvar3725 < (1'h1)); forvar3725 = (forvar3725 + (1'h1)))
                    begin
                      reg3726 <= reg21[(1'h0):(1'h0)];
                      reg3727 <= reg3646[(4'he):(3'h4)];
                      reg3728 <= reg46;
                    end
                  for (forvar3729 = (1'h0); (forvar3729 < (2'h2)); forvar3729 = (forvar3729 + (1'h1)))
                    begin
                      reg3730 <= {reg61[(1'h1):(1'h0)]};
                      reg3731 <= reg3640[(1'h0):(1'h0)];
                    end
                  for (forvar3732 = (1'h0); (forvar3732 < (2'h2)); forvar3732 = (forvar3732 + (1'h1)))
                    begin
                      reg3733 <= ((+$signed(reg3655)) >> $unsigned((8'ha1)));
                      reg3734 <= $signed($unsigned(reg64));
                      reg3735 <= $unsigned(reg3651);
                    end
                  if ($unsigned(($signed($unsigned(reg3656)) ?
                      {$signed(reg3695)} : ($unsigned(reg3735) << {reg3683}))))
                    begin
                      reg3736 <= ((($signed(reg13) ? reg76 : $unsigned(reg59)) ?
                              reg73[(3'h4):(1'h1)] : {$signed(reg3724)}) ?
                          (($signed(reg3715) && $signed(reg25)) || ((reg51 ?
                                  (8'hb0) : reg3668) ?
                              (!reg76) : (~^reg34))) : reg15[(3'h7):(1'h0)]);
                      reg3737 <= ((-reg12[(1'h0):(1'h0)]) - wire3634[(2'h3):(2'h3)]);
                      reg3738 <= {reg43};
                      reg3739 <= reg3662;
                    end
                  else
                    begin
                      reg3736 <= $unsigned(reg3653[(4'he):(4'he)]);
                      reg3737 <= reg16;
                      reg3738 <= $signed($signed($unsigned((~^reg47))));
                    end
                end
            end
          else
            begin
              reg3722 <= $signed($unsigned($signed((-(8'h9d)))));
              for (forvar3723 = (1'h0); (forvar3723 < (2'h2)); forvar3723 = (forvar3723 + (1'h1)))
                begin
                  for (forvar3724 = (1'h0); (forvar3724 < (1'h0)); forvar3724 = (forvar3724 + (1'h1)))
                    begin
                      reg3725 <= (8'hb2);
                      reg3726 <= $signed((8'ha6));
                      reg3727 <= $signed((($signed(reg3647) >> (|reg3718)) >>> $signed((^~reg77))));
                    end
                  for (forvar3728 = (1'h0); (forvar3728 < (1'h1)); forvar3728 = (forvar3728 + (1'h1)))
                    begin
                      reg3729 <= ($signed($signed($unsigned(reg84))) != ((8'hab) ?
                          $unsigned((reg74 ?
                              (8'ha0) : reg3726)) : (~^$signed(wire7))));
                      reg3730 <= (~reg3694[(3'h5):(2'h3)]);
                      reg3731 <= $signed(reg77[(4'ha):(3'h7)]);
                      reg3732 <= $signed($signed(($unsigned((8'ha9)) << $unsigned(reg3718))));
                    end
                  for (forvar3733 = (1'h0); (forvar3733 < (2'h3)); forvar3733 = (forvar3733 + (1'h1)))
                    begin
                      reg3734 <= ((+($unsigned((8'hba)) ?
                          reg3702 : (wire3720 ?
                              reg33 : (8'h9c)))) > reg3649[(2'h2):(1'h1)]);
                    end
                  for (forvar3735 = (1'h0); (forvar3735 < (2'h3)); forvar3735 = (forvar3735 + (1'h1)))
                    begin
                      reg3736 <= (reg3637[(3'h4):(2'h2)] ?
                          (reg3643[(3'h7):(3'h4)] ?
                              $signed((wire5 <= reg48)) : $unsigned((reg3670 ?
                                  (8'ha7) : reg53))) : reg3726);
                      reg3737 <= {($unsigned(reg3690) & (|(reg3710 != reg3647)))};
                      reg3738 <= (8'haf);
                      reg3739 <= (($unsigned((reg3716 ? reg49 : reg3661)) ?
                              (^~(reg3650 ?
                                  reg3646 : reg3739)) : $signed($signed(reg10))) ?
                          ((reg17[(4'h8):(1'h1)] ?
                                  (reg34 ?
                                      reg3732 : reg3736) : $unsigned(reg28)) ?
                              (&(+reg3719)) : (~&{reg3641})) : reg3653);
                    end
                end
              for (forvar3740 = (1'h0); (forvar3740 < (1'h0)); forvar3740 = (forvar3740 + (1'h1)))
                begin
                  for (forvar3741 = (1'h0); (forvar3741 < (2'h2)); forvar3741 = (forvar3741 + (1'h1)))
                    begin
                      reg3742 <= $signed({{(8'h9f)}});
                    end
                end
            end
          reg3743 <= reg15[(1'h0):(1'h0)];
          for (forvar3744 = (1'h0); (forvar3744 < (2'h2)); forvar3744 = (forvar3744 + (1'h1)))
            begin
              reg3745 <= reg49[(1'h1):(1'h1)];
              if ((8'ha2))
                begin
                  reg3746 <= {$unsigned($signed($signed((8'hb3))))};
                  if (($signed(reg3728) || reg63[(2'h2):(1'h0)]))
                    begin
                      reg3747 <= ((reg3691 ?
                          (^~$signed((8'hba))) : (~^((8'hb1) ?
                              reg3746 : (8'hb0)))) == ({$unsigned(reg60)} ?
                          $unsigned((reg54 | reg3666)) : reg3696));
                      reg3748 <= reg3637;
                      reg3749 <= $signed(wire3720);
                      reg3750 <= reg3709[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg3747 <= $signed($signed({$unsigned(reg3695)}));
                    end
                end
              else
                begin
                  if ((-{((reg3660 && reg27) <<< $unsigned((8'hb9)))}))
                    begin
                      reg3746 <= (~^($signed($unsigned(reg21)) ?
                          (reg3665[(3'h6):(2'h2)] <<< (forvar3731 ~^ reg3648)) : ($unsigned((8'ha7)) < $unsigned(reg3695))));
                      reg3747 <= $unsigned((reg3743 >= $unsigned($unsigned(reg37))));
                      reg3748 <= reg3714[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3746 <= $signed(reg20[(3'h4):(1'h0)]);
                      reg3747 <= $unsigned(($signed(reg3672[(3'h4):(3'h4)]) ?
                          reg59[(4'hb):(3'h6)] : ($signed(reg3688) ?
                              (reg3643 ? reg3717 : forvar3744) : (^reg3746))));
                      reg3748 <= reg33;
                      reg3749 <= (^~$signed($signed({reg3649})));
                    end
                  if (reg3704[(3'h5):(1'h1)])
                    begin
                      reg3750 <= (8'h9e);
                      reg3751 <= ((((reg3737 ?
                          reg3739 : forvar3729) << $unsigned(reg3746)) << ((reg3749 <= reg3699) ?
                          $signed(reg3726) : reg10)) - (^($signed(reg3738) & (reg3735 ^ forvar3725))));
                      reg3752 <= (reg3646 >> (reg80[(2'h2):(1'h0)] ?
                          reg3705 : reg40[(3'h5):(1'h0)]));
                      reg3753 <= {reg3645};
                    end
                  else
                    begin
                      reg3750 <= reg59[(4'hd):(1'h1)];
                      reg3751 <= (!reg3653[(3'h7):(1'h1)]);
                      reg3752 <= reg22;
                    end
                  for (forvar3754 = (1'h0); (forvar3754 < (1'h1)); forvar3754 = (forvar3754 + (1'h1)))
                    begin
                      reg3755 <= $signed($signed(((8'hb4) ?
                          (forvar3725 - reg3726) : (&reg3645))));
                      reg3756 <= (-($signed(reg3667) && (&reg49[(3'h7):(1'h0)])));
                      reg3757 <= (&$signed(reg80[(2'h2):(1'h0)]));
                      reg3758 <= ($signed($unsigned(reg68[(3'h6):(1'h0)])) ?
                          {$unsigned($signed(reg3745))} : reg20[(1'h0):(1'h0)]);
                    end
                end
            end
          for (forvar3759 = (1'h0); (forvar3759 < (1'h0)); forvar3759 = (forvar3759 + (1'h1)))
            begin
              for (forvar3760 = (1'h0); (forvar3760 < (2'h3)); forvar3760 = (forvar3760 + (1'h1)))
                begin
                  reg3761 <= $unsigned($signed($signed((!(8'ha7)))));
                  for (forvar3762 = (1'h0); (forvar3762 < (2'h2)); forvar3762 = (forvar3762 + (1'h1)))
                    begin
                      reg3763 <= (({reg71} ?
                              (reg3719 ? reg45 : (8'h9d)) : (+{reg3702})) ?
                          (8'hb1) : $signed(reg3647[(3'h4):(1'h1)]));
                      reg3764 <= {reg3661[(1'h0):(1'h0)]};
                    end
                  for (forvar3765 = (1'h0); (forvar3765 < (1'h0)); forvar3765 = (forvar3765 + (1'h1)))
                    begin
                      reg3766 <= (~^(reg3687 ?
                          (~|(reg3734 <<< reg3714)) : (~|(reg3665 ?
                              reg3652 : (8'h9c)))));
                      reg3767 <= reg3757;
                      reg3768 <= reg3696;
                      reg3769 <= $unsigned(reg3748[(2'h3):(2'h3)]);
                    end
                  for (forvar3770 = (1'h0); (forvar3770 < (2'h2)); forvar3770 = (forvar3770 + (1'h1)))
                    begin
                      reg3771 <= reg3767;
                      reg3772 <= reg27[(4'h8):(1'h0)];
                      reg3773 <= (((reg37 ?
                              (reg3766 ?
                                  (8'ha1) : reg12) : $signed((8'hb8))) - ((reg3660 ?
                              reg3753 : (8'hb7)) >> {reg3769})) ?
                          $unsigned($signed((|reg22))) : reg79[(2'h3):(2'h3)]);
                    end
                end
              for (forvar3774 = (1'h0); (forvar3774 < (1'h1)); forvar3774 = (forvar3774 + (1'h1)))
                begin
                  if (reg3643[(4'hc):(2'h2)])
                    begin
                      reg3775 <= (^~$signed(($signed(forvar3765) ?
                          reg3749 : reg3725)));
                      reg3776 <= ($unsigned(($signed(reg27) | (reg3756 ?
                          reg3694 : reg57))) == reg3728);
                      reg3777 <= (reg3692[(3'h4):(1'h1)] ?
                          ((((8'hb6) == reg3768) && $unsigned(reg3683)) <= ($unsigned(reg3683) ?
                              $unsigned(wire3634) : $unsigned(wire6))) : reg24[(4'hb):(4'ha)]);
                      reg3778 <= ($unsigned({$signed(reg73)}) ?
                          (-reg3642[(3'h6):(2'h2)]) : reg3685);
                    end
                  else
                    begin
                      reg3775 <= reg37;
                      reg3776 <= (reg3757 ?
                          {reg13[(3'h7):(3'h4)]} : $unsigned(reg53[(3'h5):(2'h3)]));
                      reg3777 <= $signed((~&({reg13} && (reg27 ?
                          (8'haf) : (8'haf)))));
                    end
                  reg3779 <= (8'ha2);
                  for (forvar3780 = (1'h0); (forvar3780 < (1'h1)); forvar3780 = (forvar3780 + (1'h1)))
                    begin
                      reg3781 <= ($unsigned(reg56) ~^ reg3733[(3'h7):(1'h1)]);
                    end
                end
              for (forvar3782 = (1'h0); (forvar3782 < (2'h3)); forvar3782 = (forvar3782 + (1'h1)))
                begin
                  for (forvar3783 = (1'h0); (forvar3783 < (2'h2)); forvar3783 = (forvar3783 + (1'h1)))
                    begin
                      reg3784 <= ({$unsigned((forvar3774 ?
                              (8'hb4) : reg3777))} << ((reg3669 <= (reg51 + reg3761)) == ({reg83} ?
                          $unsigned(reg15) : (reg3732 ? reg84 : reg3750))));
                    end
                  if (reg3756)
                    begin
                      reg3785 <= (((reg60 || {(8'hac)}) - $signed((reg3642 >= reg61))) | $signed($unsigned(reg3749[(1'h1):(1'h0)])));
                      reg3786 <= ($signed((8'ha4)) ?
                          (|reg68[(1'h1):(1'h0)]) : $signed((reg60 ^~ (reg17 || reg3746))));
                      reg3787 <= reg3669[(2'h3):(1'h0)];
                      reg3788 <= (^((8'hba) + (+$unsigned(reg3679))));
                    end
                  else
                    begin
                      reg3785 <= (((~reg73[(1'h1):(1'h0)]) + reg3644) ?
                          $unsigned(forvar3735[(3'h4):(2'h2)]) : $signed(((&reg3729) ?
                              reg3648 : (~^reg3771))));
                      reg3786 <= $signed((reg3660[(2'h3):(1'h1)] != (8'ha1)));
                    end
                  for (forvar3789 = (1'h0); (forvar3789 < (2'h2)); forvar3789 = (forvar3789 + (1'h1)))
                    begin
                      reg3790 <= $signed(reg3764);
                    end
                end
              reg3791 <= $signed({wire7[(3'h5):(2'h2)]});
            end
        end
      else
        begin
          for (forvar3722 = (1'h0); (forvar3722 < (2'h3)); forvar3722 = (forvar3722 + (1'h1)))
            begin
              for (forvar3723 = (1'h0); (forvar3723 < (2'h2)); forvar3723 = (forvar3723 + (1'h1)))
                begin
                  for (forvar3724 = (1'h0); (forvar3724 < (1'h0)); forvar3724 = (forvar3724 + (1'h1)))
                    begin
                      reg3725 <= (^$signed(((&reg3784) ?
                          (reg81 ? reg3738 : (8'hb1)) : (reg32 ^ reg48))));
                    end
                end
              reg3726 <= (^$signed(reg3660[(3'h4):(1'h1)]));
              for (forvar3727 = (1'h0); (forvar3727 < (2'h3)); forvar3727 = (forvar3727 + (1'h1)))
                begin
                  if ($unsigned(({(!reg83)} ?
                      {reg3692} : reg69[(2'h2):(1'h0)])))
                    begin
                      reg3728 <= reg31[(4'ha):(1'h1)];
                      reg3729 <= ((!(reg3723[(4'hc):(1'h1)] > {reg3729})) - (reg3668 ?
                          $signed((8'h9c)) : $unsigned((reg3639 ?
                              reg3763 : wire6))));
                    end
                  else
                    begin
                      reg3728 <= ({(reg25 ^~ (&reg81))} + ({{reg3752}} | reg3772));
                    end
                  for (forvar3730 = (1'h0); (forvar3730 < (2'h2)); forvar3730 = (forvar3730 + (1'h1)))
                    begin
                      reg3731 <= (reg61[(2'h3):(1'h0)] || (forvar3727[(1'h0):(1'h0)] && $signed($signed(reg18))));
                    end
                  reg3732 <= (&$signed((~|{forvar3730})));
                  if ((^~$unsigned(reg3709)))
                    begin
                      reg3733 <= $unsigned(((reg3712[(3'h5):(2'h3)] ?
                              $unsigned(reg12) : reg3735) ?
                          $unsigned(reg3650[(2'h2):(2'h2)]) : reg3696));
                    end
                  else
                    begin
                      reg3733 <= $unsigned(reg3704);
                      reg3734 <= (reg26[(1'h1):(1'h1)] < (~$unsigned((~|wire5))));
                    end
                end
              reg3735 <= $unsigned((~^wire3632[(3'h7):(1'h0)]));
            end
        end
      for (forvar3792 = (1'h0); (forvar3792 < (1'h0)); forvar3792 = (forvar3792 + (1'h1)))
        begin
          if ($signed((forvar3770 ? reg22 : {reg3756[(1'h0):(1'h0)]})))
            begin
              for (forvar3793 = (1'h0); (forvar3793 < (2'h2)); forvar3793 = (forvar3793 + (1'h1)))
                begin
                  if ($unsigned(reg3786[(3'h7):(2'h2)]))
                    begin
                      reg3794 <= {reg3652};
                      reg3795 <= forvar3780[(4'hd):(4'ha)];
                      reg3796 <= (!forvar3729[(3'h6):(3'h6)]);
                    end
                  else
                    begin
                      reg3794 <= (-(({wire85} ?
                          (&reg3649) : reg3737) >= ((-reg3773) ?
                          (forvar3782 ? forvar3759 : reg3784) : {reg77})));
                      reg3795 <= $signed(reg59);
                      reg3796 <= {$signed($unsigned(reg3757))};
                    end
                  for (forvar3797 = (1'h0); (forvar3797 < (2'h3)); forvar3797 = (forvar3797 + (1'h1)))
                    begin
                      reg3798 <= reg3679;
                    end
                end
              for (forvar3799 = (1'h0); (forvar3799 < (1'h0)); forvar3799 = (forvar3799 + (1'h1)))
                begin
                  reg3800 <= $signed(reg20);
                end
              for (forvar3801 = (1'h0); (forvar3801 < (2'h2)); forvar3801 = (forvar3801 + (1'h1)))
                begin
                  for (forvar3802 = (1'h0); (forvar3802 < (1'h1)); forvar3802 = (forvar3802 + (1'h1)))
                    begin
                      reg3803 <= (!reg28[(4'h8):(4'h8)]);
                      reg3804 <= reg3735[(2'h2):(2'h2)];
                      reg3805 <= {reg46[(1'h1):(1'h0)]};
                    end
                  if ((((reg3736[(2'h3):(2'h2)] ?
                      (reg74 ?
                          reg3749 : reg3637) : reg3709) == $signed($signed(reg3665))) != reg18))
                    begin
                      reg3806 <= (-(-$signed($unsigned(reg3768))));
                      reg3807 <= $unsigned($unsigned(wire3632[(3'h7):(3'h5)]));
                      reg3808 <= (reg3736[(4'h8):(4'h8)] <<< $signed(((forvar3724 <<< reg3692) ?
                          $signed(wire8) : reg34)));
                      reg3809 <= reg3644[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3806 <= forvar3783[(3'h6):(1'h0)];
                      reg3807 <= (forvar3801[(3'h4):(1'h1)] ?
                          (-{{reg31}}) : $signed((|(reg3667 - (8'hb3)))));
                      reg3808 <= ((!(!reg3657)) == $unsigned((8'had)));
                    end
                  for (forvar3810 = (1'h0); (forvar3810 < (2'h3)); forvar3810 = (forvar3810 + (1'h1)))
                    begin
                      reg3811 <= reg67[(1'h0):(1'h0)];
                      reg3812 <= $signed(forvar3724);
                      reg3813 <= $signed($unsigned({$unsigned(reg50)}));
                      reg3814 <= (~&(reg3804[(3'h4):(3'h4)] != $unsigned(((8'hb8) < reg3728))));
                    end
                  if (((8'h9d) >> ((8'ha5) ?
                      (&$signed((8'ha8))) : $signed(reg3692[(3'h4):(2'h2)]))))
                    begin
                      reg3815 <= $unsigned((+$unsigned($signed(forvar3793))));
                      reg3816 <= reg3651;
                      reg3817 <= (~^$signed(reg14[(1'h1):(1'h1)]));
                      reg3818 <= {$unsigned({(^~reg3738)})};
                    end
                  else
                    begin
                      reg3815 <= (^~$signed(((~|(8'haa)) && (wire5 - reg3731))));
                      reg3816 <= (-reg26[(1'h0):(1'h0)]);
                    end
                end
            end
          else
            begin
              for (forvar3793 = (1'h0); (forvar3793 < (1'h1)); forvar3793 = (forvar3793 + (1'h1)))
                begin
                  for (forvar3794 = (1'h0); (forvar3794 < (2'h3)); forvar3794 = (forvar3794 + (1'h1)))
                    begin
                      reg3795 <= reg3803;
                      reg3796 <= $signed((forvar3794[(4'hc):(3'h4)] >= {(&wire8)}));
                      reg3797 <= (|(^$unsigned({reg3654})));
                      reg3798 <= $unsigned((-$unsigned(reg3771)));
                    end
                  if ((((~^$unsigned(forvar3810)) ?
                      ($unsigned(reg3779) ?
                          reg3733 : (forvar3760 ?
                              (8'hb3) : reg3786)) : (reg3709[(3'h4):(2'h3)] ?
                          $signed(reg43) : reg3813[(2'h2):(1'h0)])) * $signed($signed(reg3688))))
                    begin
                      reg3799 <= $unsigned(((forvar3735 ?
                              $unsigned(reg3696) : (reg3650 >> forvar3731)) ?
                          {$unsigned(reg3657)} : wire3720[(4'h8):(3'h7)]));
                      reg3800 <= $unsigned(((reg3799 < reg3731[(2'h3):(1'h0)]) ?
                          (8'h9c) : reg45[(4'h8):(2'h3)]));
                      reg3801 <= ((-$unsigned($signed(reg3713))) ?
                          ({reg3778} & reg3726) : $signed($signed((!reg3643))));
                    end
                  else
                    begin
                      reg3799 <= (~&(reg15 == ((forvar3793 ?
                          reg34 : reg3648) > $unsigned(forvar3725))));
                      reg3800 <= $unsigned({(^~reg3786[(3'h7):(1'h1)])});
                    end
                  if ({(^{reg77})})
                    begin
                      reg3802 <= {(((-(8'ha0)) == reg3693) ?
                              wire3720 : (!forvar3793[(3'h6):(2'h2)]))};
                      reg3803 <= (+{(+(8'h9d))});
                      reg3804 <= $signed(reg70[(2'h3):(1'h0)]);
                    end
                  else
                    begin
                      reg3802 <= ((reg28 ?
                              ($signed((8'hb7)) ?
                                  (8'ha1) : $signed((8'ha3))) : {(&reg80)}) ?
                          reg18 : reg18);
                    end
                  reg3805 <= reg3734[(1'h1):(1'h0)];
                end
              if ($unsigned($signed((^(~|reg3712)))))
                begin
                  for (forvar3806 = (1'h0); (forvar3806 < (1'h0)); forvar3806 = (forvar3806 + (1'h1)))
                    begin
                      reg3807 <= (~reg3723);
                    end
                end
              else
                begin
                  if ((-(8'hb5)))
                    begin
                      reg3806 <= reg3775;
                      reg3807 <= reg3757;
                      reg3808 <= reg3814;
                      reg3809 <= (~&reg3737);
                    end
                  else
                    begin
                      reg3806 <= (-(~|((^reg3689) ? (&wire3721) : (+reg3658))));
                      reg3807 <= {$signed($unsigned((~&reg46)))};
                      reg3808 <= (reg69 ?
                          (((reg26 != reg10) ?
                              (+reg3727) : $unsigned(reg73)) < (reg3756[(2'h2):(1'h1)] ?
                              {reg3777} : (reg3800 ?
                                  forvar3723 : (8'h9f)))) : reg3785);
                      reg3809 <= $unsigned((~&$unsigned(reg77)));
                    end
                  reg3810 <= (~(|{forvar3722[(3'h4):(1'h1)]}));
                end
            end
          for (forvar3819 = (1'h0); (forvar3819 < (1'h0)); forvar3819 = (forvar3819 + (1'h1)))
            begin
              for (forvar3820 = (1'h0); (forvar3820 < (1'h0)); forvar3820 = (forvar3820 + (1'h1)))
                begin
                  for (forvar3821 = (1'h0); (forvar3821 < (1'h1)); forvar3821 = (forvar3821 + (1'h1)))
                    begin
                      reg3822 <= ((+((reg47 ?
                              reg3653 : wire3632) >= $unsigned(reg13))) ?
                          {$signed((~|reg3745))} : reg3811[(4'h8):(3'h5)]);
                    end
                  if (reg43[(2'h3):(1'h1)])
                    begin
                      reg3823 <= $signed(((~&(^~reg3773)) ?
                          $unsigned($signed((8'hba))) : wire3720));
                      reg3824 <= $unsigned($signed($signed(reg79[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg3823 <= $unsigned($unsigned((^(forvar3732 + (8'hab)))));
                      reg3824 <= ($signed($unsigned($unsigned(reg3699))) ?
                          reg3702[(3'h6):(3'h6)] : $unsigned({$signed(reg3736)}));
                      reg3825 <= (!$unsigned((8'ha7)));
                    end
                  if ((((!(+reg54)) ?
                          (!(8'ha9)) : ($unsigned(reg3758) == (reg54 ~^ (8'haf)))) ?
                      {$signed(reg3771)} : {{reg3732[(4'hb):(4'hb)]}}))
                    begin
                      reg3826 <= $unsigned($unsigned((~&$signed(reg3733))));
                      reg3827 <= forvar3723;
                      reg3828 <= $unsigned($signed((8'haa)));
                    end
                  else
                    begin
                      reg3826 <= {{$unsigned((8'ha0))}};
                      reg3827 <= reg45;
                      reg3828 <= (8'hb0);
                      reg3829 <= reg3719;
                    end
                  reg3830 <= reg3771;
                end
              if (reg3757)
                begin
                  for (forvar3831 = (1'h0); (forvar3831 < (2'h3)); forvar3831 = (forvar3831 + (1'h1)))
                    begin
                      reg3832 <= (^~($signed((~^reg28)) ?
                          ((reg3652 ?
                              reg25 : (8'hae)) >= wire3634[(2'h3):(1'h1)]) : forvar3731));
                      reg3833 <= reg16;
                      reg3834 <= reg3734;
                      reg3835 <= $unsigned((((wire3720 ?
                          reg43 : reg3706) - $signed(reg3803)) < reg3803));
                    end
                end
              else
                begin
                  for (forvar3831 = (1'h0); (forvar3831 < (2'h3)); forvar3831 = (forvar3831 + (1'h1)))
                    begin
                      reg3832 <= (($signed($unsigned(forvar3783)) ^~ (|reg3690[(1'h0):(1'h0)])) ?
                          {$signed((~^reg3715))} : $signed($signed((8'haf))));
                    end
                  for (forvar3833 = (1'h0); (forvar3833 < (2'h3)); forvar3833 = (forvar3833 + (1'h1)))
                    begin
                      reg3834 <= (reg59[(4'hb):(3'h5)] + reg3735);
                      reg3835 <= (reg3784[(1'h0):(1'h0)] >> (~&reg3726));
                      reg3836 <= (({(^reg3667)} >>> reg3745) ?
                          (((!reg3715) ?
                                  (reg3728 > (8'ha4)) : (reg45 & forvar3789)) ?
                              $signed({reg3688}) : (((8'hb6) ?
                                      (8'h9e) : (8'hac)) ?
                                  $signed(reg3738) : (reg3641 ?
                                      reg20 : (8'hb0)))) : $unsigned((&$signed(reg3690))));
                      reg3837 <= ($unsigned(reg3667) != {(~(reg3705 ?
                              (8'haa) : reg3717))});
                    end
                end
            end
          for (forvar3838 = (1'h0); (forvar3838 < (2'h2)); forvar3838 = (forvar3838 + (1'h1)))
            begin
              if ($signed((^~$unsigned((|reg3776)))))
                begin
                  if ($unsigned($signed((reg75[(3'h4):(1'h1)] ~^ (reg3693 ?
                      reg3718 : reg3697)))))
                    begin
                      reg3839 <= ($unsigned((8'ha4)) ?
                          (((reg57 ? reg3761 : reg3826) ?
                              (~&reg3729) : $unsigned(reg3643)) >>> reg59) : (|(reg3703 * ((8'hb2) >> reg52))));
                      reg3840 <= ({$unsigned((8'ha3))} >> forvar3789);
                      reg3841 <= ($unsigned($signed((reg3812 ~^ reg3751))) == (~reg3660));
                    end
                  else
                    begin
                      reg3839 <= $unsigned((~^$signed((forvar3782 <<< (8'h9d)))));
                      reg3840 <= reg3836;
                    end
                  reg3842 <= forvar3838;
                  for (forvar3843 = (1'h0); (forvar3843 < (2'h3)); forvar3843 = (forvar3843 + (1'h1)))
                    begin
                      reg3844 <= reg3668;
                      reg3845 <= (~|((^(reg3822 ?
                          reg3732 : reg3658)) - reg3809));
                    end
                  reg3846 <= (($unsigned((8'hb8)) ?
                      ((reg25 ?
                          (8'ha6) : reg3652) >> (^~(8'hb6))) : reg54) ^~ (+($unsigned(reg56) ?
                      {reg3641} : (reg3835 - forvar3794))));
                end
              else
                begin
                  for (forvar3839 = (1'h0); (forvar3839 < (2'h2)); forvar3839 = (forvar3839 + (1'h1)))
                    begin
                      reg3840 <= (|reg3763[(1'h0):(1'h0)]);
                      reg3841 <= ((((8'ha9) ?
                          (forvar3797 ^ reg54) : $signed((8'ha2))) != (^~$unsigned((8'h9c)))) ^~ (!$unsigned(reg67[(4'h8):(4'h8)])));
                    end
                  for (forvar3842 = (1'h0); (forvar3842 < (1'h1)); forvar3842 = (forvar3842 + (1'h1)))
                    begin
                      reg3843 <= $signed($unsigned((~&{reg3749})));
                      reg3844 <= reg3685[(2'h3):(1'h1)];
                      reg3845 <= ((8'haa) ?
                          $signed($unsigned($unsigned(reg68))) : ((+(~&reg45)) * $signed(((8'hab) ?
                              reg72 : (8'hb1)))));
                    end
                  for (forvar3846 = (1'h0); (forvar3846 < (1'h0)); forvar3846 = (forvar3846 + (1'h1)))
                    begin
                      reg3847 <= $signed(reg3714[(2'h2):(2'h2)]);
                      reg3848 <= (reg3786[(3'h4):(2'h2)] <= $signed(reg3781));
                      reg3849 <= $unsigned($unsigned(reg3699));
                      reg3850 <= ($unsigned(reg3817) ^~ (!((reg3692 != reg3710) ?
                          (~&(8'ha0)) : reg83[(3'h5):(2'h2)])));
                    end
                end
              for (forvar3851 = (1'h0); (forvar3851 < (2'h2)); forvar3851 = (forvar3851 + (1'h1)))
                begin
                  if ({$unsigned($unsigned(reg3769[(3'h6):(2'h2)]))})
                    begin
                      reg3852 <= reg50[(4'ha):(3'h5)];
                    end
                  else
                    begin
                      reg3852 <= $unsigned(reg3639[(3'h4):(2'h3)]);
                      reg3853 <= (8'hb9);
                    end
                  reg3854 <= ({(8'had)} ?
                      $signed(forvar3730[(3'h4):(2'h2)]) : reg3648[(3'h6):(3'h5)]);
                  reg3855 <= (+$signed(forvar3762[(4'hd):(4'ha)]));
                end
              for (forvar3856 = (1'h0); (forvar3856 < (2'h2)); forvar3856 = (forvar3856 + (1'h1)))
                begin
                  if ((reg3850 + $unsigned($signed((reg46 ?
                      reg3781 : (8'hac))))))
                    begin
                      reg3857 <= ((~&{(^~reg3854)}) <= ({(forvar3735 < reg31)} ?
                          $unsigned($unsigned(reg3810)) : {reg3797[(2'h3):(2'h2)]}));
                      reg3858 <= {reg3825[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg3857 <= reg3669;
                    end
                end
            end
          if (((^~reg3798[(3'h6):(1'h0)]) - (reg27[(3'h6):(3'h5)] ^ $unsigned((~|reg3853)))))
            begin
              for (forvar3859 = (1'h0); (forvar3859 < (2'h2)); forvar3859 = (forvar3859 + (1'h1)))
                begin
                  if ($unsigned(((8'ha2) != {{reg15}})))
                    begin
                      reg3860 <= ((+forvar3774[(1'h1):(1'h1)]) | (~&(reg3787 ?
                          (reg3650 ?
                              reg3842 : reg3852) : forvar3838[(2'h3):(2'h3)])));
                    end
                  else
                    begin
                      reg3860 <= {reg3725};
                      reg3861 <= reg3652[(4'h8):(2'h2)];
                    end
                  for (forvar3862 = (1'h0); (forvar3862 < (1'h0)); forvar3862 = (forvar3862 + (1'h1)))
                    begin
                      reg3863 <= ((|$unsigned(((8'ha4) << reg50))) ?
                          ((&reg3681[(2'h3):(2'h2)]) | ({reg3662} >> {reg3826})) : ((~&$signed(reg3668)) ?
                              ($signed(forvar3831) ^~ reg15[(3'h4):(3'h4)]) : $unsigned(reg12[(3'h4):(3'h4)])));
                      reg3864 <= forvar3725;
                      reg3865 <= reg80;
                    end
                end
              reg3866 <= (forvar3789[(4'hc):(1'h0)] ?
                  ($signed((^(8'ha0))) >= reg3818[(1'h0):(1'h0)]) : reg45);
              reg3867 <= reg22;
            end
          else
            begin
              if ($signed(reg3639))
                begin
                  if (({reg3735[(2'h2):(2'h2)]} || reg3742))
                    begin
                      reg3859 <= $signed($signed($unsigned((reg84 ^~ reg3807))));
                    end
                  else
                    begin
                      reg3859 <= {$unsigned((reg53 ?
                              reg64[(2'h2):(1'h0)] : wire6[(3'h6):(1'h0)]))};
                      reg3860 <= reg3844[(4'hb):(2'h3)];
                      reg3861 <= $signed(((reg3827[(3'h6):(2'h2)] ?
                              ((8'h9d) >> (8'ha6)) : $unsigned(reg63)) ?
                          ((reg3771 ?
                              reg3655 : reg3742) - $signed(forvar3799)) : $signed(reg3839)));
                    end
                end
              else
                begin
                  if (($signed({(reg3727 <= reg3714)}) ?
                      $unsigned(reg81) : $signed((8'hb3))))
                    begin
                      reg3859 <= forvar3856;
                      reg3860 <= ($unsigned($unsigned(reg3670[(4'hb):(3'h7)])) >= {((reg61 < reg3643) && (reg3807 && reg3751))});
                    end
                  else
                    begin
                      reg3859 <= ($signed(($unsigned((8'hac)) ?
                          reg21[(3'h4):(1'h0)] : $unsigned(reg3666))) ^ forvar3780);
                      reg3860 <= ({(^$unsigned(reg3733))} ?
                          forvar3760 : {forvar3793});
                      reg3861 <= (~|$unsigned((~|reg3784)));
                    end
                  for (forvar3862 = (1'h0); (forvar3862 < (1'h0)); forvar3862 = (forvar3862 + (1'h1)))
                    begin
                      reg3863 <= (($unsigned({reg3675}) ?
                          (+{reg63}) : ((forvar3728 ?
                              reg3725 : (8'ha9)) >>> reg3738)) ^ {$unsigned($unsigned(reg20))});
                      reg3864 <= $signed({(!(reg3730 <= reg3701))});
                    end
                  for (forvar3865 = (1'h0); (forvar3865 < (2'h3)); forvar3865 = (forvar3865 + (1'h1)))
                    begin
                      reg3866 <= (~(($unsigned((8'hb6)) > $unsigned(reg70)) >>> $signed(wire85)));
                      reg3867 <= $signed({reg3700});
                      reg3868 <= (^~(-reg3662));
                      reg3869 <= ((8'hb7) >> $unsigned((~&(forvar3789 - forvar3740))));
                    end
                  for (forvar3870 = (1'h0); (forvar3870 < (1'h1)); forvar3870 = (forvar3870 + (1'h1)))
                    begin
                      reg3871 <= reg3763;
                      reg3872 <= ({$unsigned($unsigned(forvar3851))} == reg57[(1'h0):(1'h0)]);
                      reg3873 <= (&$unsigned(($unsigned(reg3679) != (~forvar3870))));
                    end
                end
              if ($unsigned(($signed(((8'ha7) ^~ (8'ha7))) ?
                  $unsigned((+(8'h9d))) : (reg3645 & $unsigned((8'ha3))))))
                begin
                  if ((~|{(^(reg3769 ? reg3745 : reg51))}))
                    begin
                      reg3874 <= reg3812;
                      reg3875 <= (+{$signed((!(8'hae)))});
                    end
                  else
                    begin
                      reg3874 <= {reg3786[(2'h3):(2'h3)]};
                      reg3875 <= (!reg3643[(3'h7):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar3874 = (1'h0); (forvar3874 < (2'h2)); forvar3874 = (forvar3874 + (1'h1)))
                    begin
                      reg3875 <= (!reg3718);
                      reg3876 <= $signed($signed(((reg3700 ^ reg3657) <<< reg3739[(2'h3):(1'h0)])));
                      reg3877 <= reg3717[(2'h2):(1'h1)];
                    end
                  if ((|(forvar3810 | ($unsigned(reg3855) ?
                      $signed(reg3848) : (reg3810 || reg3745)))))
                    begin
                      reg3878 <= reg3679[(3'h5):(2'h2)];
                      reg3879 <= $signed($unsigned(reg3794[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg3878 <= wire85[(3'h5):(1'h0)];
                      reg3879 <= ((!$unsigned(reg3844)) & reg3827[(2'h3):(2'h3)]);
                      reg3880 <= (({$signed(reg3644)} ?
                              forvar3831 : (!(forvar3870 ~^ reg3748))) ?
                          $signed((~reg3716)) : {(+(reg3758 ?
                                  reg3669 : (8'hb1)))});
                    end
                end
              for (forvar3881 = (1'h0); (forvar3881 < (1'h0)); forvar3881 = (forvar3881 + (1'h1)))
                begin
                  if ($signed((8'hb9)))
                    begin
                      reg3882 <= reg3643[(3'h4):(1'h1)];
                      reg3883 <= reg3761[(1'h0):(1'h0)];
                      reg3884 <= reg53;
                    end
                  else
                    begin
                      reg3882 <= wire85;
                      reg3883 <= forvar3729;
                    end
                end
            end
        end
      for (forvar3885 = (1'h0); (forvar3885 < (2'h3)); forvar3885 = (forvar3885 + (1'h1)))
        begin
          reg3886 <= $signed(({$signed(reg52)} ?
              $unsigned(reg3808[(2'h2):(1'h0)]) : ($signed(reg3843) ~^ (|reg3829))));
        end
      for (forvar3887 = (1'h0); (forvar3887 < (2'h2)); forvar3887 = (forvar3887 + (1'h1)))
        begin
          for (forvar3888 = (1'h0); (forvar3888 < (1'h1)); forvar3888 = (forvar3888 + (1'h1)))
            begin
              for (forvar3889 = (1'h0); (forvar3889 < (2'h2)); forvar3889 = (forvar3889 + (1'h1)))
                begin
                  for (forvar3890 = (1'h0); (forvar3890 < (1'h0)); forvar3890 = (forvar3890 + (1'h1)))
                    begin
                      reg3891 <= $unsigned((reg69 >> (((8'h9c) < reg3731) ^~ (reg3772 && reg56))));
                      reg3892 <= $unsigned((((reg3805 - reg3725) | (reg3771 - reg3877)) & (&{reg43})));
                    end
                  for (forvar3893 = (1'h0); (forvar3893 < (1'h0)); forvar3893 = (forvar3893 + (1'h1)))
                    begin
                      reg3894 <= $signed(reg3687);
                      reg3895 <= {$signed(reg14[(2'h3):(1'h0)])};
                    end
                  if ((~&(~&(forvar3722 << (reg14 >>> reg3840)))))
                    begin
                      reg3896 <= forvar3862;
                      reg3897 <= ({$unsigned(reg61)} ?
                          ((forvar3888 ?
                              $unsigned(reg19) : ((8'ha5) < wire6)) >> $signed((-forvar3865))) : ((|reg3643[(3'h5):(2'h2)]) | reg3696));
                      reg3898 <= $unsigned(reg3859[(4'h9):(4'h8)]);
                    end
                  else
                    begin
                      reg3896 <= ($unsigned(wire6) == (-reg57[(2'h3):(2'h3)]));
                      reg3897 <= reg3657[(1'h1):(1'h1)];
                      reg3898 <= (({reg3692} ?
                          $signed($unsigned(reg3892)) : reg28) ^~ (reg3804[(4'h8):(4'h8)] >>> $signed($unsigned(reg3709))));
                    end
                  reg3899 <= reg3678;
                end
              for (forvar3900 = (1'h0); (forvar3900 < (1'h0)); forvar3900 = (forvar3900 + (1'h1)))
                begin
                  for (forvar3901 = (1'h0); (forvar3901 < (1'h0)); forvar3901 = (forvar3901 + (1'h1)))
                    begin
                      reg3902 <= forvar3874[(3'h6):(2'h2)];
                      reg3903 <= $signed((^$unsigned((reg3652 ?
                          reg3745 : reg3791))));
                    end
                  for (forvar3904 = (1'h0); (forvar3904 < (1'h0)); forvar3904 = (forvar3904 + (1'h1)))
                    begin
                      reg3905 <= (((8'haf) <= $unsigned((~forvar3889))) ?
                          forvar3783[(4'hb):(4'h9)] : (~reg3884[(1'h1):(1'h1)]));
                    end
                  if ($unsigned(reg3651))
                    begin
                      reg3906 <= $unsigned(((+(reg3682 ^~ reg19)) >>> reg56));
                      reg3907 <= (+(forvar3799 * reg83));
                      reg3908 <= reg72;
                      reg3909 <= ($signed($unsigned(reg70)) > ($unsigned($signed(reg3876)) ?
                          forvar3725 : reg3860));
                    end
                  else
                    begin
                      reg3906 <= {$unsigned(reg3736[(3'h5):(3'h4)])};
                      reg3907 <= (reg3694 <<< (&$signed((reg15 != reg17))));
                    end
                end
            end
          for (forvar3910 = (1'h0); (forvar3910 < (2'h3)); forvar3910 = (forvar3910 + (1'h1)))
            begin
              if ((~|$unsigned((&(forvar3851 ? (8'hb2) : forvar3782)))))
                begin
                  for (forvar3911 = (1'h0); (forvar3911 < (2'h3)); forvar3911 = (forvar3911 + (1'h1)))
                    begin
                      reg3912 <= $unsigned((8'ha3));
                      reg3913 <= $signed($unsigned(($unsigned(reg3677) ?
                          reg3816[(3'h4):(2'h3)] : (8'ha3))));
                      reg3914 <= (reg3775[(4'h9):(2'h3)] ?
                          (reg3731[(2'h2):(1'h1)] && reg3908) : {forvar3821[(4'h8):(2'h3)]});
                    end
                  if ($unsigned(reg3758[(1'h1):(1'h1)]))
                    begin
                      reg3915 <= $signed(reg3877);
                      reg3916 <= ($unsigned($signed($unsigned(reg3795))) ?
                          $unsigned($signed(reg3656[(3'h7):(2'h3)])) : {reg3858[(3'h6):(2'h3)]});
                    end
                  else
                    begin
                      reg3915 <= ($signed(reg3813) <<< reg3646);
                      reg3916 <= reg46[(3'h4):(1'h1)];
                    end
                end
              else
                begin
                  if ({(~{forvar3889[(2'h3):(1'h0)]})})
                    begin
                      reg3911 <= $unsigned(reg3785[(2'h3):(2'h2)]);
                      reg3912 <= $unsigned(reg3678[(4'h8):(3'h6)]);
                      reg3913 <= {reg3700};
                      reg3914 <= reg3875;
                    end
                  else
                    begin
                      reg3911 <= (forvar3733 ?
                          $unsigned((^~$signed(reg3841))) : (~^$signed((reg14 ^~ forvar3842))));
                      reg3912 <= (($signed({forvar3810}) ~^ (8'ha5)) == reg3863);
                    end
                  if ($signed($unsigned((!$signed(reg3837)))))
                    begin
                      reg3915 <= reg3908;
                      reg3916 <= ((+$signed((8'hb7))) && (&((reg3826 ?
                          reg3898 : reg3697) ~^ $unsigned(forvar3838))));
                      reg3917 <= $unsigned((!reg3807));
                    end
                  else
                    begin
                      reg3915 <= $signed({{(^forvar3765)}});
                      reg3916 <= $unsigned(((8'haf) ?
                          reg3677[(3'h7):(3'h7)] : reg3656));
                      reg3917 <= (forvar3762[(4'h8):(3'h4)] <<< (reg3785 << reg3728[(1'h1):(1'h1)]));
                      reg3918 <= reg3828;
                    end
                end
            end
        end
    end
  assign wire3919 = reg3814[(2'h3):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar3920 = (1'h0); (forvar3920 < (2'h3)); forvar3920 = (forvar3920 + (1'h1)))
        begin
          for (forvar3921 = (1'h0); (forvar3921 < (2'h2)); forvar3921 = (forvar3921 + (1'h1)))
            begin
              for (forvar3922 = (1'h0); (forvar3922 < (2'h3)); forvar3922 = (forvar3922 + (1'h1)))
                begin
                  if ($unsigned((~&(&(~reg3710)))))
                    begin
                      reg3923 <= reg3651[(4'h8):(4'h8)];
                      reg3924 <= reg3781[(4'h8):(4'h8)];
                      reg3925 <= reg3723[(4'hb):(3'h6)];
                    end
                  else
                    begin
                      reg3923 <= $unsigned($unsigned({$signed((8'ha4))}));
                      reg3924 <= (reg3837 == reg3745);
                    end
                  for (forvar3926 = (1'h0); (forvar3926 < (1'h1)); forvar3926 = (forvar3926 + (1'h1)))
                    begin
                      reg3927 <= $signed((^$signed(reg3748[(4'h9):(3'h5)])));
                    end
                end
            end
          for (forvar3928 = (1'h0); (forvar3928 < (2'h3)); forvar3928 = (forvar3928 + (1'h1)))
            begin
              for (forvar3929 = (1'h0); (forvar3929 < (1'h0)); forvar3929 = (forvar3929 + (1'h1)))
                begin
                  for (forvar3930 = (1'h0); (forvar3930 < (2'h3)); forvar3930 = (forvar3930 + (1'h1)))
                    begin
                      reg3931 <= $unsigned(($signed(reg3913[(3'h7):(2'h3)]) ?
                          $unsigned(reg3731) : reg3817[(1'h1):(1'h0)]));
                      reg3932 <= (($unsigned($signed((8'had))) ?
                              reg54[(4'h8):(4'h8)] : (!{reg68})) ?
                          (($signed(reg3674) < reg3865) ?
                              reg24 : (reg3669[(3'h7):(3'h7)] >>> ((8'h9f) ?
                                  reg3727 : (8'ha5)))) : $signed(reg3874));
                    end
                  if ($signed((-{$signed(reg59)})))
                    begin
                      reg3933 <= ($signed(($signed((8'hb5)) <= $unsigned(reg3797))) >= ((reg3826[(1'h0):(1'h0)] & forvar3928) ?
                          reg3657 : $unsigned($unsigned(reg12))));
                      reg3934 <= (^~(((reg28 ?
                          reg3854 : reg3659) >>> (|reg61)) + ((reg3723 >= reg3918) | $signed(reg3815))));
                      reg3935 <= ({((~&reg3764) ?
                                  $signed(reg22) : (+reg3879))} ?
                          $signed(((reg3802 != reg3647) ?
                              (^~reg77) : (reg3694 * reg37))) : $unsigned((~|reg3656[(3'h4):(2'h3)])));
                      reg3936 <= reg3875[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg3933 <= $unsigned((8'hb1));
                    end
                  if ($signed(reg3869))
                    begin
                      reg3937 <= ((8'had) != $signed((reg3738[(1'h0):(1'h0)] && (8'hb7))));
                      reg3938 <= (((&(~|reg77)) ? reg3670 : (8'ha9)) ?
                          ($unsigned($unsigned(reg63)) || ((reg21 <= reg3858) >> (^reg3846))) : $unsigned({$signed(reg3718)}));
                      reg3939 <= {$unsigned({(~|(8'ha1))})};
                      reg3940 <= (reg3654[(3'h7):(1'h1)] ?
                          reg76[(1'h0):(1'h0)] : (|($signed(reg3731) <= $unsigned(reg3670))));
                    end
                  else
                    begin
                      reg3937 <= $unsigned(((reg3758[(1'h1):(1'h1)] > reg3825) & reg3832[(4'hb):(3'h7)]));
                      reg3938 <= reg3785;
                      reg3939 <= (($unsigned({reg3787}) == (+{reg3931})) - (reg3761[(3'h6):(3'h6)] ?
                          (!(~reg3882)) : $signed((reg76 ?
                              reg3701 : reg3755))));
                      reg3940 <= reg3864;
                    end
                  if ((reg3835[(1'h1):(1'h0)] ~^ (reg69 * ((reg3811 | reg3813) ~^ (~reg34)))))
                    begin
                      reg3941 <= (($unsigned($unsigned((8'haa))) << (^~$unsigned(wire8))) ?
                          $unsigned($unsigned($unsigned((8'ha8)))) : $signed({reg3822}));
                      reg3942 <= $unsigned(reg3742[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg3941 <= reg3835[(3'h4):(3'h4)];
                      reg3942 <= reg3872[(5'h10):(4'h9)];
                      reg3943 <= $signed($unsigned($unsigned((~^reg17))));
                    end
                end
              if (reg24)
                begin
                  if (reg3932[(3'h6):(2'h2)])
                    begin
                      reg3944 <= $signed({(^~((8'h9d) - reg40))});
                      reg3945 <= $unsigned(reg3828);
                      reg3946 <= $unsigned((^((reg53 ? reg3724 : reg3641) ?
                          {reg3880} : reg3902[(4'h9):(2'h2)])));
                    end
                  else
                    begin
                      reg3944 <= $unsigned($unsigned($unsigned(reg3660[(4'ha):(4'h8)])));
                    end
                end
              else
                begin
                  if ($unsigned(reg3937))
                    begin
                      reg3944 <= reg20[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg3944 <= reg3877[(3'h5):(1'h0)];
                      reg3945 <= $unsigned(($signed((reg3652 == reg3737)) ?
                          reg3895[(3'h6):(3'h4)] : ({reg3802} ?
                              (^reg3884) : $unsigned((8'hab)))));
                      reg3946 <= $unsigned($unsigned((forvar3921 >>> $signed(reg3894))));
                      reg3947 <= reg3799[(1'h1):(1'h0)];
                    end
                end
              reg3948 <= {$unsigned(reg3753[(3'h5):(3'h5)])};
            end
          if ($unsigned((($signed(reg3748) + (reg3924 & reg3675)) ?
              reg50 : (8'ha5))))
            begin
              for (forvar3949 = (1'h0); (forvar3949 < (1'h1)); forvar3949 = (forvar3949 + (1'h1)))
                begin
                  for (forvar3950 = (1'h0); (forvar3950 < (2'h3)); forvar3950 = (forvar3950 + (1'h1)))
                    begin
                      reg3951 <= $signed($signed(((reg77 ? reg3833 : (8'hb5)) ?
                          (reg3647 ? reg31 : reg25) : (reg3781 * reg3742))));
                      reg3952 <= (reg3715 > ($signed((reg3947 + wire8)) ?
                          (^~$signed(reg50)) : reg43));
                      reg3953 <= {(~|reg3777)};
                    end
                  for (forvar3954 = (1'h0); (forvar3954 < (1'h1)); forvar3954 = (forvar3954 + (1'h1)))
                    begin
                      reg3955 <= {$signed((~&{reg3826}))};
                    end
                  if ((reg45[(4'h8):(2'h3)] ?
                      reg3899 : $signed(reg3824[(1'h0):(1'h0)])))
                    begin
                      reg3956 <= $signed($signed(((|reg3894) ?
                          forvar3920[(2'h3):(2'h3)] : reg3859)));
                      reg3957 <= (reg25[(3'h5):(2'h2)] ?
                          $unsigned(((forvar3926 - reg3643) ^~ (reg3828 ?
                              reg17 : reg3906))) : ((~|$unsigned(reg3818)) ?
                              ($signed(reg3715) <<< (reg3701 < reg3737)) : ((reg3652 << reg3769) ?
                                  (reg77 ?
                                      reg12 : reg3824) : $unsigned(reg3834))));
                      reg3958 <= $signed((((reg3742 <<< reg3835) <= (|reg3752)) ?
                          (8'h9d) : reg3768[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg3956 <= $signed($unsigned(((forvar3920 ?
                              reg3847 : reg3940) ?
                          $unsigned(reg34) : (reg76 >= reg3727))));
                      reg3957 <= {reg73[(3'h4):(1'h0)]};
                    end
                  for (forvar3959 = (1'h0); (forvar3959 < (2'h3)); forvar3959 = (forvar3959 + (1'h1)))
                    begin
                      reg3960 <= $unsigned(reg54[(3'h7):(3'h5)]);
                      reg3961 <= $unsigned(($unsigned((~|(8'ha5))) ^ ($unsigned(reg3857) < reg3649)));
                      reg3962 <= {{(^reg3686[(1'h0):(1'h0)])}};
                    end
                end
              for (forvar3963 = (1'h0); (forvar3963 < (2'h3)); forvar3963 = (forvar3963 + (1'h1)))
                begin
                  if ($signed({((~|reg3795) && (reg15 ? reg3645 : (8'hac)))}))
                    begin
                      reg3964 <= ((8'hb1) ?
                          (~^{(reg3961 ~^ reg3716)}) : (~|reg49));
                      reg3965 <= $unsigned(($signed((reg3863 + (8'hb1))) > ($signed(reg3767) <= reg46[(1'h1):(1'h0)])));
                      reg3966 <= ((reg12 ^~ (^~$signed(reg3796))) || (8'hba));
                      reg3967 <= ($unsigned($unsigned(reg3685)) ^ ($signed(reg3677[(4'ha):(4'h8)]) < reg3639[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg3964 <= reg3809;
                    end
                  if ($signed($signed(($signed(reg3813) - reg3937))))
                    begin
                      reg3968 <= reg3822[(1'h0):(1'h0)];
                      reg3969 <= $unsigned(((((8'hb4) ?
                          reg3864 : (8'hac)) ^~ reg3730) && (8'ha4)));
                    end
                  else
                    begin
                      reg3968 <= $signed((~^(8'hb6)));
                      reg3969 <= reg3698;
                    end
                  if (reg3662)
                    begin
                      reg3970 <= $unsigned(reg48[(4'h8):(4'h8)]);
                      reg3971 <= $signed($unsigned(reg3817));
                      reg3972 <= $signed($signed((8'ha1)));
                    end
                  else
                    begin
                      reg3970 <= reg3830;
                      reg3971 <= reg3935;
                      reg3972 <= (-$unsigned($signed((|(8'had)))));
                    end
                end
              reg3973 <= (~^reg3697[(4'h8):(3'h4)]);
            end
          else
            begin
              reg3949 <= $unsigned((8'ha4));
              reg3950 <= $signed($unsigned(reg3661[(4'hb):(4'h9)]));
              if (reg3679)
                begin
                  for (forvar3951 = (1'h0); (forvar3951 < (2'h2)); forvar3951 = (forvar3951 + (1'h1)))
                    begin
                      reg3952 <= (((~|$signed(reg3909)) ?
                              (reg24[(4'hf):(2'h3)] ?
                                  {reg3834} : (reg3813 | reg3675)) : (((8'h9e) ?
                                      reg13 : reg3973) ?
                                  $signed((8'hab)) : $signed(reg3726))) ?
                          ($signed((8'ha6)) << reg3962) : {reg3884[(1'h1):(1'h1)]});
                    end
                  for (forvar3953 = (1'h0); (forvar3953 < (2'h3)); forvar3953 = (forvar3953 + (1'h1)))
                    begin
                      reg3954 <= {$signed(reg3743)};
                      reg3955 <= reg3912;
                      reg3956 <= $signed(({(reg3642 ? reg3854 : forvar3953)} ?
                          $signed((8'haa)) : $signed($unsigned(reg68))));
                    end
                  for (forvar3957 = (1'h0); (forvar3957 < (1'h0)); forvar3957 = (forvar3957 + (1'h1)))
                    begin
                      reg3958 <= $unsigned($signed($signed($signed(reg3949))));
                      reg3959 <= reg3839;
                      reg3960 <= ((&reg3706) & (((reg3699 ? reg3853 : (8'hb2)) ?
                          $unsigned(reg77) : reg3947) + (reg3863[(4'h9):(3'h5)] ?
                          reg3869 : (reg3840 >>> reg3699))));
                      reg3961 <= $signed($signed($signed((reg3702 | (8'ha9)))));
                    end
                end
              else
                begin
                  reg3951 <= reg3897;
                  if ($unsigned({reg3753[(2'h3):(2'h3)]}))
                    begin
                      reg3952 <= ($unsigned($unsigned($unsigned((8'hb6)))) & (8'hba));
                    end
                  else
                    begin
                      reg3952 <= reg3752[(1'h0):(1'h0)];
                      reg3953 <= ($signed(reg3710) | ((forvar3951[(2'h3):(2'h2)] ?
                          (reg3691 ~^ (8'ha5)) : (reg57 & reg15)) >>> $unsigned((~|reg3958))));
                      reg3954 <= (^~($unsigned($signed(reg70)) == (8'haa)));
                      reg3955 <= (|(((forvar3929 ? reg3718 : reg3791) ?
                          (reg3951 ?
                              reg3952 : reg3784) : reg3750[(3'h4):(2'h3)]) - ($signed(reg3684) || (reg3909 ?
                          reg3824 : reg3837))));
                    end
                  if (((~&$unsigned(reg3897)) + $signed(($unsigned(reg3684) ?
                      (reg3773 ? (8'ha0) : reg3946) : reg3790[(4'h8):(3'h7)]))))
                    begin
                      reg3956 <= $signed($unsigned((((8'hb7) > (8'ha2)) ?
                          (~^reg3691) : (-reg3683))));
                      reg3957 <= reg3734[(1'h1):(1'h1)];
                      reg3958 <= {(~$signed((reg45 == reg3859)))};
                    end
                  else
                    begin
                      reg3956 <= reg3949[(2'h2):(1'h0)];
                      reg3957 <= reg60;
                      reg3958 <= $unsigned({$signed({(8'hb3)})});
                      reg3959 <= $signed(reg48);
                    end
                  if ($signed((~|((reg3950 != forvar3922) ?
                      $signed(reg3841) : {(8'hb6)}))))
                    begin
                      reg3960 <= $unsigned(reg3745);
                    end
                  else
                    begin
                      reg3960 <= $unsigned(reg3849);
                      reg3961 <= $unsigned(($unsigned((&reg3809)) <= (((8'hb8) ^ reg3950) ?
                          (reg3750 + (8'hb0)) : $signed(reg3880))));
                    end
                end
              for (forvar3962 = (1'h0); (forvar3962 < (1'h0)); forvar3962 = (forvar3962 + (1'h1)))
                begin
                  for (forvar3963 = (1'h0); (forvar3963 < (2'h2)); forvar3963 = (forvar3963 + (1'h1)))
                    begin
                      reg3964 <= {(((wire3634 >> (8'hb9)) ?
                              {(8'hb8)} : $unsigned(reg3973)) - (~&(wire85 >> reg3942)))};
                      reg3965 <= (forvar3929[(1'h1):(1'h0)] ?
                          $signed((~{reg3939})) : $unsigned(((-reg3852) + (reg3805 ?
                              forvar3920 : reg3931))));
                    end
                end
            end
        end
      if ((8'hac))
        begin
          for (forvar3974 = (1'h0); (forvar3974 < (1'h0)); forvar3974 = (forvar3974 + (1'h1)))
            begin
              for (forvar3975 = (1'h0); (forvar3975 < (2'h3)); forvar3975 = (forvar3975 + (1'h1)))
                begin
                  if (wire5)
                    begin
                      reg3976 <= ({forvar3962} >> reg3911[(1'h1):(1'h1)]);
                      reg3977 <= $unsigned($signed($signed(reg3827[(1'h1):(1'h1)])));
                      reg3978 <= $unsigned((&(((8'hb6) ? (8'ha9) : wire3632) ?
                          reg3666[(4'he):(3'h5)] : reg3836)));
                    end
                  else
                    begin
                      reg3976 <= $unsigned((|(|$unsigned(reg3815))));
                      reg3977 <= (reg3841 ?
                          ((+reg3972[(3'h7):(3'h6)]) ?
                              $unsigned((reg3948 ?
                                  reg3681 : reg3972)) : reg51) : reg56);
                      reg3978 <= $unsigned(($signed((~reg12)) ?
                          $unsigned((&reg68)) : (^~(reg3719 ?
                              reg3960 : (8'ha7)))));
                    end
                  reg3979 <= $unsigned(forvar3920[(1'h0):(1'h0)]);
                  for (forvar3980 = (1'h0); (forvar3980 < (2'h3)); forvar3980 = (forvar3980 + (1'h1)))
                    begin
                      reg3981 <= (^($unsigned($signed(reg3971)) == (reg3729[(3'h4):(2'h3)] * (reg3696 ?
                          reg27 : reg3886))));
                      reg3982 <= reg3725;
                      reg3983 <= ($unsigned({$unsigned(reg3895)}) | (~|(~$signed(reg3716))));
                      reg3984 <= {$unsigned($unsigned((reg3652 ?
                              reg3810 : reg69)))};
                    end
                  if ($signed((reg3752 ?
                      $signed($unsigned(reg3859)) : $signed((reg19 ?
                          reg73 : reg3659)))))
                    begin
                      reg3985 <= {$unsigned($unsigned((~reg3746)))};
                      reg3986 <= ({reg3925} ^~ $signed(reg3854[(3'h6):(2'h3)]));
                      reg3987 <= reg3815;
                      reg3988 <= (8'hb5);
                    end
                  else
                    begin
                      reg3985 <= $unsigned($signed($unsigned($unsigned(reg10))));
                      reg3986 <= (!{((+reg3687) ^~ $unsigned(reg31))});
                      reg3987 <= $signed((reg81 ?
                          $unsigned(reg3973[(2'h2):(1'h1)]) : reg3847));
                      reg3988 <= reg3841[(4'hb):(1'h1)];
                    end
                end
              if (forvar3922[(2'h2):(1'h1)])
                begin
                  for (forvar3989 = (1'h0); (forvar3989 < (1'h1)); forvar3989 = (forvar3989 + (1'h1)))
                    begin
                      reg3990 <= (~&(^$signed(wire7)));
                      reg3991 <= (|(-$signed(reg3835)));
                      reg3992 <= (reg3864 ?
                          (($signed(reg3914) <= $unsigned(reg3879)) ?
                              reg3840[(4'h8):(3'h4)] : (((8'haa) - reg3933) ?
                                  $signed(reg81) : ((8'ha2) <<< reg3958))) : reg3672[(1'h0):(1'h0)]);
                      reg3993 <= (~{{(&reg18)}});
                    end
                  reg3994 <= reg3982;
                  if (reg3737)
                    begin
                      reg3995 <= (reg3992 ?
                          $unsigned(((reg3864 ?
                              reg3902 : (8'hab)) < reg40)) : ($unsigned(reg3661) ?
                              $unsigned($signed(reg3712)) : reg3643[(2'h3):(2'h3)]));
                      reg3996 <= $signed((reg3955 ?
                          (~|((8'hb2) ?
                              reg3695 : forvar3929)) : $signed((-reg3915))));
                    end
                  else
                    begin
                      reg3995 <= $unsigned(reg3902[(3'h5):(2'h3)]);
                      reg3996 <= {reg3696[(4'ha):(2'h2)]};
                    end
                end
              else
                begin
                  if (reg64)
                    begin
                      reg3989 <= reg3777;
                      reg3990 <= $unsigned(reg50[(3'h7):(3'h6)]);
                      reg3991 <= (reg3846 ?
                          reg68 : $unsigned(((reg3992 ?
                              (8'ha5) : reg3903) && {reg3787})));
                    end
                  else
                    begin
                      reg3989 <= reg3822;
                      reg3990 <= ((($signed(reg3954) && {reg3681}) | $signed(((8'ha1) ?
                              reg3700 : (8'hb8)))) ?
                          (^(reg3959 >>> $signed(reg3964))) : (~|reg80[(2'h3):(1'h0)]));
                    end
                end
            end
        end
      else
        begin
          reg3974 <= reg3991[(4'hc):(2'h3)];
          for (forvar3975 = (1'h0); (forvar3975 < (1'h1)); forvar3975 = (forvar3975 + (1'h1)))
            begin
              if ($unsigned($signed((+$unsigned((8'hae))))))
                begin
                  for (forvar3976 = (1'h0); (forvar3976 < (2'h3)); forvar3976 = (forvar3976 + (1'h1)))
                    begin
                      reg3977 <= $unsigned($unsigned(($signed(reg3943) * ((8'had) ?
                          (8'h9d) : wire3720))));
                      reg3978 <= ({(+$signed(reg3937))} >> (forvar3922[(3'h4):(1'h1)] >= reg3824));
                      reg3979 <= ((reg83[(4'hb):(1'h1)] ?
                          $unsigned((reg3647 ^~ reg32)) : $signed((!reg3936))) != $signed((reg3679 ~^ (reg3657 < reg79))));
                    end
                  for (forvar3980 = (1'h0); (forvar3980 < (1'h0)); forvar3980 = (forvar3980 + (1'h1)))
                    begin
                      reg3981 <= reg3845;
                    end
                end
              else
                begin
                  for (forvar3976 = (1'h0); (forvar3976 < (1'h1)); forvar3976 = (forvar3976 + (1'h1)))
                    begin
                      reg3977 <= $signed($unsigned((8'hb9)));
                      reg3978 <= $signed($signed($signed((!(8'hb2)))));
                      reg3979 <= (reg3790[(4'hf):(1'h0)] ?
                          (8'hab) : (({reg3729} ?
                                  (|reg3742) : (reg3978 * reg3931)) ?
                              ((reg3974 ?
                                  (8'hb8) : reg20) >> $unsigned(reg3786)) : $unsigned(reg31)));
                      reg3980 <= reg3951;
                    end
                  for (forvar3981 = (1'h0); (forvar3981 < (1'h0)); forvar3981 = (forvar3981 + (1'h1)))
                    begin
                      reg3982 <= reg3950[(2'h3):(1'h0)];
                      reg3983 <= (~((|reg3791) ?
                          ($unsigned(reg3943) ?
                              {reg3882} : {reg3849}) : reg3918[(1'h0):(1'h0)]));
                      reg3984 <= $unsigned((((forvar3962 ? reg3776 : (8'ha7)) ?
                              $unsigned(reg3698) : (!reg26)) ?
                          reg3685[(2'h2):(1'h1)] : (wire8[(2'h3):(2'h2)] ?
                              (reg3834 ? reg3925 : reg44) : (!reg3876))));
                      reg3985 <= reg3730[(1'h0):(1'h0)];
                    end
                end
              for (forvar3986 = (1'h0); (forvar3986 < (1'h0)); forvar3986 = (forvar3986 + (1'h1)))
                begin
                  for (forvar3987 = (1'h0); (forvar3987 < (2'h2)); forvar3987 = (forvar3987 + (1'h1)))
                    begin
                      reg3988 <= reg3969;
                      reg3989 <= $signed(reg3755[(4'hc):(4'hb)]);
                      reg3990 <= (reg3662 <<< wire6[(3'h6):(2'h2)]);
                    end
                  for (forvar3991 = (1'h0); (forvar3991 < (2'h3)); forvar3991 = (forvar3991 + (1'h1)))
                    begin
                      reg3992 <= reg3719;
                      reg3993 <= (((forvar3987[(4'ha):(2'h2)] + (reg44 ?
                              reg3693 : reg3731)) ?
                          (8'hb1) : (~^reg3860[(1'h1):(1'h1)])) && reg3871[(1'h0):(1'h0)]);
                    end
                  for (forvar3994 = (1'h0); (forvar3994 < (2'h3)); forvar3994 = (forvar3994 + (1'h1)))
                    begin
                      reg3995 <= reg3943;
                      reg3996 <= {wire3636};
                      reg3997 <= $signed($unsigned((&$unsigned(reg3826))));
                      reg3998 <= {(!((reg3798 && reg3872) ?
                              (-(8'had)) : $signed(reg3791)))};
                    end
                end
              if ((+reg3682))
                begin
                  for (forvar3999 = (1'h0); (forvar3999 < (2'h2)); forvar3999 = (forvar3999 + (1'h1)))
                    begin
                      reg4000 <= (!reg63[(1'h1):(1'h1)]);
                      reg4001 <= (-(reg3751[(4'hf):(4'hd)] != $unsigned($unsigned(forvar3987))));
                      reg4002 <= ((($signed(reg3784) ?
                          $unsigned(reg3971) : (reg3722 ~^ reg3958)) <= (^~(reg3996 ?
                          reg3758 : forvar3987))) || {(8'h9f)});
                    end
                  for (forvar4003 = (1'h0); (forvar4003 < (2'h3)); forvar4003 = (forvar4003 + (1'h1)))
                    begin
                      reg4004 <= $signed((((reg3766 ? reg14 : reg3756) ?
                          {reg3847} : {forvar3951}) <<< {(^reg3777)}));
                      reg4005 <= $unsigned($signed((reg3993 + reg25)));
                    end
                  if ($unsigned(reg3955))
                    begin
                      reg4006 <= (((reg46[(3'h5):(2'h3)] ?
                                  (~|reg3847) : $signed(reg3713)) ?
                              (reg3946[(1'h0):(1'h0)] ?
                                  $signed(reg3983) : (reg3869 ?
                                      reg73 : (8'hb8))) : reg3952[(3'h6):(3'h4)]) ?
                          ((forvar3922[(2'h2):(2'h2)] & $signed(reg3738)) == reg3970) : $signed((~|reg3804[(3'h7):(3'h4)])));
                      reg4007 <= forvar3949;
                    end
                  else
                    begin
                      reg4006 <= ((({(8'ha4)} >= (reg3864 ?
                                  reg4004 : reg3717)) ?
                              reg3679 : $signed((reg3709 ?
                                  reg3994 : reg3766))) ?
                          (+reg3943[(4'hc):(4'h8)]) : {((~&reg3697) ?
                                  (8'h9e) : $unsigned((8'ha2)))});
                      reg4007 <= $signed($unsigned(reg60));
                    end
                  if ($signed(({reg32[(3'h4):(1'h0)]} != $signed(forvar3975[(2'h3):(1'h1)]))))
                    begin
                      reg4008 <= $signed((((8'ha2) ?
                          forvar3999 : (reg3908 << reg3995)) <= ({reg4007} | $signed(reg3854))));
                    end
                  else
                    begin
                      reg4008 <= {$signed($unsigned((reg3916 ^ reg3697)))};
                      reg4009 <= (($signed($unsigned(reg3992)) ~^ (8'ha2)) <= (^~{{reg3841}}));
                      reg4010 <= ((-((^~reg40) | (reg3841 == reg4004))) | (!(~|forvar3950[(2'h3):(1'h0)])));
                      reg4011 <= forvar3954;
                    end
                end
              else
                begin
                  if ((~^$unsigned(reg84)))
                    begin
                      reg3999 <= $unsigned((((wire6 < reg3847) ?
                          $unsigned(reg3872) : reg63[(1'h0):(1'h0)]) >>> {$unsigned(forvar3999)}));
                      reg4000 <= reg3980[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg3999 <= $signed(((reg3932 <= wire3919) != (reg3667 - {reg4001})));
                      reg4000 <= (($unsigned(reg3994) ?
                          (&(reg3937 && (8'h9c))) : {(forvar3920 ?
                                  reg3726 : reg3662)}) ^ {((8'ha2) <<< $unsigned((8'hb8)))});
                      reg4001 <= $signed({$unsigned((^~reg31))});
                      reg4002 <= $unsigned((8'ha6));
                    end
                  for (forvar4003 = (1'h0); (forvar4003 < (2'h3)); forvar4003 = (forvar4003 + (1'h1)))
                    begin
                      reg4004 <= $signed((reg80[(1'h1):(1'h1)] ?
                          reg49[(2'h3):(2'h2)] : reg3815[(1'h1):(1'h0)]));
                      reg4005 <= (({(reg3805 == reg3841)} + $unsigned(((8'haf) ?
                              reg3991 : reg3939))) ?
                          (reg3728[(3'h4):(2'h3)] ?
                              (^(forvar3994 ?
                                  (8'ha2) : reg3794)) : reg3960) : reg31[(2'h3):(1'h0)]);
                      reg4006 <= $signed({((reg3764 > wire8) <<< reg3705[(3'h7):(2'h2)])});
                    end
                  if (($signed($signed((reg3816 ? forvar3962 : reg3999))) ?
                      $signed($unsigned($unsigned(reg3925))) : ({$unsigned(reg3790)} ?
                          (^reg4008) : forvar3999)))
                    begin
                      reg4007 <= reg3863[(3'h6):(3'h5)];
                      reg4008 <= ((-$unsigned((reg27 ?
                          reg52 : reg3675))) >>> $signed((~|reg61)));
                    end
                  else
                    begin
                      reg4007 <= ((((!reg24) || reg3748) | reg3994[(3'h6):(3'h6)]) ?
                          $signed($signed(reg46)) : reg3855);
                      reg4008 <= (reg3697 ?
                          (reg64[(2'h2):(2'h2)] ?
                              $signed({reg3931}) : ((reg3739 ?
                                  reg3811 : reg3966) << $unsigned(reg3895))) : {{(~&reg3895)}});
                    end
                  if ((^~$signed($signed($unsigned(reg3748)))))
                    begin
                      reg4009 <= $signed(reg3824);
                    end
                  else
                    begin
                      reg4009 <= $unsigned(($signed((~|(8'ha0))) ?
                          (+reg3714[(1'h1):(1'h0)]) : reg3753[(3'h5):(3'h5)]));
                      reg4010 <= (8'hb5);
                      reg4011 <= {($signed((reg3733 && (8'hba))) ?
                              reg53 : $signed(reg3691[(2'h3):(1'h1)]))};
                    end
                end
              if ((reg4011 && $signed(((reg3942 | reg3916) <<< reg3998[(2'h2):(1'h1)]))))
                begin
                  if (reg3755[(3'h5):(1'h1)])
                    begin
                      reg4012 <= reg3976[(3'h4):(1'h1)];
                      reg4013 <= {reg3804};
                      reg4014 <= (~$signed($signed((reg3694 ?
                          (8'hb5) : reg3674))));
                      reg4015 <= ({$signed((8'h9c))} || (reg3772 ?
                          ((reg63 > reg3902) < (reg77 ?
                              reg3805 : reg3907)) : (8'haa)));
                    end
                  else
                    begin
                      reg4012 <= ((~|($unsigned(forvar3953) ?
                              $signed(reg3706) : $signed(reg20))) ?
                          (&{reg44[(2'h2):(1'h1)]}) : $unsigned(reg3906[(2'h3):(1'h0)]));
                      reg4013 <= (reg16[(3'h4):(2'h2)] <<< $unsigned(reg3886));
                      reg4014 <= (8'hb6);
                      reg4015 <= ({$signed((8'ha8))} ?
                          $signed(((reg3867 ^~ reg3942) != $unsigned(reg76))) : {($unsigned(reg3830) || (!reg4014))});
                    end
                end
              else
                begin
                  for (forvar4012 = (1'h0); (forvar4012 < (2'h2)); forvar4012 = (forvar4012 + (1'h1)))
                    begin
                      reg4013 <= $signed({({reg15} ?
                              (reg3713 == reg3999) : reg3876[(1'h1):(1'h1)])});
                      reg4014 <= reg3936;
                      reg4015 <= $unsigned(reg3748[(3'h5):(2'h2)]);
                      reg4016 <= $signed($signed(reg17));
                    end
                  reg4017 <= $signed($signed(($unsigned(reg3938) >> (reg52 ?
                      reg60 : reg3677))));
                  for (forvar4018 = (1'h0); (forvar4018 < (2'h2)); forvar4018 = (forvar4018 + (1'h1)))
                    begin
                      reg4019 <= $unsigned(forvar3962);
                      reg4020 <= reg3698[(2'h2):(1'h0)];
                      reg4021 <= $unsigned(reg51[(4'h9):(1'h1)]);
                      reg4022 <= reg3651;
                    end
                end
            end
          for (forvar4023 = (1'h0); (forvar4023 < (1'h1)); forvar4023 = (forvar4023 + (1'h1)))
            begin
              for (forvar4024 = (1'h0); (forvar4024 < (1'h0)); forvar4024 = (forvar4024 + (1'h1)))
                begin
                  if ($signed((!{reg56})))
                    begin
                      reg4025 <= (!$unsigned($unsigned((8'hb9))));
                    end
                  else
                    begin
                      reg4025 <= (reg68 ?
                          ($unsigned(reg3723) > $signed(reg49)) : $unsigned(((forvar3926 || reg3690) ?
                              $signed(reg4010) : (reg3840 * reg31))));
                      reg4026 <= ({reg3855[(4'h8):(3'h7)]} ?
                          forvar3950[(2'h3):(1'h1)] : ($unsigned((&forvar3926)) ?
                              {(reg3836 == (8'hb5))} : ((reg3667 ^ reg3658) ?
                                  $signed((8'haf)) : (reg15 >> reg3850))));
                      reg4027 <= (^~$unsigned($unsigned((reg3719 ?
                          reg3864 : reg3865))));
                      reg4028 <= (reg3776 ?
                          reg3947[(4'h9):(3'h4)] : {$unsigned(reg3652)});
                    end
                  for (forvar4029 = (1'h0); (forvar4029 < (1'h1)); forvar4029 = (forvar4029 + (1'h1)))
                    begin
                      reg4030 <= reg3806;
                      reg4031 <= reg3651;
                      reg4032 <= (($signed(((8'h9f) && (8'hb4))) >>> (^~$unsigned(reg3723))) <= forvar3991);
                      reg4033 <= {$unsigned(reg3797)};
                    end
                  reg4034 <= $signed((reg15 ?
                      reg3703[(2'h3):(1'h1)] : reg4017[(1'h1):(1'h1)]));
                  for (forvar4035 = (1'h0); (forvar4035 < (1'h1)); forvar4035 = (forvar4035 + (1'h1)))
                    begin
                      reg4036 <= ($signed(((^reg3846) ?
                          wire3634 : reg3863[(3'h7):(1'h1)])) - reg4013);
                      reg4037 <= $signed((reg4001[(2'h2):(2'h2)] ?
                          {wire6} : {{reg3877}}));
                      reg4038 <= (!((~|{(8'hb1)}) < (!(~|reg3973))));
                    end
                end
            end
          reg4039 <= $signed(($signed($signed(reg3811)) ?
              $signed(reg60[(3'h4):(2'h3)]) : $unsigned({reg3945})));
        end
    end
  always
    @(posedge clk) begin
      if ({$unsigned($unsigned(reg54))})
        begin
          reg4040 <= reg4014;
        end
      else
        begin
          reg4040 <= ($signed($signed($signed((8'hb8)))) ?
              reg3644[(1'h0):(1'h0)] : $signed((reg3697[(2'h2):(2'h2)] ^ $signed(reg4027))));
          for (forvar4041 = (1'h0); (forvar4041 < (2'h2)); forvar4041 = (forvar4041 + (1'h1)))
            begin
              if (reg3877[(3'h6):(3'h6)])
                begin
                  reg4042 <= ((8'hb1) < (^reg3872[(2'h3):(1'h0)]));
                  reg4043 <= (^~reg3712);
                  for (forvar4044 = (1'h0); (forvar4044 < (2'h3)); forvar4044 = (forvar4044 + (1'h1)))
                    begin
                      reg4045 <= ((reg3970[(3'h6):(3'h4)] ?
                              $unsigned(reg3659[(3'h4):(3'h4)]) : reg3858[(3'h7):(1'h1)]) ?
                          (reg3857[(3'h5):(1'h1)] == reg10) : $signed({((8'hac) * reg3800)}));
                    end
                end
              else
                begin
                  for (forvar4042 = (1'h0); (forvar4042 < (1'h1)); forvar4042 = (forvar4042 + (1'h1)))
                    begin
                      reg4043 <= reg3997[(2'h2):(2'h2)];
                    end
                  for (forvar4044 = (1'h0); (forvar4044 < (1'h1)); forvar4044 = (forvar4044 + (1'h1)))
                    begin
                      reg4045 <= reg3797;
                      reg4046 <= $unsigned((&{$signed(reg3795)}));
                      reg4047 <= $unsigned((({reg3738} + $signed(reg4008)) ?
                          $signed(reg3949) : reg3994));
                    end
                end
              if ((&$unsigned((8'ha0))))
                begin
                  for (forvar4048 = (1'h0); (forvar4048 < (2'h2)); forvar4048 = (forvar4048 + (1'h1)))
                    begin
                      reg4049 <= (~&(|{((8'haa) >= reg3994)}));
                      reg4050 <= {(!$signed($signed(reg17)))};
                      reg4051 <= $signed(($unsigned(reg3934[(4'ha):(3'h7)]) | $unsigned((reg3836 ?
                          reg3815 : reg3767))));
                    end
                  if (reg4039)
                    begin
                      reg4052 <= $unsigned(reg3818[(3'h7):(2'h3)]);
                      reg4053 <= $unsigned(($unsigned((~reg28)) ?
                          reg18[(3'h5):(3'h4)] : (reg4012 <= $unsigned(reg3786))));
                      reg4054 <= (~reg72);
                      reg4055 <= {$signed(reg3834[(3'h7):(3'h7)])};
                    end
                  else
                    begin
                      reg4052 <= $unsigned((($unsigned(reg3688) ?
                              (forvar4044 ~^ reg4050) : (-reg3998)) ?
                          reg3818[(3'h5):(3'h4)] : $signed((~&(8'hba)))));
                      reg4053 <= reg3850;
                    end
                  reg4056 <= (({(wire6 ^ reg25)} ?
                      (reg71[(4'hc):(4'h8)] >>> (~reg3877)) : {(~&reg3953)}) & reg3723);
                  if ((|((~^$unsigned(reg4001)) ?
                      reg3658 : ($unsigned((8'hb2)) ?
                          $unsigned(reg3769) : reg28))))
                    begin
                      reg4057 <= reg3875;
                      reg4058 <= ({reg3718} != ((-(reg3988 ?
                              reg3737 : reg3666)) ?
                          ($signed(reg4004) + (reg3844 ?
                              wire85 : reg3956)) : (((8'haf) >> reg3952) ?
                              (~reg18) : $signed(reg3842))));
                    end
                  else
                    begin
                      reg4057 <= $signed(reg47[(1'h0):(1'h0)]);
                      reg4058 <= (reg4005 || $unsigned(((reg3653 <<< reg3764) ?
                          $signed(reg3971) : $unsigned(reg4058))));
                      reg4059 <= reg3827[(4'hb):(4'ha)];
                    end
                end
              else
                begin
                  for (forvar4048 = (1'h0); (forvar4048 < (1'h0)); forvar4048 = (forvar4048 + (1'h1)))
                    begin
                      reg4049 <= $signed((reg3751[(4'hd):(1'h1)] == ($signed(reg3895) + (reg3868 || reg3653))));
                      reg4050 <= (&$unsigned(reg3933[(2'h2):(1'h1)]));
                      reg4051 <= $signed(reg3755);
                    end
                  if ($signed((reg3977 >> reg3956[(4'h8):(1'h1)])))
                    begin
                      reg4052 <= reg3766;
                      reg4053 <= {reg3992};
                    end
                  else
                    begin
                      reg4052 <= $signed((reg3980[(2'h3):(1'h1)] ?
                          reg3946[(1'h1):(1'h1)] : (+(wire3636 | reg3769))));
                      reg4053 <= reg3742;
                      reg4054 <= reg3666;
                    end
                  for (forvar4055 = (1'h0); (forvar4055 < (2'h2)); forvar4055 = (forvar4055 + (1'h1)))
                    begin
                      reg4056 <= {($signed((|reg3804)) ?
                              ((reg3995 && reg3757) - {reg3726}) : reg3681)};
                      reg4057 <= reg3681[(1'h0):(1'h0)];
                      reg4058 <= ($unsigned((!$signed(reg3902))) ~^ $signed((~reg3993)));
                      reg4059 <= reg3704[(4'hb):(3'h4)];
                    end
                end
            end
          for (forvar4060 = (1'h0); (forvar4060 < (2'h3)); forvar4060 = (forvar4060 + (1'h1)))
            begin
              for (forvar4061 = (1'h0); (forvar4061 < (1'h1)); forvar4061 = (forvar4061 + (1'h1)))
                begin
                  for (forvar4062 = (1'h0); (forvar4062 < (1'h0)); forvar4062 = (forvar4062 + (1'h1)))
                    begin
                      reg4063 <= ({$unsigned((^~reg3937))} >>> reg3944[(1'h0):(1'h0)]);
                      reg4064 <= $signed(({reg3879} * $signed($unsigned(reg3982))));
                    end
                end
              reg4065 <= ({(!(reg3848 * (8'ha8)))} | (+($signed((8'haa)) + $unsigned(reg3906))));
              if (reg3906[(2'h3):(2'h2)])
                begin
                  for (forvar4066 = (1'h0); (forvar4066 < (2'h3)); forvar4066 = (forvar4066 + (1'h1)))
                    begin
                      reg4067 <= $unsigned($unsigned(reg3736));
                    end
                end
              else
                begin
                  for (forvar4066 = (1'h0); (forvar4066 < (2'h3)); forvar4066 = (forvar4066 + (1'h1)))
                    begin
                      reg4067 <= (^{$unsigned((8'ha0))});
                    end
                  reg4068 <= {reg3728};
                end
              if ((reg16 ?
                  ((&(reg3988 & reg3809)) == ($signed(reg3835) ?
                      (reg3882 == reg3840) : {reg3681})) : $unsigned(reg4040)))
                begin
                  for (forvar4069 = (1'h0); (forvar4069 < (2'h2)); forvar4069 = (forvar4069 + (1'h1)))
                    begin
                      reg4070 <= reg4021[(4'h9):(3'h7)];
                      reg4071 <= $signed((reg20 > {reg3699}));
                      reg4072 <= reg3733[(3'h6):(3'h4)];
                    end
                end
              else
                begin
                  if ($unsigned(((~reg3974) ^~ reg4030[(2'h2):(2'h2)])))
                    begin
                      reg4069 <= (-(^~reg3725));
                      reg4070 <= $unsigned($signed((~&reg4050[(4'h9):(2'h3)])));
                      reg4071 <= reg3647[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg4069 <= (8'hb2);
                      reg4070 <= (8'hac);
                      reg4071 <= reg3713[(3'h6):(2'h3)];
                      reg4072 <= reg3692;
                    end
                end
            end
          for (forvar4073 = (1'h0); (forvar4073 < (2'h2)); forvar4073 = (forvar4073 + (1'h1)))
            begin
              if (({reg3696[(1'h0):(1'h0)]} ?
                  (|$unsigned((reg3687 ? reg81 : reg3709))) : reg4045))
                begin
                  reg4074 <= reg3656;
                  if ((^~(!reg80)))
                    begin
                      reg4075 <= (reg3786 || reg4000);
                      reg4076 <= (reg3946[(3'h5):(2'h3)] + reg3991[(4'he):(3'h7)]);
                    end
                  else
                    begin
                      reg4075 <= (~^((~^$signed(reg13)) <= reg3934[(1'h1):(1'h1)]));
                    end
                end
              else
                begin
                  if (reg4057)
                    begin
                      reg4074 <= $unsigned((8'hab));
                    end
                  else
                    begin
                      reg4074 <= $signed($signed({(reg3798 ?
                              reg3844 : reg3786)}));
                      reg4075 <= ($unsigned($signed({reg3935})) <= (&$unsigned({reg3936})));
                      reg4076 <= reg4036[(4'hd):(4'h8)];
                    end
                  if (reg3951[(1'h1):(1'h1)])
                    begin
                      reg4077 <= reg3834[(3'h4):(1'h1)];
                      reg4078 <= wire8;
                      reg4079 <= (reg31 ? reg3687 : (~^reg3640[(2'h2):(1'h0)]));
                      reg4080 <= (($signed($signed(wire3720)) ?
                          (~|(!reg3817)) : reg4045[(1'h1):(1'h1)]) >= ($signed((reg3899 ^~ reg4045)) ?
                          (-(reg3839 ? (8'ha7) : reg3757)) : (reg3878 ?
                              (reg3698 ? (8'ha7) : reg3874) : (reg3815 ?
                                  reg3796 : forvar4041))));
                    end
                  else
                    begin
                      reg4077 <= {reg3692};
                      reg4078 <= reg4045[(4'h9):(4'h8)];
                      reg4079 <= (reg3913 ~^ {$signed(reg3914[(3'h4):(1'h0)])});
                      reg4080 <= reg3669;
                    end
                end
              for (forvar4081 = (1'h0); (forvar4081 < (2'h2)); forvar4081 = (forvar4081 + (1'h1)))
                begin
                  if ({{reg3829[(4'h8):(3'h4)]}})
                    begin
                      reg4082 <= $unsigned($signed($unsigned((reg3850 || reg3658))));
                      reg4083 <= ($signed((~^$unsigned(reg3705))) ?
                          reg3943 : ((|$signed((8'ha1))) ?
                              reg3755 : $unsigned((reg3865 && reg36))));
                      reg4084 <= ($signed(((^reg3871) != $signed(reg3716))) <<< {((reg4031 > reg70) ?
                              ((8'ha0) ? reg3923 : reg3775) : {reg3915})});
                    end
                  else
                    begin
                      reg4082 <= $unsigned({$unsigned({reg36})});
                    end
                  for (forvar4085 = (1'h0); (forvar4085 < (2'h3)); forvar4085 = (forvar4085 + (1'h1)))
                    begin
                      reg4086 <= $signed((~|$unsigned((-reg3871))));
                      reg4087 <= ((($unsigned(reg3738) ^ reg3661[(4'h9):(3'h4)]) ?
                          ($unsigned(wire5) & reg3665[(4'hb):(4'ha)]) : reg3689[(1'h1):(1'h1)]) ~^ reg3835[(2'h3):(2'h3)]);
                    end
                  reg4088 <= (reg3950 || (reg3739[(4'h9):(1'h0)] ?
                      wire3632[(1'h0):(1'h0)] : (~^$signed((8'haa)))));
                end
              reg4089 <= (((+{reg3784}) >= {$signed(reg3683)}) ?
                  ($signed((reg3717 ? (8'ha5) : reg4088)) ?
                      ((reg72 ? reg3988 : reg3673) ?
                          $unsigned(reg3806) : (reg74 & (8'hb4))) : $signed((8'hb3))) : ($unsigned($unsigned(reg3882)) > (reg3824 ?
                      (forvar4069 ? reg4014 : reg3909) : (reg3960 || reg45))));
              for (forvar4090 = (1'h0); (forvar4090 < (2'h2)); forvar4090 = (forvar4090 + (1'h1)))
                begin
                  for (forvar4091 = (1'h0); (forvar4091 < (1'h0)); forvar4091 = (forvar4091 + (1'h1)))
                    begin
                      reg4092 <= reg3757;
                      reg4093 <= $signed($signed($signed((~reg3899))));
                      reg4094 <= $unsigned(((8'h9c) ?
                          ($unsigned(reg3684) ?
                              {reg53} : (reg4017 + reg3863)) : ($unsigned(reg3786) ?
                              reg3931 : $signed(reg3996))));
                      reg4095 <= (($signed($signed(reg3668)) ?
                              (-(reg3738 >= reg3797)) : {(!reg3939)}) ?
                          $signed((~|(~|reg84))) : ($signed(reg3650) <= $unsigned($unsigned(forvar4073))));
                    end
                end
            end
        end
    end
  assign wire4096 = reg3767;
  assign wire4097 = {reg4038[(4'hb):(2'h3)]};
  assign wire4098 = reg3795[(4'h9):(2'h2)];
  assign wire4099 = {(reg4017 > (!(reg3643 != reg3966)))};
  assign wire4100 = reg3739;
  always
    @(posedge clk) begin
      if ($signed($signed((8'hb6))))
        begin
          if ((^(-reg3852)))
            begin
              if ({$unsigned((~|$signed(reg3670)))})
                begin
                  reg4101 <= ({$unsigned(reg51)} || (8'hb5));
                end
              else
                begin
                  reg4101 <= (~&(&(&(reg3815 ? reg3959 : reg3953))));
                end
            end
          else
            begin
              if (reg3805[(4'h8):(2'h2)])
                begin
                  for (forvar4101 = (1'h0); (forvar4101 < (1'h0)); forvar4101 = (forvar4101 + (1'h1)))
                    begin
                      reg4102 <= reg4038[(3'h7):(2'h3)];
                    end
                  for (forvar4103 = (1'h0); (forvar4103 < (1'h1)); forvar4103 = (forvar4103 + (1'h1)))
                    begin
                      reg4104 <= {$signed($unsigned($signed(reg56)))};
                      reg4105 <= (8'hba);
                      reg4106 <= $signed({reg3689[(2'h2):(1'h1)]});
                      reg4107 <= ($signed(reg3850) ?
                          ((^~{reg3643}) ?
                              ($signed(reg4078) ^ $signed(reg3905)) : (~(reg21 + reg3674))) : ({$signed((8'ha2))} & ((reg3641 ?
                              reg3690 : reg3734) | reg74)));
                    end
                  for (forvar4108 = (1'h0); (forvar4108 < (2'h2)); forvar4108 = (forvar4108 + (1'h1)))
                    begin
                      reg4109 <= $signed(((~^((8'hb3) >>> reg4088)) ?
                          reg3985 : (((8'h9e) ? reg4080 : (8'ha3)) ?
                              reg3659 : (reg59 || reg3984))));
                    end
                  if ((8'ha3))
                    begin
                      reg4110 <= reg44;
                      reg4111 <= $unsigned(reg4110[(1'h0):(1'h0)]);
                      reg4112 <= $signed((8'hae));
                      reg4113 <= (!(!(8'hba)));
                    end
                  else
                    begin
                      reg4110 <= ((reg43[(3'h5):(1'h1)] >>> (8'hac)) | reg73[(3'h4):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar4101 = (1'h0); (forvar4101 < (1'h0)); forvar4101 = (forvar4101 + (1'h1)))
                    begin
                      reg4102 <= reg4016;
                      reg4103 <= reg3784[(3'h7):(3'h4)];
                      reg4104 <= (8'ha2);
                    end
                  for (forvar4105 = (1'h0); (forvar4105 < (2'h3)); forvar4105 = (forvar4105 + (1'h1)))
                    begin
                      reg4106 <= ((reg3898 <= (reg3653[(4'ha):(4'h9)] ?
                              {reg3734} : reg3986[(1'h0):(1'h0)])) ?
                          $signed(reg3974[(1'h0):(1'h0)]) : (+$signed(reg3823)));
                      reg4107 <= $unsigned($signed(((reg3897 ?
                              reg3724 : reg3639) ?
                          (reg4046 << (8'h9d)) : (reg3790 >= reg3654))));
                      reg4108 <= ($signed($unsigned(((8'hb5) ?
                              (8'ha2) : reg19))) ?
                          $signed({(reg74 ? reg3933 : wire4097)}) : (reg3984 ?
                              $unsigned({(8'hb7)}) : reg3951));
                      reg4109 <= reg3898;
                    end
                end
              reg4114 <= reg3659[(3'h7):(2'h2)];
            end
        end
      else
        begin
          reg4101 <= (reg57[(1'h1):(1'h1)] ?
              $signed($unsigned(reg3764[(1'h0):(1'h0)])) : $unsigned($unsigned(reg3908[(3'h5):(1'h1)])));
          for (forvar4102 = (1'h0); (forvar4102 < (2'h3)); forvar4102 = (forvar4102 + (1'h1)))
            begin
              for (forvar4103 = (1'h0); (forvar4103 < (1'h0)); forvar4103 = (forvar4103 + (1'h1)))
                begin
                  for (forvar4104 = (1'h0); (forvar4104 < (1'h1)); forvar4104 = (forvar4104 + (1'h1)))
                    begin
                      reg4105 <= reg3771[(3'h7):(3'h7)];
                      reg4106 <= $unsigned($signed(reg3839[(2'h3):(2'h2)]));
                    end
                  for (forvar4107 = (1'h0); (forvar4107 < (1'h1)); forvar4107 = (forvar4107 + (1'h1)))
                    begin
                      reg4108 <= reg81;
                      reg4109 <= ({($unsigned(reg4092) || (reg3697 ?
                                  reg3983 : reg3646))} ?
                          reg3716[(2'h2):(1'h0)] : $unsigned($signed(reg3665[(3'h5):(2'h3)])));
                    end
                  reg4110 <= reg4014;
                end
              for (forvar4111 = (1'h0); (forvar4111 < (2'h3)); forvar4111 = (forvar4111 + (1'h1)))
                begin
                  reg4112 <= (reg3696 <<< ($signed((reg3795 ?
                          reg3743 : reg3927)) ?
                      (8'ha3) : reg3848));
                  for (forvar4113 = (1'h0); (forvar4113 < (1'h0)); forvar4113 = (forvar4113 + (1'h1)))
                    begin
                      reg4114 <= ($signed(((reg3873 | wire4098) <<< (+reg3705))) ?
                          $unsigned($unsigned((reg3955 - reg3806))) : (|{reg14}));
                    end
                  for (forvar4115 = (1'h0); (forvar4115 < (2'h2)); forvar4115 = (forvar4115 + (1'h1)))
                    begin
                      reg4116 <= (reg4008 ?
                          (($signed(reg3758) - reg3722[(3'h4):(3'h4)]) ?
                              reg3818[(1'h0):(1'h0)] : (forvar4101[(2'h2):(1'h1)] == reg3978)) : (8'hb3));
                      reg4117 <= reg75;
                      reg4118 <= reg3996[(4'ha):(3'h6)];
                    end
                end
              for (forvar4119 = (1'h0); (forvar4119 < (2'h2)); forvar4119 = (forvar4119 + (1'h1)))
                begin
                  for (forvar4120 = (1'h0); (forvar4120 < (2'h2)); forvar4120 = (forvar4120 + (1'h1)))
                    begin
                      reg4121 <= $signed({reg3670[(4'h8):(3'h5)]});
                      reg4122 <= (reg3935[(3'h4):(1'h0)] ?
                          $signed(reg3948) : (reg3641 ?
                              (~&reg3656[(3'h5):(3'h5)]) : $signed($signed((8'ha6)))));
                    end
                end
            end
          for (forvar4123 = (1'h0); (forvar4123 < (2'h2)); forvar4123 = (forvar4123 + (1'h1)))
            begin
              if ({reg3967[(3'h5):(3'h4)]})
                begin
                  if ((~^{(+$signed(reg47))}))
                    begin
                      reg4124 <= reg4009[(1'h1):(1'h1)];
                      reg4125 <= {$unsigned($signed(reg3837))};
                    end
                  else
                    begin
                      reg4124 <= (-($unsigned((^reg3739)) ?
                          ($signed(reg3933) & reg3849[(1'h1):(1'h0)]) : reg3942[(4'hb):(1'h1)]));
                    end
                  for (forvar4126 = (1'h0); (forvar4126 < (2'h2)); forvar4126 = (forvar4126 + (1'h1)))
                    begin
                      reg4127 <= $signed(reg3982);
                      reg4128 <= $unsigned({reg3771});
                    end
                end
              else
                begin
                  if ((^reg3911))
                    begin
                      reg4124 <= reg4072;
                      reg4125 <= $unsigned((($unsigned(reg3682) ~^ $signed(reg3927)) >>> reg4038[(1'h1):(1'h1)]));
                      reg4126 <= reg3959[(3'h6):(1'h1)];
                      reg4127 <= $signed($unsigned((~&reg4056)));
                    end
                  else
                    begin
                      reg4124 <= reg3730[(4'ha):(3'h6)];
                      reg4125 <= reg3968[(4'h9):(4'h8)];
                    end
                  if ($unsigned(reg3704))
                    begin
                      reg4128 <= reg4111[(3'h7):(3'h6)];
                      reg4129 <= reg4006;
                      reg4130 <= $signed($unsigned((&{reg3845})));
                    end
                  else
                    begin
                      reg4128 <= reg4079[(3'h6):(3'h5)];
                    end
                end
              for (forvar4131 = (1'h0); (forvar4131 < (2'h3)); forvar4131 = (forvar4131 + (1'h1)))
                begin
                  for (forvar4132 = (1'h0); (forvar4132 < (1'h0)); forvar4132 = (forvar4132 + (1'h1)))
                    begin
                      reg4133 <= reg3843[(1'h0):(1'h0)];
                      reg4134 <= ($unsigned($unsigned((!reg3777))) ?
                          $unsigned($unsigned((reg50 && reg16))) : wire4100[(2'h3):(1'h0)]);
                      reg4135 <= reg79[(2'h2):(1'h1)];
                      reg4136 <= $signed($signed(forvar4103[(2'h2):(1'h1)]));
                    end
                  if ((~&reg3943[(4'h8):(2'h3)]))
                    begin
                      reg4137 <= reg4093[(3'h6):(3'h4)];
                    end
                  else
                    begin
                      reg4137 <= reg3960[(4'hb):(3'h4)];
                    end
                  for (forvar4138 = (1'h0); (forvar4138 < (1'h1)); forvar4138 = (forvar4138 + (1'h1)))
                    begin
                      reg4139 <= ($signed(reg3785[(1'h1):(1'h0)]) ?
                          forvar4111 : ($signed(reg3815[(2'h2):(1'h0)]) >= (reg3864[(1'h1):(1'h0)] ?
                              (~^reg3964) : (reg4054 ? (8'ha2) : reg4124))));
                      reg4140 <= reg3785;
                      reg4141 <= ({(&reg3834[(2'h2):(1'h1)])} >>> (reg3729 <<< reg3773[(1'h1):(1'h1)]));
                      reg4142 <= ((reg3748 * ({reg3659} >>> reg4007)) ?
                          wire6[(2'h2):(2'h2)] : reg4013);
                    end
                end
              for (forvar4143 = (1'h0); (forvar4143 < (1'h0)); forvar4143 = (forvar4143 + (1'h1)))
                begin
                  for (forvar4144 = (1'h0); (forvar4144 < (1'h0)); forvar4144 = (forvar4144 + (1'h1)))
                    begin
                      reg4145 <= ((|$signed((8'ha9))) ?
                          ((|$unsigned(reg3849)) ?
                              $signed((reg3724 ?
                                  reg3871 : reg3794)) : $unsigned((reg3909 ?
                                  wire6 : reg3948))) : $unsigned({$unsigned(reg4039)}));
                    end
                  reg4146 <= reg3869;
                  for (forvar4147 = (1'h0); (forvar4147 < (2'h3)); forvar4147 = (forvar4147 + (1'h1)))
                    begin
                      reg4148 <= ((+(reg50 ? reg33 : (~reg3729))) ?
                          (~|reg3730[(3'h5):(3'h4)]) : ((~reg3665[(3'h7):(2'h2)]) + reg3982[(2'h3):(2'h2)]));
                    end
                  for (forvar4149 = (1'h0); (forvar4149 < (2'h3)); forvar4149 = (forvar4149 + (1'h1)))
                    begin
                      reg4150 <= ((8'hb6) ?
                          reg4067 : {$unsigned($unsigned(reg3877))});
                      reg4151 <= ({(!reg4002)} << {((reg3649 - reg3993) ?
                              {reg43} : reg76)});
                      reg4152 <= {$unsigned({(|(8'h9d))})};
                    end
                end
              reg4153 <= reg4032[(4'hb):(1'h1)];
            end
          for (forvar4154 = (1'h0); (forvar4154 < (1'h1)); forvar4154 = (forvar4154 + (1'h1)))
            begin
              for (forvar4155 = (1'h0); (forvar4155 < (1'h1)); forvar4155 = (forvar4155 + (1'h1)))
                begin
                  reg4156 <= ({((reg3749 ?
                          reg4021 : (8'hab)) ^ $signed(reg3935))} == $signed($unsigned((reg63 ?
                      reg3714 : (8'ha9)))));
                end
              reg4157 <= $signed((reg26[(3'h5):(3'h5)] ?
                  $unsigned((reg3763 > reg4036)) : $signed((|(8'ha5)))));
              reg4158 <= reg4114[(2'h2):(1'h1)];
              if ((-$unsigned((^~reg4025))))
                begin
                  reg4159 <= {$unsigned({((8'ha8) > reg3688)})};
                  for (forvar4160 = (1'h0); (forvar4160 < (2'h2)); forvar4160 = (forvar4160 + (1'h1)))
                    begin
                      reg4161 <= $unsigned($unsigned(reg3933));
                      reg4162 <= {(8'h9d)};
                      reg4163 <= reg3908[(2'h3):(1'h1)];
                    end
                  if (((((reg3902 > reg3927) < reg3709[(1'h0):(1'h0)]) ?
                      ((~^forvar4119) < reg4017) : $signed($unsigned((8'h9c)))) ^~ (|(!reg3980))))
                    begin
                      reg4164 <= reg3794;
                    end
                  else
                    begin
                      reg4164 <= reg3737;
                      reg4165 <= ({$unsigned({reg4014})} ?
                          (~|{$unsigned(reg3769)}) : reg3886[(1'h0):(1'h0)]);
                      reg4166 <= $signed((((~&reg4108) ?
                              (reg4010 && (8'ha0)) : reg3784[(4'hd):(3'h5)]) ?
                          $signed(reg4083) : $signed($unsigned(reg3827))));
                      reg4167 <= reg4101[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  if (({((~|reg3826) <= $signed((8'hb4)))} >= reg3811))
                    begin
                      reg4159 <= reg3786;
                    end
                  else
                    begin
                      reg4159 <= (forvar4149[(1'h1):(1'h1)] ?
                          (-{reg3988[(1'h1):(1'h0)]}) : (({reg83} | (reg4040 <<< reg3814)) ?
                              forvar4111[(3'h7):(1'h0)] : reg3976[(3'h7):(3'h6)]));
                      reg4160 <= $unsigned(reg4117);
                      reg4161 <= (reg4106 << $signed($unsigned($signed(reg3646))));
                      reg4162 <= ((~&$unsigned($signed(reg3981))) && $unsigned(reg57));
                    end
                  for (forvar4163 = (1'h0); (forvar4163 < (1'h1)); forvar4163 = (forvar4163 + (1'h1)))
                    begin
                      reg4164 <= ((8'hb3) ?
                          {{forvar4149[(2'h2):(2'h2)]}} : {$unsigned((reg4116 ?
                                  reg4057 : (8'ha7)))});
                      reg4165 <= reg4116;
                      reg4166 <= reg4118[(2'h2):(1'h1)];
                      reg4167 <= reg4117[(2'h3):(1'h0)];
                    end
                  for (forvar4168 = (1'h0); (forvar4168 < (1'h1)); forvar4168 = (forvar4168 + (1'h1)))
                    begin
                      reg4169 <= (~|(reg3932[(4'h8):(1'h0)] ?
                          ({reg4015} ?
                              $unsigned(wire8) : reg59) : reg3728[(1'h1):(1'h1)]));
                      reg4170 <= (8'hb4);
                      reg4171 <= (reg3739 ^~ $unsigned(($signed(reg4129) ?
                          reg4113[(1'h1):(1'h0)] : (reg3981 ? reg33 : reg69))));
                    end
                  if ($signed({$signed(reg3811[(2'h3):(1'h1)])}))
                    begin
                      reg4172 <= $unsigned(reg3706);
                      reg4173 <= ($unsigned({(reg3699 ? reg4063 : reg3796)}) ?
                          $signed(({reg4127} == $unsigned(reg3945))) : ($unsigned((reg3685 << wire8)) * $unsigned($signed(reg3656))));
                      reg4174 <= (reg3673 ?
                          (|reg4158[(2'h2):(1'h0)]) : $unsigned((~^reg4126)));
                      reg4175 <= (reg3952[(3'h4):(1'h0)] ^ reg4001[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg4172 <= $unsigned(((8'ha1) ?
                          (~&(~|(8'hb9))) : (((8'ha1) || reg3684) * (reg4173 ?
                              reg3642 : reg50))));
                      reg4173 <= (($signed(reg3915) || reg4031[(1'h1):(1'h0)]) * $signed($unsigned((reg3807 ~^ reg3987))));
                    end
                end
            end
        end
      for (forvar4176 = (1'h0); (forvar4176 < (1'h0)); forvar4176 = (forvar4176 + (1'h1)))
        begin
          for (forvar4177 = (1'h0); (forvar4177 < (1'h1)); forvar4177 = (forvar4177 + (1'h1)))
            begin
              if ($signed($signed($signed($unsigned(reg3706)))))
                begin
                  for (forvar4178 = (1'h0); (forvar4178 < (1'h1)); forvar4178 = (forvar4178 + (1'h1)))
                    begin
                      reg4179 <= reg3979;
                      reg4180 <= (reg3849 ^~ (((reg3644 > wire4098) ?
                          reg3802 : {(8'h9d)}) && $signed(reg4163)));
                      reg4181 <= $signed((($signed(reg4012) | forvar4154[(5'h10):(4'h9)]) << (8'ha9)));
                      reg4182 <= {$unsigned((reg3909 ? reg3794 : (|(8'ha9))))};
                    end
                  reg4183 <= $signed(((~|reg4153) ?
                      (reg3767 > (reg3832 ? reg3729 : reg3757)) : (reg3785 ?
                          (reg3942 ? (8'ha9) : reg4034) : (reg3939 ?
                              reg3880 : forvar4143))));
                  reg4184 <= $signed({reg4110[(1'h1):(1'h0)]});
                  if ({$signed((~&$signed(reg67)))})
                    begin
                      reg4185 <= (($unsigned((reg3916 ~^ reg3925)) ?
                          reg84 : reg3667[(2'h3):(1'h0)]) & (($unsigned(reg4174) ~^ (reg3882 >>> reg4125)) ?
                          reg4077 : reg3696[(3'h7):(3'h7)]));
                    end
                  else
                    begin
                      reg4185 <= $unsigned(($unsigned(reg3966[(3'h5):(2'h2)]) ?
                          (!{reg4009}) : $unsigned($unsigned(reg3879))));
                      reg4186 <= (8'hb4);
                      reg4187 <= ($signed($unsigned(reg3810[(2'h2):(1'h1)])) + $unsigned(reg3876));
                    end
                end
              else
                begin
                  reg4178 <= ($unsigned($signed(reg3734)) >= reg3886[(4'h8):(1'h0)]);
                  for (forvar4179 = (1'h0); (forvar4179 < (1'h1)); forvar4179 = (forvar4179 + (1'h1)))
                    begin
                      reg4180 <= ($signed((-reg3884)) ~^ $unsigned($unsigned($signed(reg3735))));
                      reg4181 <= (~(reg4101 ?
                          reg3706 : reg3852[(2'h2):(1'h1)]));
                      reg4182 <= ({$signed($signed(reg3692))} * reg4074);
                      reg4183 <= (reg4162 ?
                          (-{$unsigned(reg3949)}) : reg4021[(3'h5):(2'h2)]);
                    end
                  if ({$signed({((8'ha8) == reg4158)})})
                    begin
                      reg4184 <= ({((forvar4160 >>> reg4118) != $signed((8'h9f)))} > $unsigned($signed(reg3858[(3'h5):(2'h3)])));
                      reg4185 <= forvar4176[(1'h1):(1'h1)];
                      reg4186 <= ({(reg3964 >= reg4117)} ?
                          ({reg4071[(2'h3):(2'h3)]} ^~ ((reg3739 ~^ reg3990) + (~^reg4092))) : forvar4179);
                      reg4187 <= ((((reg3805 + (8'hb3)) ?
                          reg3882 : reg4057) ~^ reg79) ^ (|((reg3824 - (8'haf)) ~^ (reg3779 > reg3646))));
                    end
                  else
                    begin
                      reg4184 <= reg3804[(4'hb):(2'h3)];
                      reg4185 <= wire4096[(2'h2):(2'h2)];
                      reg4186 <= {$unsigned(reg4001)};
                      reg4187 <= (((^(~&reg3709)) << $signed(reg15)) ?
                          ((reg3991[(2'h2):(1'h0)] > $signed(reg26)) ?
                              ((reg3768 >>> reg3978) ?
                                  reg67 : {reg3886}) : $signed((reg3697 || reg3660))) : $signed(((!reg4152) ?
                              (forvar4163 < reg3983) : $unsigned(reg3827))));
                    end
                end
            end
          if ($signed(reg52))
            begin
              if (reg3964[(3'h5):(1'h0)])
                begin
                  for (forvar4188 = (1'h0); (forvar4188 < (2'h3)); forvar4188 = (forvar4188 + (1'h1)))
                    begin
                      reg4189 <= reg4088;
                      reg4190 <= $signed(((8'ha7) < {(reg4094 <= (8'ha7))}));
                      reg4191 <= wire3720;
                    end
                  reg4192 <= (|(!$unsigned({(8'ha5)})));
                  for (forvar4193 = (1'h0); (forvar4193 < (2'h3)); forvar4193 = (forvar4193 + (1'h1)))
                    begin
                      reg4194 <= $unsigned((~^(|(~^reg4055))));
                    end
                end
              else
                begin
                  for (forvar4188 = (1'h0); (forvar4188 < (2'h3)); forvar4188 = (forvar4188 + (1'h1)))
                    begin
                      reg4189 <= (^$signed(reg4106));
                      reg4190 <= ({(reg3993 << forvar4104)} & $unsigned((~^reg4114[(2'h2):(1'h1)])));
                    end
                  for (forvar4191 = (1'h0); (forvar4191 < (1'h1)); forvar4191 = (forvar4191 + (1'h1)))
                    begin
                      reg4192 <= $signed({(-reg3842)});
                      reg4193 <= $unsigned($signed(($unsigned(wire5) > ((8'hba) <= wire4096))));
                      reg4194 <= (reg4194 ?
                          $signed((!$signed(reg3781))) : $signed((~|(forvar4193 - reg4148))));
                    end
                  if (reg4193)
                    begin
                      reg4195 <= reg3785[(2'h2):(1'h0)];
                      reg4196 <= reg75[(4'h8):(3'h5)];
                      reg4197 <= (({(reg49 ? forvar4188 : (8'hac))} ?
                          reg3800[(4'he):(1'h1)] : reg4032[(2'h3):(1'h0)]) + (reg3942 >= ((reg3873 < (8'hb7)) ?
                          ((8'ha5) ? reg3855 : wire8) : (~^reg83))));
                    end
                  else
                    begin
                      reg4195 <= $unsigned($unsigned($unsigned($signed(reg4004))));
                      reg4196 <= ({wire3632} ? reg4089 : (8'h9e));
                      reg4197 <= ($signed(reg3737) & {(8'ha9)});
                    end
                end
              reg4198 <= (+({(reg67 || (8'ha5))} >>> ($unsigned(reg4192) && ((8'hb0) ^ reg4068))));
              for (forvar4199 = (1'h0); (forvar4199 < (1'h0)); forvar4199 = (forvar4199 + (1'h1)))
                begin
                  if (reg31)
                    begin
                      reg4200 <= reg3730;
                    end
                  else
                    begin
                      reg4200 <= ((reg3717[(3'h6):(2'h3)] >>> ((reg3858 >>> reg3863) != reg3983[(1'h1):(1'h0)])) ?
                          (!((reg4055 >> reg4198) & (reg3729 || forvar4191))) : (((reg4069 - forvar4138) ^ (reg3891 ^~ reg17)) == $signed($signed(reg3909))));
                      reg4201 <= $signed(reg4171);
                      reg4202 <= reg4112;
                    end
                  if (($signed($unsigned(((8'hb0) && reg3906))) ?
                      $signed((|{reg4127})) : {{(reg3748 ?
                                  reg3824 : reg3874)}}))
                    begin
                      reg4203 <= ((&(^~{reg4094})) ^ $unsigned((reg3979 >>> reg3816[(1'h0):(1'h0)])));
                      reg4204 <= ((($signed(reg3802) ?
                              reg3976[(2'h2):(2'h2)] : (|reg3771)) - reg3808) ?
                          $signed(reg83) : reg3799);
                    end
                  else
                    begin
                      reg4203 <= (8'hae);
                      reg4204 <= $signed($unsigned($signed(reg3969[(4'h8):(3'h5)])));
                      reg4205 <= (8'hab);
                      reg4206 <= $unsigned($unsigned((reg3939 ?
                          reg3936 : $unsigned(reg34))));
                    end
                end
              if ($unsigned(reg4068))
                begin
                  for (forvar4207 = (1'h0); (forvar4207 < (2'h2)); forvar4207 = (forvar4207 + (1'h1)))
                    begin
                      reg4208 <= $unsigned($unsigned((~^$signed((8'haf)))));
                      reg4209 <= (reg3880[(3'h6):(3'h5)] ?
                          (-(reg3684 ?
                              wire4097[(1'h0):(1'h0)] : (~reg3965))) : $unsigned((~&reg3687[(4'hc):(4'hc)])));
                      reg4210 <= reg3941;
                      reg4211 <= reg3973[(1'h0):(1'h0)];
                    end
                  for (forvar4212 = (1'h0); (forvar4212 < (1'h0)); forvar4212 = (forvar4212 + (1'h1)))
                    begin
                      reg4213 <= {$signed($unsigned((~^(8'h9e))))};
                    end
                end
              else
                begin
                  if ($signed($unsigned(($signed(reg4172) ?
                      {forvar4108} : reg4104[(4'hc):(4'hc)]))))
                    begin
                      reg4207 <= $signed(reg4152[(1'h0):(1'h0)]);
                      reg4208 <= (8'hac);
                      reg4209 <= ({$signed((&reg3859))} > $unsigned($signed((reg31 | reg4160))));
                      reg4210 <= ((-reg3824) ?
                          {reg49} : (~^(((8'h9e) ^ reg46) || (~reg3709))));
                    end
                  else
                    begin
                      reg4207 <= reg3766;
                    end
                  reg4211 <= (($unsigned(((8'hac) | forvar4113)) ?
                          reg27[(4'hc):(1'h1)] : (+(reg4128 > reg3989))) ?
                      reg3674[(2'h2):(1'h0)] : wire4097[(2'h2):(1'h1)]);
                  for (forvar4212 = (1'h0); (forvar4212 < (2'h2)); forvar4212 = (forvar4212 + (1'h1)))
                    begin
                      reg4213 <= (~&($signed(reg3743[(1'h1):(1'h0)]) ?
                          reg3825[(4'hb):(3'h5)] : reg3704));
                      reg4214 <= reg4206[(2'h3):(2'h3)];
                    end
                end
            end
          else
            begin
              for (forvar4188 = (1'h0); (forvar4188 < (2'h3)); forvar4188 = (forvar4188 + (1'h1)))
                begin
                  if ($unsigned(reg4030[(3'h5):(1'h1)]))
                    begin
                      reg4189 <= (8'ha1);
                      reg4190 <= (8'hb9);
                      reg4191 <= reg3801[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg4189 <= reg4001;
                      reg4190 <= ((~&(((8'ha1) ?
                              (8'haa) : reg3701) ^ (wire3632 ?
                              reg3818 : reg3715))) ?
                          (reg4049 ?
                              ($signed(reg4078) ?
                                  $unsigned((8'h9c)) : reg4051[(3'h7):(2'h3)]) : reg3809) : reg24);
                      reg4191 <= ((8'h9d) <<< reg3986);
                      reg4192 <= reg4053;
                    end
                  if (reg3939[(2'h3):(1'h0)])
                    begin
                      reg4193 <= $unsigned(reg50);
                      reg4194 <= ((reg4007[(4'hd):(3'h4)] >>> reg4117) ?
                          ($signed(reg4184[(2'h2):(1'h0)]) - reg3745[(3'h6):(3'h5)]) : (^~reg3639));
                      reg4195 <= $signed((reg4148 > ((^~reg3662) ^~ {(8'ha2)})));
                    end
                  else
                    begin
                      reg4193 <= reg3850[(3'h6):(3'h6)];
                      reg4194 <= (~((^~(8'ha0)) ?
                          ((reg3701 ?
                              reg3941 : reg3940) - $unsigned(reg3839)) : (^(reg4055 ?
                              reg3701 : reg57))));
                    end
                  for (forvar4196 = (1'h0); (forvar4196 < (2'h3)); forvar4196 = (forvar4196 + (1'h1)))
                    begin
                      reg4197 <= (~|reg3988);
                      reg4198 <= ($unsigned($signed((8'h9e))) >>> ((8'h9e) ?
                          $signed((^~reg4116)) : ((reg4204 || reg28) - (reg4013 << reg4065))));
                    end
                  for (forvar4199 = (1'h0); (forvar4199 < (1'h0)); forvar4199 = (forvar4199 + (1'h1)))
                    begin
                      reg4200 <= (((&(|reg3669)) && reg3840[(4'hc):(4'hc)]) << $unsigned($unsigned($unsigned(reg3662))));
                      reg4201 <= reg3687[(4'ha):(2'h2)];
                      reg4202 <= ((reg4017 * ((reg3924 <<< (8'hab)) == $unsigned(reg4159))) > $signed(($signed(reg3857) >> reg3652[(3'h6):(2'h3)])));
                      reg4203 <= $signed((($unsigned(reg3961) ?
                          (reg4126 ?
                              reg4009 : wire3721) : {reg3940}) > $signed((8'ha4))));
                    end
                end
              if ($unsigned(reg3877[(1'h1):(1'h1)]))
                begin
                  if ((^~(~^reg4043[(3'h5):(1'h0)])))
                    begin
                      reg4204 <= reg4101;
                      reg4205 <= $unsigned((!forvar4101));
                      reg4206 <= (reg3763[(3'h5):(2'h2)] ^ ((reg4017[(2'h2):(1'h1)] ?
                          $signed(reg3902) : reg3880) >> {$signed(forvar4132)}));
                      reg4207 <= ($signed(($unsigned((8'ha2)) - $signed(reg4116))) & $unsigned(($unsigned(reg3967) ?
                          (!(8'hb2)) : $unsigned(forvar4196))));
                    end
                  else
                    begin
                      reg4204 <= (reg3726[(1'h1):(1'h0)] << $unsigned(((reg3730 ^~ reg63) ?
                          reg84[(3'h6):(2'h2)] : (!forvar4188))));
                      reg4205 <= (^((8'h9f) <= ($unsigned(reg3666) * reg4182[(4'h9):(2'h2)])));
                    end
                  for (forvar4208 = (1'h0); (forvar4208 < (1'h0)); forvar4208 = (forvar4208 + (1'h1)))
                    begin
                      reg4209 <= $signed((8'haf));
                      reg4210 <= (((~^$signed(reg3899)) ?
                              ($unsigned(reg3832) ^ (!reg3943)) : (-((8'h9d) ?
                                  (8'hb3) : reg3958))) ?
                          (((forvar4120 ? reg3639 : reg3876) ?
                              (forvar4102 - reg4151) : $signed(wire3919)) & ($signed(forvar4147) >>> (reg4069 ?
                              reg4059 : reg3859))) : (-$unsigned({reg3673})));
                      reg4211 <= (($signed($unsigned(reg4182)) ^ $unsigned($unsigned(reg3704))) ?
                          $unsigned($unsigned((reg3814 ^ reg4122))) : $signed(reg3641));
                      reg4212 <= $unsigned((({reg3805} == $unsigned((8'h9e))) << ($unsigned(forvar4138) ~^ (|(8'haa)))));
                    end
                end
              else
                begin
                  if ((forvar4212 & {$unsigned(((8'hb4) ? reg3936 : reg4187))}))
                    begin
                      reg4204 <= ($signed(reg3722[(1'h0):(1'h0)]) ?
                          ((wire7 ?
                                  (+reg3694) : (reg3948 ? (8'ha4) : reg4065)) ?
                              {reg3731} : $signed((reg3933 ^ reg3979))) : (^~({reg3750} ?
                              $signed(reg3747) : (reg3938 ?
                                  reg4124 : reg3962))));
                      reg4205 <= $signed((reg3690 >>> $signed(reg4086)));
                      reg4206 <= forvar4199[(4'h8):(3'h4)];
                    end
                  else
                    begin
                      reg4204 <= $signed((($signed(reg4019) >= (8'hb9)) ?
                          (~(forvar4193 ~^ reg4173)) : ($unsigned(reg3990) == (~|reg46))));
                    end
                  for (forvar4207 = (1'h0); (forvar4207 < (2'h2)); forvar4207 = (forvar4207 + (1'h1)))
                    begin
                      reg4208 <= (($unsigned((reg3952 ? reg4178 : forvar4177)) ?
                              (^(reg3772 || reg3693)) : {(wire4099 << reg4063)}) ?
                          forvar4191[(4'hc):(3'h7)] : $unsigned(reg3748));
                    end
                end
              for (forvar4213 = (1'h0); (forvar4213 < (1'h1)); forvar4213 = (forvar4213 + (1'h1)))
                begin
                  reg4214 <= (+reg3673);
                  reg4215 <= $unsigned(($unsigned((+(8'hb3))) == reg3724[(2'h3):(1'h0)]));
                  for (forvar4216 = (1'h0); (forvar4216 < (1'h1)); forvar4216 = (forvar4216 + (1'h1)))
                    begin
                      reg4217 <= reg3844[(4'he):(4'he)];
                      reg4218 <= (($unsigned((&reg4118)) | (&(~reg3806))) + $signed($unsigned($unsigned(reg3956))));
                    end
                  for (forvar4219 = (1'h0); (forvar4219 < (2'h2)); forvar4219 = (forvar4219 + (1'h1)))
                    begin
                      reg4220 <= (((((8'ha1) >= reg3704) ?
                              $unsigned(reg4125) : {reg3788}) ?
                          ($signed(reg3673) + $unsigned(reg3733)) : reg3794) ^~ ({$unsigned(reg3781)} ?
                          $signed($unsigned(forvar4132)) : (~&reg3954[(4'hb):(3'h5)])));
                      reg4221 <= (({(~^forvar4154)} ?
                          reg4134[(3'h7):(3'h5)] : reg76) && reg4130[(1'h0):(1'h0)]);
                    end
                end
              if ({((reg3806[(3'h5):(2'h3)] + (^reg3989)) >= reg3727)})
                begin
                  for (forvar4222 = (1'h0); (forvar4222 < (1'h1)); forvar4222 = (forvar4222 + (1'h1)))
                    begin
                      reg4223 <= reg3724[(1'h1):(1'h0)];
                      reg4224 <= $signed(reg13);
                    end
                  for (forvar4225 = (1'h0); (forvar4225 < (1'h0)); forvar4225 = (forvar4225 + (1'h1)))
                    begin
                      reg4226 <= {((^(-reg4049)) < reg3805[(3'h4):(1'h0)])};
                      reg4227 <= {(^$unsigned($signed(reg3761)))};
                    end
                end
              else
                begin
                  if ($signed(reg3812))
                    begin
                      reg4222 <= $unsigned($signed(reg4034[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg4222 <= reg4192[(3'h6):(3'h5)];
                      reg4223 <= {$unsigned(reg3871[(2'h2):(1'h0)])};
                      reg4224 <= $unsigned(reg44[(1'h0):(1'h0)]);
                      reg4225 <= {(((8'ha5) + (-(8'hb6))) && reg52)};
                    end
                  reg4226 <= reg4017[(1'h0):(1'h0)];
                  if ((($unsigned((reg3955 ?
                          reg3717 : wire3721)) ~^ wire4096[(3'h4):(1'h1)]) ?
                      (($signed(reg4124) ?
                          (^(8'ha5)) : (-reg3665)) == $unsigned($signed(reg3724))) : ((reg81[(3'h5):(3'h5)] ?
                          reg3766[(1'h0):(1'h0)] : {reg3665}) + $unsigned((reg3979 ?
                          forvar4177 : (8'hb3))))))
                    begin
                      reg4227 <= $signed(reg3941[(4'hc):(3'h5)]);
                      reg4228 <= reg3987;
                      reg4229 <= (8'ha3);
                      reg4230 <= reg4075[(3'h6):(3'h4)];
                    end
                  else
                    begin
                      reg4227 <= $unsigned((((+reg3878) >> $unsigned(reg4213)) ?
                          (~(reg22 ? reg3796 : (8'hb3))) : (|(reg3679 ?
                              reg3698 : reg4212))));
                      reg4228 <= reg4092[(1'h0):(1'h0)];
                      reg4229 <= wire3632[(3'h6):(3'h6)];
                    end
                  if (reg3699[(4'hb):(2'h3)])
                    begin
                      reg4231 <= ({((reg3966 ^ reg3981) == reg3858)} < $unsigned(reg3985[(3'h4):(2'h2)]));
                      reg4232 <= (((~&(reg3712 <<< reg3983)) ?
                              $signed($signed(reg40)) : (reg3911[(3'h4):(1'h0)] ?
                                  (wire5 ?
                                      reg3948 : reg3661) : $unsigned(reg74))) ?
                          {(8'ha7)} : (((reg4108 ? reg4051 : reg4204) ?
                                  reg3973 : reg3769) ?
                              reg3771 : $signed(reg3730)));
                    end
                  else
                    begin
                      reg4231 <= reg3830[(1'h0):(1'h0)];
                      reg4232 <= reg3830[(2'h3):(2'h3)];
                      reg4233 <= (reg3912[(2'h3):(1'h0)] >>> reg3940);
                      reg4234 <= ($unsigned(({reg4046} ~^ ((8'h9d) ?
                              reg4116 : forvar4207))) ?
                          (reg4175[(3'h6):(3'h6)] <<< $signed(reg3846[(4'ha):(3'h4)])) : (|$unsigned((reg4095 < (8'hac)))));
                    end
                end
            end
          if ({(8'hab)})
            begin
              for (forvar4235 = (1'h0); (forvar4235 < (1'h1)); forvar4235 = (forvar4235 + (1'h1)))
                begin
                  reg4236 <= $unsigned(((!reg4220[(2'h2):(1'h1)]) ?
                      $signed((!wire4096)) : (~&(!reg3883))));
                  for (forvar4237 = (1'h0); (forvar4237 < (2'h2)); forvar4237 = (forvar4237 + (1'h1)))
                    begin
                      reg4238 <= $unsigned((wire7[(3'h5):(1'h1)] ?
                          reg4179 : ($unsigned(reg4150) ?
                              reg3911[(3'h4):(1'h0)] : reg3815[(1'h1):(1'h0)])));
                    end
                  for (forvar4239 = (1'h0); (forvar4239 < (2'h3)); forvar4239 = (forvar4239 + (1'h1)))
                    begin
                      reg4240 <= ((|(reg4201 ? {reg3876} : (!reg3984))) ?
                          reg4030 : ((reg3791 ?
                              reg3810[(1'h1):(1'h1)] : wire4098) && $unsigned((reg3872 ?
                              (8'hb1) : reg3990))));
                      reg4241 <= (reg4026[(4'hc):(4'h8)] ?
                          ((|reg19[(2'h2):(2'h2)]) ?
                              (reg3879[(1'h1):(1'h1)] - $signed(reg81)) : reg3832[(4'ha):(3'h7)]) : (~(~$signed(reg3808))));
                      reg4242 <= $unsigned((^~$unsigned({reg4086})));
                      reg4243 <= reg4027[(2'h3):(2'h2)];
                    end
                  if (wire7)
                    begin
                      reg4244 <= $unsigned(reg46);
                      reg4245 <= (8'hab);
                      reg4246 <= ((($unsigned(reg3917) || ((8'ha2) | (8'ha4))) ?
                              $unsigned((reg3859 ?
                                  reg3674 : reg4001)) : reg3730[(3'h6):(2'h3)]) ?
                          reg3995[(2'h2):(1'h0)] : $unsigned(({reg3771} ^ (8'hb3))));
                      reg4247 <= {$signed(($unsigned(reg19) >> (^(8'ha8))))};
                    end
                  else
                    begin
                      reg4244 <= reg3700;
                      reg4245 <= $signed(($signed($unsigned(reg25)) ^~ (~|$unsigned(reg3656))));
                      reg4246 <= reg3993;
                    end
                end
              for (forvar4248 = (1'h0); (forvar4248 < (1'h1)); forvar4248 = (forvar4248 + (1'h1)))
                begin
                  for (forvar4249 = (1'h0); (forvar4249 < (1'h1)); forvar4249 = (forvar4249 + (1'h1)))
                    begin
                      reg4250 <= ($signed((+(wire4097 ?
                          forvar4235 : (8'ha5)))) > ($unsigned(forvar4249) ?
                          reg3837[(1'h1):(1'h0)] : (8'hb0)));
                      reg4251 <= reg3886;
                    end
                  for (forvar4252 = (1'h0); (forvar4252 < (1'h1)); forvar4252 = (forvar4252 + (1'h1)))
                    begin
                      reg4253 <= {$signed((~^reg4225))};
                    end
                  if ((~reg3848))
                    begin
                      reg4254 <= ((~(8'hb5)) >= reg4167[(2'h3):(2'h3)]);
                      reg4255 <= $unsigned(forvar4115[(4'ha):(4'ha)]);
                      reg4256 <= $unsigned((~|$signed((reg3863 ?
                          reg4214 : forvar4252))));
                      reg4257 <= $signed((reg3667 ?
                          ((^reg45) >= $unsigned(reg4038)) : reg3649));
                    end
                  else
                    begin
                      reg4254 <= $unsigned((-reg4157[(3'h4):(1'h1)]));
                    end
                end
            end
          else
            begin
              for (forvar4235 = (1'h0); (forvar4235 < (1'h0)); forvar4235 = (forvar4235 + (1'h1)))
                begin
                  reg4236 <= ($unsigned(($signed(reg3991) ?
                          (~&(8'ha8)) : (reg3739 > (8'hab)))) ?
                      {$unsigned(reg4134)} : (!reg3701));
                  for (forvar4237 = (1'h0); (forvar4237 < (1'h0)); forvar4237 = (forvar4237 + (1'h1)))
                    begin
                      reg4238 <= reg3726[(4'ha):(3'h5)];
                      reg4239 <= $unsigned((!reg3728));
                      reg4240 <= reg3650;
                    end
                  for (forvar4241 = (1'h0); (forvar4241 < (2'h2)); forvar4241 = (forvar4241 + (1'h1)))
                    begin
                      reg4242 <= $signed((!reg4233));
                      reg4243 <= $signed((reg3977[(3'h4):(1'h1)] || reg4242));
                    end
                  if ((^~(($signed(reg4196) ?
                      $unsigned((8'hb3)) : (forvar4191 | reg4244)) > ({reg4203} > (reg3662 ~^ reg3823)))))
                    begin
                      reg4244 <= reg34;
                      reg4245 <= $signed($signed(($unsigned(reg4253) ?
                          ((8'ha4) == (8'h9e)) : (~|wire4099))));
                      reg4246 <= $signed(reg3753[(3'h5):(1'h1)]);
                    end
                  else
                    begin
                      reg4244 <= $signed(({reg3954} > $unsigned(((8'ha0) - reg3763))));
                      reg4245 <= (~^(reg3685[(4'hb):(1'h1)] ?
                          reg4134 : forvar4131));
                      reg4246 <= (8'hb4);
                      reg4247 <= reg3941[(3'h6):(2'h3)];
                    end
                end
              if (reg4157[(1'h0):(1'h0)])
                begin
                  if ($unsigned($signed($unsigned((^~reg4242)))))
                    begin
                      reg4248 <= ({$signed((forvar4207 ? reg43 : (8'ha4)))} ?
                          reg3805[(3'h4):(1'h0)] : (!((!reg3841) ?
                              (reg3704 ?
                                  reg3690 : (8'ha6)) : ((8'ha9) <= reg4204))));
                    end
                  else
                    begin
                      reg4248 <= $signed(($signed({reg4021}) ?
                          reg3683[(2'h2):(1'h0)] : reg4105[(3'h5):(1'h1)]));
                      reg4249 <= (($unsigned(reg3696) ?
                          $signed((reg4105 - reg4160)) : reg3978) << reg4070[(4'hf):(2'h2)]);
                    end
                  reg4250 <= ((!$signed((|reg3998))) ?
                      forvar4107[(2'h3):(1'h0)] : (-(~^reg3818)));
                end
              else
                begin
                  reg4248 <= reg4007;
                end
              reg4251 <= $unsigned($unsigned($signed((wire7 & reg3701))));
              for (forvar4252 = (1'h0); (forvar4252 < (1'h0)); forvar4252 = (forvar4252 + (1'h1)))
                begin
                  for (forvar4253 = (1'h0); (forvar4253 < (1'h1)); forvar4253 = (forvar4253 + (1'h1)))
                    begin
                      reg4254 <= ($signed($unsigned(reg3757)) >= ((8'h9f) ^~ ($unsigned((8'ha5)) != {(8'ha5)})));
                      reg4255 <= $signed(reg3874[(4'h8):(3'h7)]);
                      reg4256 <= {$unsigned({$signed(reg3849)})};
                      reg4257 <= {forvar4119[(2'h2):(1'h1)]};
                    end
                  if ((reg4172[(4'hb):(3'h5)] < ($signed(reg3728) + ({reg3751} ?
                      (reg3810 - reg4056) : reg3909))))
                    begin
                      reg4258 <= $unsigned(reg3828);
                    end
                  else
                    begin
                      reg4258 <= reg3653;
                      reg4259 <= (~(((|reg4034) ?
                          (reg3652 ?
                              reg3719 : reg3846) : {reg3678}) * ($signed(reg4137) ?
                          (-(8'ha2)) : reg4136)));
                      reg4260 <= (reg3835 ?
                          (-reg4166) : $unsigned($unsigned(reg3659)));
                      reg4261 <= (+reg4089);
                    end
                end
            end
        end
      for (forvar4262 = (1'h0); (forvar4262 < (1'h1)); forvar4262 = (forvar4262 + (1'h1)))
        begin
          for (forvar4263 = (1'h0); (forvar4263 < (2'h3)); forvar4263 = (forvar4263 + (1'h1)))
            begin
              for (forvar4264 = (1'h0); (forvar4264 < (2'h2)); forvar4264 = (forvar4264 + (1'h1)))
                begin
                  reg4265 <= $signed($signed((reg4046 ?
                      (reg3818 != forvar4219) : (reg4070 - reg3815))));
                end
              for (forvar4266 = (1'h0); (forvar4266 < (2'h2)); forvar4266 = (forvar4266 + (1'h1)))
                begin
                  for (forvar4267 = (1'h0); (forvar4267 < (1'h1)); forvar4267 = (forvar4267 + (1'h1)))
                    begin
                      reg4268 <= (((&(^reg4180)) ?
                              reg3996[(4'ha):(3'h7)] : (reg70[(3'h6):(1'h0)] + {forvar4196})) ?
                          reg4169 : (&reg3859));
                    end
                  for (forvar4269 = (1'h0); (forvar4269 < (1'h0)); forvar4269 = (forvar4269 + (1'h1)))
                    begin
                      reg4270 <= $signed($unsigned($signed({reg3878})));
                      reg4271 <= $signed($signed(((|(8'hb5)) ^~ (8'ha2))));
                    end
                end
              if (($signed(forvar4105[(3'h5):(3'h4)]) > $unsigned(((-(8'hb8)) ^~ (|reg3844)))))
                begin
                  if ($signed(reg4183))
                    begin
                      reg4272 <= (reg3937[(4'ha):(2'h2)] >>> reg4242[(1'h0):(1'h0)]);
                      reg4273 <= $unsigned(reg3814);
                      reg4274 <= ((8'haa) ? reg3924 : (~&$signed((~^reg3766))));
                      reg4275 <= $signed({{(-reg4265)}});
                    end
                  else
                    begin
                      reg4272 <= ((((~reg4039) ?
                              $signed((8'hb7)) : $signed(reg4271)) ?
                          (~^(~reg3637)) : $unsigned((forvar4262 ?
                              (8'h9d) : (8'hb5)))) | (reg4114[(2'h3):(2'h2)] ~^ ((reg4163 <= forvar4168) > {reg3965})));
                      reg4273 <= ($unsigned((reg4049[(4'h9):(3'h5)] ?
                          (forvar4103 ?
                              reg3848 : reg3912) : reg3951[(2'h3):(1'h0)])) >= (-reg3761[(1'h0):(1'h0)]));
                    end
                  for (forvar4276 = (1'h0); (forvar4276 < (2'h2)); forvar4276 = (forvar4276 + (1'h1)))
                    begin
                      reg4277 <= reg3912[(4'hc):(3'h5)];
                      reg4278 <= (&((-(^reg3767)) ?
                          ((!reg3884) ?
                              (^~reg4074) : (~forvar4252)) : (-((8'ha3) ?
                              reg4070 : reg3661))));
                      reg4279 <= (($unsigned((reg4141 ?
                              reg3989 : reg3709)) | reg4242[(3'h4):(2'h3)]) ?
                          (((reg3849 || (8'hb3)) ?
                              $unsigned(reg3681) : (reg3879 >> wire3636)) ~^ reg3863[(3'h7):(2'h2)]) : reg4064[(1'h1):(1'h0)]);
                      reg4280 <= $unsigned((-$signed((reg4170 ?
                          reg3845 : reg3832))));
                    end
                end
              else
                begin
                  if (reg77[(4'ha):(4'h9)])
                    begin
                      reg4272 <= (^~reg3841[(4'he):(4'he)]);
                      reg4273 <= $unsigned((^$unsigned((8'hba))));
                      reg4274 <= ((&reg3657[(1'h1):(1'h0)]) ?
                          {$signed(reg4170[(3'h4):(1'h1)])} : reg4231[(3'h5):(3'h5)]);
                    end
                  else
                    begin
                      reg4272 <= $signed((+(^~(^~reg3669))));
                    end
                  reg4275 <= ($signed($unsigned($unsigned(reg3644))) & $unsigned((((8'h9c) ~^ reg4196) && $signed(reg3848))));
                  for (forvar4276 = (1'h0); (forvar4276 < (2'h3)); forvar4276 = (forvar4276 + (1'h1)))
                    begin
                      reg4277 <= (reg20[(2'h3):(2'h2)] && {$signed((reg3730 & reg4017))});
                      reg4278 <= (reg3667 <<< reg3844[(3'h5):(1'h0)]);
                    end
                end
            end
          reg4281 <= ((+(8'hb1)) ? {(^~reg25)} : reg4250[(3'h6):(1'h1)]);
          for (forvar4282 = (1'h0); (forvar4282 < (1'h0)); forvar4282 = (forvar4282 + (1'h1)))
            begin
              if ((($signed((~reg4006)) ?
                  reg3661 : ((8'hb2) || (reg4021 && (8'ha0)))) <= (&(|reg4109[(1'h1):(1'h1)]))))
                begin
                  for (forvar4283 = (1'h0); (forvar4283 < (2'h3)); forvar4283 = (forvar4283 + (1'h1)))
                    begin
                      reg4284 <= (reg4277 > (~&$signed((8'hab))));
                      reg4285 <= (((reg3894[(4'hb):(2'h2)] ?
                              reg3675 : reg3966) < reg14[(3'h4):(2'h3)]) ?
                          $signed(reg3990) : $signed($unsigned($unsigned(reg4095))));
                    end
                  for (forvar4286 = (1'h0); (forvar4286 < (1'h0)); forvar4286 = (forvar4286 + (1'h1)))
                    begin
                      reg4287 <= reg3654[(3'h6):(2'h2)];
                      reg4288 <= $signed($unsigned((+((8'hb4) ^~ reg3745))));
                    end
                  reg4289 <= reg3858;
                end
              else
                begin
                  if (reg4247)
                    begin
                      reg4283 <= (({(reg45 ?
                              reg3962 : reg4181)} <<< $signed((reg4190 - reg3696))) != (~((reg3925 >>> (8'ha5)) ?
                          (reg3937 ?
                              reg3791 : (8'ha5)) : $signed(forvar4155))));
                      reg4284 <= ($signed($unsigned((^reg3950))) ?
                          forvar4102 : (~&($unsigned(reg27) + reg3878)));
                      reg4285 <= {$signed({$signed(reg4238)})};
                    end
                  else
                    begin
                      reg4283 <= $unsigned((reg71 - reg4016[(1'h0):(1'h0)]));
                      reg4284 <= reg3972;
                      reg4285 <= $unsigned(((~&reg3698[(3'h7):(1'h1)]) + $signed((~reg4118))));
                      reg4286 <= (reg4084 ?
                          ($signed(reg3810) ?
                              $unsigned((reg3880 ?
                                  reg3797 : (8'h9d))) : $signed($unsigned((8'hb2)))) : $unsigned(reg4222));
                    end
                  reg4287 <= (($unsigned($unsigned((8'ha8))) ?
                      reg3832[(4'he):(4'h9)] : reg73) == $signed($unsigned((-(8'hb4)))));
                  if ($signed(reg3897))
                    begin
                      reg4288 <= $unsigned($signed(($unsigned(reg4275) ?
                          $unsigned((8'h9f)) : $unsigned(reg4283))));
                      reg4289 <= reg4139;
                    end
                  else
                    begin
                      reg4288 <= reg4160[(4'h9):(4'h8)];
                      reg4289 <= reg4106[(3'h6):(3'h4)];
                      reg4290 <= reg4170[(2'h2):(1'h0)];
                      reg4291 <= forvar4120;
                    end
                  for (forvar4292 = (1'h0); (forvar4292 < (1'h0)); forvar4292 = (forvar4292 + (1'h1)))
                    begin
                      reg4293 <= (^~(|$unsigned((reg18 >>> reg4006))));
                      reg4294 <= (^reg4173);
                      reg4295 <= {$signed(reg3826[(3'h4):(1'h1)])};
                    end
                end
              reg4296 <= {(((reg3832 ? reg3968 : reg4215) ?
                      reg3879[(2'h3):(1'h0)] : reg3934[(4'ha):(1'h0)]) <<< $signed($signed(reg4174)))};
            end
          for (forvar4297 = (1'h0); (forvar4297 < (2'h2)); forvar4297 = (forvar4297 + (1'h1)))
            begin
              if ($unsigned($signed(reg4056)))
                begin
                  reg4298 <= (8'hb7);
                  reg4299 <= (8'hb9);
                  reg4300 <= $signed(({$unsigned(reg4071)} ?
                      (|(^reg3940)) : $signed(reg3853)));
                  if (((&$signed(reg37[(2'h2):(1'h0)])) ?
                      ($signed({reg4206}) ?
                          reg3652[(2'h3):(1'h1)] : reg4169) : $unsigned(((forvar4178 ?
                              (8'hb0) : reg4289) ?
                          reg4104[(4'ha):(3'h7)] : reg3718[(2'h3):(1'h1)]))))
                    begin
                      reg4301 <= $unsigned($signed({reg4005[(4'hc):(3'h5)]}));
                    end
                  else
                    begin
                      reg4301 <= $unsigned((reg4248 ^ reg3778));
                      reg4302 <= reg3658[(3'h6):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar4298 = (1'h0); (forvar4298 < (2'h3)); forvar4298 = (forvar4298 + (1'h1)))
                    begin
                      reg4299 <= (reg3983[(1'h1):(1'h1)] ^~ reg3852);
                    end
                end
              for (forvar4303 = (1'h0); (forvar4303 < (2'h2)); forvar4303 = (forvar4303 + (1'h1)))
                begin
                  if (($unsigned($signed((forvar4168 ? reg3823 : wire6))) ?
                      ((&$signed(reg3993)) ?
                          ((reg3748 <<< forvar4123) ^ $signed(reg3749)) : {reg3837[(2'h3):(1'h1)]}) : ($unsigned(forvar4132) ?
                          {reg3858} : $signed((wire3632 ? reg4068 : reg3699)))))
                    begin
                      reg4304 <= reg4260[(4'hd):(4'hb)];
                    end
                  else
                    begin
                      reg4304 <= $unsigned((reg72 ?
                          (reg4053[(2'h2):(2'h2)] < $unsigned((8'haa))) : $signed((reg3828 ?
                              reg4043 : reg3966))));
                      reg4305 <= (reg4165 ?
                          $unsigned(((^~reg3667) ?
                              (reg3988 <<< reg3647) : {forvar4193})) : reg3639[(3'h7):(2'h2)]);
                      reg4306 <= (8'haa);
                      reg4307 <= $unsigned({{(~(8'ha4))}});
                    end
                  for (forvar4308 = (1'h0); (forvar4308 < (1'h0)); forvar4308 = (forvar4308 + (1'h1)))
                    begin
                      reg4309 <= $signed((((^~reg3645) > (reg4247 ?
                          wire4097 : reg4180)) * $unsigned((reg4201 >>> reg4020))));
                      reg4310 <= (|((^(8'ha2)) == (reg3757[(2'h3):(2'h2)] && $unsigned(reg4253))));
                    end
                  for (forvar4311 = (1'h0); (forvar4311 < (1'h0)); forvar4311 = (forvar4311 + (1'h1)))
                    begin
                      reg4312 <= $unsigned(reg4165[(2'h3):(2'h2)]);
                      reg4313 <= reg34[(2'h2):(2'h2)];
                      reg4314 <= (!(((reg3905 ?
                          reg4116 : (8'hb8)) >>> {reg4242}) < $unsigned((reg3903 ?
                          reg3839 : reg4256))));
                    end
                end
            end
        end
      reg4315 <= reg4301;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module86
#(parameter param3631 = (8'ha1))
(y, clk, wire90, wire89, wire88, wire87);
  output wire [(32'h1085):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire90;
  input wire signed [(3'h4):(1'h0)] wire89;
  input wire [(3'h5):(1'h0)] wire88;
  input wire signed [(4'h8):(1'h0)] wire87;
  wire [(3'h7):(1'h0)] wire3629;
  wire signed [(4'ha):(1'h0)] wire721;
  wire signed [(4'hb):(1'h0)] wire720;
  wire [(4'h9):(1'h0)] wire718;
  wire signed [(4'h8):(1'h0)] wire512;
  wire signed [(3'h6):(1'h0)] wire511;
  wire [(5'h10):(1'h0)] wire510;
  wire signed [(3'h4):(1'h0)] wire93;
  wire [(3'h6):(1'h0)] wire92;
  wire signed [(3'h5):(1'h0)] wire91;
  reg signed [(3'h6):(1'h0)] reg509 = (1'h0);
  reg [(4'h9):(1'h0)] reg508 = (1'h0);
  reg [(4'h9):(1'h0)] reg507 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg506 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg505 = (1'h0);
  reg [(4'he):(1'h0)] reg504 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg503 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg502 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg501 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg500 = (1'h0);
  reg [(4'hc):(1'h0)] reg499 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg498 = (1'h0);
  reg [(3'h7):(1'h0)] reg497 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg496 = (1'h0);
  reg [(2'h3):(1'h0)] reg495 = (1'h0);
  reg [(4'hd):(1'h0)] reg494 = (1'h0);
  reg [(4'hc):(1'h0)] reg493 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg488 = (1'h0);
  reg [(2'h2):(1'h0)] reg492 = (1'h0);
  reg [(5'h10):(1'h0)] reg491 = (1'h0);
  reg [(4'hc):(1'h0)] reg490 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg489 = (1'h0);
  reg [(4'h8):(1'h0)] reg486 = (1'h0);
  reg [(3'h4):(1'h0)] reg485 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg484 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg483 = (1'h0);
  reg [(4'he):(1'h0)] reg482 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg480 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg479 = (1'h0);
  reg [(4'he):(1'h0)] reg478 = (1'h0);
  reg [(4'he):(1'h0)] reg477 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg475 = (1'h0);
  reg signed [(4'he):(1'h0)] reg474 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg473 = (1'h0);
  reg [(2'h3):(1'h0)] reg470 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg469 = (1'h0);
  reg [(4'h8):(1'h0)] reg466 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg462 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg468 = (1'h0);
  reg [(4'h8):(1'h0)] reg467 = (1'h0);
  reg [(3'h4):(1'h0)] reg465 = (1'h0);
  reg [(4'hb):(1'h0)] reg464 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg463 = (1'h0);
  reg [(4'hd):(1'h0)] reg461 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg459 = (1'h0);
  reg [(2'h2):(1'h0)] reg458 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg457 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg456 = (1'h0);
  reg [(4'h9):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg452 = (1'h0);
  reg [(2'h3):(1'h0)] reg451 = (1'h0);
  reg [(4'hd):(1'h0)] reg450 = (1'h0);
  reg [(3'h6):(1'h0)] reg449 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg447 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg446 = (1'h0);
  reg [(4'h9):(1'h0)] reg445 = (1'h0);
  reg [(4'hf):(1'h0)] reg444 = (1'h0);
  reg [(5'h10):(1'h0)] reg443 = (1'h0);
  reg [(4'hc):(1'h0)] reg441 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg440 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg439 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg438 = (1'h0);
  reg [(4'hd):(1'h0)] reg437 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg436 = (1'h0);
  reg [(3'h6):(1'h0)] reg435 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg434 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg430 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg427 = (1'h0);
  reg [(2'h2):(1'h0)] reg426 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg425 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg424 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg422 = (1'h0);
  reg [(2'h2):(1'h0)] reg421 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg420 = (1'h0);
  reg [(5'h10):(1'h0)] reg419 = (1'h0);
  reg [(3'h6):(1'h0)] reg418 = (1'h0);
  reg [(3'h4):(1'h0)] reg417 = (1'h0);
  reg [(2'h2):(1'h0)] reg416 = (1'h0);
  reg [(4'h9):(1'h0)] reg414 = (1'h0);
  reg [(4'h8):(1'h0)] reg413 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg412 = (1'h0);
  reg [(3'h4):(1'h0)] reg409 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg408 = (1'h0);
  reg [(4'hf):(1'h0)] reg407 = (1'h0);
  reg [(4'hf):(1'h0)] reg406 = (1'h0);
  reg [(5'h10):(1'h0)] reg404 = (1'h0);
  reg [(4'hb):(1'h0)] reg402 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg401 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg400 = (1'h0);
  reg [(4'hf):(1'h0)] reg399 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg397 = (1'h0);
  reg signed [(4'he):(1'h0)] reg396 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg393 = (1'h0);
  reg [(4'hd):(1'h0)] reg392 = (1'h0);
  reg [(4'h9):(1'h0)] reg391 = (1'h0);
  reg [(3'h4):(1'h0)] reg390 = (1'h0);
  reg [(3'h4):(1'h0)] reg389 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg388 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg386 = (1'h0);
  reg [(4'hd):(1'h0)] reg385 = (1'h0);
  reg [(4'h8):(1'h0)] reg384 = (1'h0);
  reg [(3'h7):(1'h0)] reg383 = (1'h0);
  reg [(5'h10):(1'h0)] reg380 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg378 = (1'h0);
  reg [(2'h3):(1'h0)] reg377 = (1'h0);
  reg [(4'hd):(1'h0)] reg376 = (1'h0);
  reg [(3'h5):(1'h0)] reg375 = (1'h0);
  reg [(4'hc):(1'h0)] reg374 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg373 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg363 = (1'h0);
  reg [(3'h7):(1'h0)] reg362 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg358 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg356 = (1'h0);
  reg [(4'h9):(1'h0)] reg351 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg371 = (1'h0);
  reg signed [(4'he):(1'h0)] reg370 = (1'h0);
  reg [(4'h9):(1'h0)] reg369 = (1'h0);
  reg [(4'h8):(1'h0)] reg368 = (1'h0);
  reg [(4'hb):(1'h0)] reg367 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg366 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg365 = (1'h0);
  reg [(4'h9):(1'h0)] reg364 = (1'h0);
  reg [(4'hd):(1'h0)] reg361 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg360 = (1'h0);
  reg [(3'h5):(1'h0)] reg359 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg357 = (1'h0);
  reg [(3'h6):(1'h0)] reg355 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg354 = (1'h0);
  reg [(4'hf):(1'h0)] reg353 = (1'h0);
  reg signed [(4'he):(1'h0)] reg350 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg349 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg348 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg345 = (1'h0);
  reg [(4'he):(1'h0)] reg347 = (1'h0);
  reg [(2'h2):(1'h0)] reg346 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg344 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg343 = (1'h0);
  reg [(3'h5):(1'h0)] reg342 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg341 = (1'h0);
  reg signed [(4'he):(1'h0)] reg339 = (1'h0);
  reg [(3'h4):(1'h0)] reg338 = (1'h0);
  reg [(4'h9):(1'h0)] reg337 = (1'h0);
  reg [(4'he):(1'h0)] reg336 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg334 = (1'h0);
  reg [(5'h10):(1'h0)] reg333 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg332 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg331 = (1'h0);
  reg [(4'h9):(1'h0)] reg330 = (1'h0);
  reg [(3'h4):(1'h0)] reg329 = (1'h0);
  reg [(4'hb):(1'h0)] reg328 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg327 = (1'h0);
  reg [(4'ha):(1'h0)] reg324 = (1'h0);
  reg [(3'h4):(1'h0)] reg323 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg322 = (1'h0);
  reg [(3'h4):(1'h0)] reg321 = (1'h0);
  reg [(4'ha):(1'h0)] reg320 = (1'h0);
  reg [(4'ha):(1'h0)] reg318 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg319 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg317 = (1'h0);
  reg [(5'h10):(1'h0)] reg316 = (1'h0);
  reg [(4'hd):(1'h0)] reg315 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg314 = (1'h0);
  reg [(2'h2):(1'h0)] reg313 = (1'h0);
  reg [(2'h2):(1'h0)] reg311 = (1'h0);
  reg [(3'h7):(1'h0)] reg310 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg304 = (1'h0);
  reg [(4'he):(1'h0)] reg292 = (1'h0);
  reg [(3'h5):(1'h0)] reg287 = (1'h0);
  reg [(3'h6):(1'h0)] reg284 = (1'h0);
  reg [(3'h4):(1'h0)] reg283 = (1'h0);
  reg [(4'hd):(1'h0)] reg303 = (1'h0);
  reg [(5'h10):(1'h0)] reg302 = (1'h0);
  reg [(4'ha):(1'h0)] reg301 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg300 = (1'h0);
  reg [(4'hb):(1'h0)] reg299 = (1'h0);
  reg [(4'ha):(1'h0)] reg296 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg295 = (1'h0);
  reg [(2'h2):(1'h0)] reg294 = (1'h0);
  reg [(3'h5):(1'h0)] reg293 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg291 = (1'h0);
  reg [(4'hd):(1'h0)] reg290 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg289 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg288 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg286 = (1'h0);
  reg [(4'h8):(1'h0)] reg285 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg278 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg274 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg272 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg282 = (1'h0);
  reg [(4'he):(1'h0)] reg281 = (1'h0);
  reg [(4'hf):(1'h0)] reg280 = (1'h0);
  reg [(2'h2):(1'h0)] reg279 = (1'h0);
  reg [(4'he):(1'h0)] reg277 = (1'h0);
  reg [(3'h7):(1'h0)] reg276 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg275 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg273 = (1'h0);
  reg [(4'ha):(1'h0)] reg271 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg270 = (1'h0);
  reg [(3'h7):(1'h0)] reg269 = (1'h0);
  reg [(4'hd):(1'h0)] reg268 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg267 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg264 = (1'h0);
  reg [(4'h8):(1'h0)] reg263 = (1'h0);
  reg [(5'h10):(1'h0)] reg262 = (1'h0);
  reg [(4'hb):(1'h0)] reg261 = (1'h0);
  reg [(4'h8):(1'h0)] reg260 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg258 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg256 = (1'h0);
  reg [(4'hc):(1'h0)] reg255 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg254 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg253 = (1'h0);
  reg [(3'h4):(1'h0)] reg252 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg250 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg249 = (1'h0);
  reg [(4'hc):(1'h0)] reg248 = (1'h0);
  reg [(2'h2):(1'h0)] reg247 = (1'h0);
  reg [(4'h8):(1'h0)] reg246 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg244 = (1'h0);
  reg [(3'h7):(1'h0)] reg243 = (1'h0);
  reg [(4'hf):(1'h0)] reg242 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg241 = (1'h0);
  reg [(4'hd):(1'h0)] reg240 = (1'h0);
  reg [(4'hf):(1'h0)] reg239 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg238 = (1'h0);
  reg [(4'hb):(1'h0)] reg237 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg236 = (1'h0);
  reg [(4'ha):(1'h0)] reg234 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg233 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg232 = (1'h0);
  reg [(4'hd):(1'h0)] reg231 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg219 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg229 = (1'h0);
  reg [(4'hf):(1'h0)] reg227 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg226 = (1'h0);
  reg [(4'hb):(1'h0)] reg225 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg223 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg222 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg221 = (1'h0);
  reg [(4'h9):(1'h0)] reg220 = (1'h0);
  reg [(3'h4):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg217 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg216 = (1'h0);
  reg [(4'hd):(1'h0)] reg215 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg213 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg212 = (1'h0);
  reg [(5'h10):(1'h0)] reg211 = (1'h0);
  reg [(4'hb):(1'h0)] reg209 = (1'h0);
  reg [(2'h3):(1'h0)] reg208 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg207 = (1'h0);
  reg [(3'h4):(1'h0)] reg205 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg204 = (1'h0);
  reg [(5'h10):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg202 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg201 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg200 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg199 = (1'h0);
  reg [(4'hf):(1'h0)] reg198 = (1'h0);
  reg [(4'h9):(1'h0)] reg197 = (1'h0);
  reg [(2'h2):(1'h0)] reg196 = (1'h0);
  reg [(5'h10):(1'h0)] reg195 = (1'h0);
  reg [(2'h2):(1'h0)] reg194 = (1'h0);
  reg [(4'h9):(1'h0)] reg193 = (1'h0);
  reg [(4'hc):(1'h0)] reg192 = (1'h0);
  reg [(3'h6):(1'h0)] reg191 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg187 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg186 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg185 = (1'h0);
  reg signed [(4'he):(1'h0)] reg184 = (1'h0);
  reg [(5'h10):(1'h0)] reg183 = (1'h0);
  reg signed [(4'he):(1'h0)] reg182 = (1'h0);
  reg [(3'h5):(1'h0)] reg180 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg178 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg177 = (1'h0);
  reg [(3'h4):(1'h0)] reg176 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg175 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg174 = (1'h0);
  reg [(4'hc):(1'h0)] reg172 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg171 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg169 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg168 = (1'h0);
  reg [(4'h8):(1'h0)] reg167 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg166 = (1'h0);
  reg [(4'hc):(1'h0)] reg165 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg160 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg157 = (1'h0);
  reg [(4'hd):(1'h0)] reg156 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg155 = (1'h0);
  reg [(4'h8):(1'h0)] reg154 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg153 = (1'h0);
  reg [(3'h7):(1'h0)] reg148 = (1'h0);
  reg [(4'hc):(1'h0)] reg147 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg146 = (1'h0);
  reg [(4'hc):(1'h0)] reg145 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg144 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg143 = (1'h0);
  reg signed [(4'he):(1'h0)] reg142 = (1'h0);
  reg [(4'ha):(1'h0)] reg141 = (1'h0);
  reg [(3'h6):(1'h0)] reg140 = (1'h0);
  reg [(5'h10):(1'h0)] reg139 = (1'h0);
  reg [(3'h7):(1'h0)] reg138 = (1'h0);
  reg signed [(4'he):(1'h0)] reg136 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg135 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg134 = (1'h0);
  reg [(2'h3):(1'h0)] reg131 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg129 = (1'h0);
  reg [(4'h8):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg127 = (1'h0);
  reg [(4'h8):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg125 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg124 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg123 = (1'h0);
  reg [(3'h5):(1'h0)] reg122 = (1'h0);
  reg [(4'he):(1'h0)] reg121 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg118 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg117 = (1'h0);
  reg [(4'hb):(1'h0)] reg116 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg115 = (1'h0);
  reg [(4'hc):(1'h0)] reg114 = (1'h0);
  reg [(2'h2):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg112 = (1'h0);
  reg signed [(4'he):(1'h0)] reg111 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg110 = (1'h0);
  reg [(4'hf):(1'h0)] reg109 = (1'h0);
  reg [(3'h7):(1'h0)] reg107 = (1'h0);
  reg [(2'h3):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg104 = (1'h0);
  reg [(4'hf):(1'h0)] reg103 = (1'h0);
  reg [(4'hf):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg100 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg99 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg98 = (1'h0);
  reg [(3'h6):(1'h0)] reg97 = (1'h0);
  reg [(4'h9):(1'h0)] forvar506 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar496 = (1'h0);
  reg [(2'h2):(1'h0)] forvar488 = (1'h0);
  reg [(5'h10):(1'h0)] forvar487 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar481 = (1'h0);
  reg [(3'h6):(1'h0)] forvar476 = (1'h0);
  reg [(4'hb):(1'h0)] forvar472 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar471 = (1'h0);
  reg [(2'h2):(1'h0)] forvar467 = (1'h0);
  reg [(4'he):(1'h0)] forvar465 = (1'h0);
  reg [(4'hd):(1'h0)] forvar466 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar462 = (1'h0);
  reg [(4'h9):(1'h0)] forvar460 = (1'h0);
  reg [(4'hd):(1'h0)] forvar455 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar453 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar445 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar448 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar442 = (1'h0);
  reg [(4'h8):(1'h0)] forvar433 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar432 = (1'h0);
  reg [(2'h2):(1'h0)] forvar431 = (1'h0);
  reg [(4'hb):(1'h0)] forvar429 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar428 = (1'h0);
  reg [(2'h2):(1'h0)] forvar423 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar415 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar411 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar410 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar405 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar403 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar398 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar395 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar394 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar389 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar387 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar382 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar381 = (1'h0);
  reg [(4'ha):(1'h0)] forvar372 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar371 = (1'h0);
  reg [(4'hd):(1'h0)] forvar370 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar364 = (1'h0);
  reg [(4'h9):(1'h0)] forvar350 = (1'h0);
  reg [(4'hf):(1'h0)] forvar344 = (1'h0);
  reg [(3'h7):(1'h0)] forvar341 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar363 = (1'h0);
  reg [(2'h3):(1'h0)] forvar362 = (1'h0);
  reg [(3'h5):(1'h0)] forvar358 = (1'h0);
  reg [(3'h5):(1'h0)] forvar356 = (1'h0);
  reg [(4'he):(1'h0)] forvar352 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar351 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar345 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar340 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar289 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar335 = (1'h0);
  reg [(3'h5):(1'h0)] forvar326 = (1'h0);
  reg [(4'hf):(1'h0)] forvar325 = (1'h0);
  reg [(2'h2):(1'h0)] forvar318 = (1'h0);
  reg [(2'h2):(1'h0)] forvar312 = (1'h0);
  reg [(4'hf):(1'h0)] forvar309 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar307 = (1'h0);
  reg [(4'h9):(1'h0)] forvar306 = (1'h0);
  reg [(2'h3):(1'h0)] forvar305 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar293 = (1'h0);
  reg [(3'h7):(1'h0)] forvar285 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar281 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar298 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar297 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar292 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar287 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar284 = (1'h0);
  reg [(3'h7):(1'h0)] forvar283 = (1'h0);
  reg [(2'h2):(1'h0)] forvar276 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar271 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar278 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar274 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar272 = (1'h0);
  reg [(4'hc):(1'h0)] forvar266 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar265 = (1'h0);
  reg [(4'he):(1'h0)] forvar259 = (1'h0);
  reg [(4'hb):(1'h0)] forvar257 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar245 = (1'h0);
  reg [(5'h10):(1'h0)] forvar242 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar235 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar230 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar217 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar228 = (1'h0);
  reg [(3'h6):(1'h0)] forvar224 = (1'h0);
  reg [(3'h4):(1'h0)] forvar219 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar214 = (1'h0);
  reg [(4'hb):(1'h0)] forvar210 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar206 = (1'h0);
  reg [(5'h10):(1'h0)] forvar190 = (1'h0);
  reg [(4'he):(1'h0)] forvar189 = (1'h0);
  reg [(2'h2):(1'h0)] forvar188 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar181 = (1'h0);
  reg [(4'ha):(1'h0)] forvar179 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar173 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar170 = (1'h0);
  reg [(3'h7):(1'h0)] forvar164 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar163 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar161 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar158 = (1'h0);
  reg [(3'h6):(1'h0)] forvar152 = (1'h0);
  reg [(3'h4):(1'h0)] forvar151 = (1'h0);
  reg [(4'hd):(1'h0)] forvar150 = (1'h0);
  reg [(4'hc):(1'h0)] forvar149 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar137 = (1'h0);
  reg [(4'hf):(1'h0)] forvar133 = (1'h0);
  reg [(3'h4):(1'h0)] forvar132 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar130 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar120 = (1'h0);
  reg [(2'h2):(1'h0)] forvar119 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar110 = (1'h0);
  reg [(3'h6):(1'h0)] forvar108 = (1'h0);
  reg [(4'he):(1'h0)] forvar106 = (1'h0);
  reg [(4'ha):(1'h0)] forvar99 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar102 = (1'h0);
  reg [(3'h4):(1'h0)] forvar96 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar95 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar94 = (1'h0);
  assign y = {wire3629,
                 wire721,
                 wire720,
                 wire718,
                 wire512,
                 wire511,
                 wire510,
                 wire93,
                 wire92,
                 wire91,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg488,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg480,
                 reg479,
                 reg478,
                 reg477,
                 reg475,
                 reg474,
                 reg473,
                 reg470,
                 reg469,
                 reg466,
                 reg462,
                 reg468,
                 reg467,
                 reg465,
                 reg464,
                 reg463,
                 reg461,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg454,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg447,
                 reg446,
                 reg445,
                 reg444,
                 reg443,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg430,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg414,
                 reg413,
                 reg412,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg404,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg397,
                 reg396,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg363,
                 reg362,
                 reg358,
                 reg356,
                 reg351,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg361,
                 reg360,
                 reg359,
                 reg357,
                 reg355,
                 reg354,
                 reg353,
                 reg350,
                 reg349,
                 reg348,
                 reg345,
                 reg347,
                 reg346,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg318,
                 reg319,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg311,
                 reg310,
                 reg308,
                 reg304,
                 reg292,
                 reg287,
                 reg284,
                 reg283,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg286,
                 reg285,
                 reg278,
                 reg274,
                 reg272,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg277,
                 reg276,
                 reg275,
                 reg273,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg258,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg219,
                 reg229,
                 reg227,
                 reg226,
                 reg225,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg213,
                 reg212,
                 reg211,
                 reg209,
                 reg208,
                 reg207,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg180,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg172,
                 reg171,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg162,
                 reg160,
                 reg159,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg136,
                 reg135,
                 reg134,
                 reg131,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg107,
                 reg105,
                 reg104,
                 reg103,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 forvar506,
                 forvar496,
                 forvar488,
                 forvar487,
                 forvar481,
                 forvar476,
                 forvar472,
                 forvar471,
                 forvar467,
                 forvar465,
                 forvar466,
                 forvar462,
                 forvar460,
                 forvar455,
                 forvar453,
                 forvar445,
                 forvar448,
                 forvar442,
                 forvar433,
                 forvar432,
                 forvar431,
                 forvar429,
                 forvar428,
                 forvar423,
                 forvar415,
                 forvar411,
                 forvar410,
                 forvar405,
                 forvar403,
                 forvar398,
                 forvar395,
                 forvar394,
                 forvar389,
                 forvar387,
                 forvar382,
                 forvar381,
                 forvar372,
                 forvar371,
                 forvar370,
                 forvar364,
                 forvar350,
                 forvar344,
                 forvar341,
                 forvar363,
                 forvar362,
                 forvar358,
                 forvar356,
                 forvar352,
                 forvar351,
                 forvar345,
                 forvar340,
                 forvar289,
                 forvar335,
                 forvar326,
                 forvar325,
                 forvar318,
                 forvar312,
                 forvar309,
                 forvar307,
                 forvar306,
                 forvar305,
                 forvar293,
                 forvar285,
                 forvar281,
                 forvar298,
                 forvar297,
                 forvar292,
                 forvar287,
                 forvar284,
                 forvar283,
                 forvar276,
                 forvar271,
                 forvar278,
                 forvar274,
                 forvar272,
                 forvar266,
                 forvar265,
                 forvar259,
                 forvar257,
                 forvar245,
                 forvar242,
                 forvar235,
                 forvar230,
                 forvar217,
                 forvar228,
                 forvar224,
                 forvar219,
                 forvar214,
                 forvar210,
                 forvar206,
                 forvar190,
                 forvar189,
                 forvar188,
                 forvar181,
                 forvar179,
                 forvar173,
                 forvar170,
                 forvar164,
                 forvar163,
                 forvar161,
                 forvar158,
                 forvar152,
                 forvar151,
                 forvar150,
                 forvar149,
                 forvar137,
                 forvar133,
                 forvar132,
                 forvar130,
                 forvar120,
                 forvar119,
                 forvar110,
                 forvar108,
                 forvar106,
                 forvar99,
                 forvar102,
                 forvar96,
                 forvar95,
                 forvar94,
                 (1'h0)};
  assign wire91 = {{$signed($unsigned(wire87))}};
  assign wire92 = $signed((~wire91[(1'h1):(1'h1)]));
  assign wire93 = wire88[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar94 = (1'h0); (forvar94 < (1'h0)); forvar94 = (forvar94 + (1'h1)))
        begin
          for (forvar95 = (1'h0); (forvar95 < (1'h0)); forvar95 = (forvar95 + (1'h1)))
            begin
              for (forvar96 = (1'h0); (forvar96 < (1'h0)); forvar96 = (forvar96 + (1'h1)))
                begin
                  reg97 <= ((-(-(~^wire91))) & wire89[(2'h3):(2'h3)]);
                end
              if ($unsigned((8'haa)))
                begin
                  if ((forvar95 || $signed(forvar94)))
                    begin
                      reg98 <= wire91;
                      reg99 <= $signed($signed((8'ha3)));
                      reg100 <= ((|($unsigned(wire91) == (wire92 ^~ wire88))) == $signed(((|wire87) ?
                          (forvar96 ?
                              wire87 : wire91) : forvar96[(1'h1):(1'h1)])));
                      reg101 <= $unsigned(((forvar96 >= reg97) ?
                          $unsigned(reg97) : wire93[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg98 <= wire88;
                      reg99 <= (8'hb5);
                      reg100 <= $unsigned(wire93);
                    end
                  for (forvar102 = (1'h0); (forvar102 < (2'h3)); forvar102 = (forvar102 + (1'h1)))
                    begin
                      reg103 <= {$signed($signed((forvar95 ?
                              wire89 : reg101)))};
                      reg104 <= $unsigned(($unsigned((reg99 ?
                          reg103 : reg100)) < $signed({reg99})));
                      reg105 <= $signed(((reg101 ?
                          forvar94[(1'h0):(1'h0)] : (wire92 + reg101)) - $unsigned((forvar96 || wire88))));
                    end
                end
              else
                begin
                  reg98 <= (&(reg101[(3'h7):(1'h0)] ?
                      (~$unsigned(wire92)) : {reg97}));
                  for (forvar99 = (1'h0); (forvar99 < (1'h1)); forvar99 = (forvar99 + (1'h1)))
                    begin
                      reg100 <= {reg100[(2'h3):(1'h1)]};
                    end
                end
              for (forvar106 = (1'h0); (forvar106 < (1'h1)); forvar106 = (forvar106 + (1'h1)))
                begin
                  reg107 <= wire93[(2'h3):(2'h2)];
                  for (forvar108 = (1'h0); (forvar108 < (1'h0)); forvar108 = (forvar108 + (1'h1)))
                    begin
                      reg109 <= $signed(wire90);
                    end
                end
            end
          if (($signed((~&$signed(forvar102))) >> $signed(wire93)))
            begin
              reg110 <= reg97;
            end
          else
            begin
              for (forvar110 = (1'h0); (forvar110 < (1'h1)); forvar110 = (forvar110 + (1'h1)))
                begin
                  reg111 <= (~(8'had));
                  if ((reg98[(4'h8):(3'h6)] ?
                      wire87 : ({{reg103}} ? reg100 : reg101[(4'h8):(2'h2)])))
                    begin
                      reg112 <= (~(((8'h9e) || (8'hb1)) ?
                          reg100[(3'h6):(3'h6)] : (^(forvar108 ?
                              reg103 : (8'ha3)))));
                      reg113 <= $unsigned((|(wire88 ?
                          $unsigned(reg99) : $unsigned(reg111))));
                      reg114 <= (~|wire90);
                      reg115 <= ($unsigned({((8'hb3) < reg98)}) ?
                          $unsigned($signed(reg111[(3'h6):(3'h5)])) : ({$signed(reg101)} ?
                              forvar95 : ($signed((8'hb6)) * wire89)));
                    end
                  else
                    begin
                      reg112 <= $unsigned((+(|(^forvar106))));
                    end
                  reg116 <= {$signed(wire88[(3'h4):(1'h1)])};
                end
              reg117 <= ((|reg101) >> ($unsigned((~wire87)) || (wire88[(2'h2):(2'h2)] ?
                  (reg114 ? forvar108 : reg107) : (forvar110 >> reg104))));
              reg118 <= ((((!reg111) * {forvar106}) ?
                      $signed(reg97) : (reg98 ? {reg99} : reg116)) ?
                  $unsigned($signed(reg99[(2'h2):(1'h0)])) : ((~^reg100[(2'h3):(1'h1)]) + reg109[(3'h6):(2'h2)]));
              for (forvar119 = (1'h0); (forvar119 < (1'h1)); forvar119 = (forvar119 + (1'h1)))
                begin
                  for (forvar120 = (1'h0); (forvar120 < (1'h0)); forvar120 = (forvar120 + (1'h1)))
                    begin
                      reg121 <= reg103;
                      reg122 <= reg114;
                      reg123 <= reg114[(4'h8):(4'h8)];
                    end
                  if (((((wire93 ?
                      reg107 : (8'h9d)) != $signed(forvar102)) && $unsigned((forvar96 ?
                      forvar95 : forvar108))) ~^ ((^~reg121) ?
                      (-reg112[(3'h4):(2'h3)]) : forvar106)))
                    begin
                      reg124 <= (reg118 ?
                          $unsigned(forvar106[(4'h8):(3'h5)]) : $unsigned(forvar102));
                    end
                  else
                    begin
                      reg124 <= reg123[(1'h0):(1'h0)];
                      reg125 <= {$unsigned(reg97)};
                      reg126 <= $unsigned(reg125);
                      reg127 <= (~$unsigned($unsigned(((8'ha4) ?
                          reg115 : reg104))));
                    end
                  reg128 <= ((forvar106[(4'hb):(3'h6)] && {$signed(wire93)}) ^ {reg117});
                  reg129 <= (reg117 > wire91[(3'h5):(3'h5)]);
                end
            end
          for (forvar130 = (1'h0); (forvar130 < (1'h0)); forvar130 = (forvar130 + (1'h1)))
            begin
              reg131 <= (+$signed($unsigned((forvar96 ? reg104 : forvar94))));
              for (forvar132 = (1'h0); (forvar132 < (2'h3)); forvar132 = (forvar132 + (1'h1)))
                begin
                  for (forvar133 = (1'h0); (forvar133 < (1'h1)); forvar133 = (forvar133 + (1'h1)))
                    begin
                      reg134 <= forvar108;
                      reg135 <= (forvar119[(1'h1):(1'h1)] ?
                          (~|reg105[(2'h3):(2'h2)]) : forvar95[(4'h9):(3'h5)]);
                      reg136 <= forvar95;
                    end
                  for (forvar137 = (1'h0); (forvar137 < (1'h1)); forvar137 = (forvar137 + (1'h1)))
                    begin
                      reg138 <= $unsigned(wire92[(1'h1):(1'h0)]);
                      reg139 <= (reg136[(2'h2):(1'h1)] < $signed((+reg113[(1'h0):(1'h0)])));
                    end
                  if ($signed(reg97[(3'h5):(3'h4)]))
                    begin
                      reg140 <= forvar108[(2'h3):(2'h2)];
                      reg141 <= ((forvar133 ?
                              {(forvar120 && forvar95)} : $unsigned(reg127[(4'hf):(4'hb)])) ?
                          (&(~^{reg111})) : (~wire90[(1'h1):(1'h0)]));
                      reg142 <= reg109;
                    end
                  else
                    begin
                      reg140 <= {(forvar108 > (reg126 == {reg135}))};
                      reg141 <= $signed({($signed(reg124) ?
                              (reg118 ? reg124 : reg128) : $unsigned(reg131))});
                    end
                  if ($signed($unsigned($unsigned($unsigned(reg118)))))
                    begin
                      reg143 <= reg136[(1'h0):(1'h0)];
                      reg144 <= reg107[(3'h7):(3'h7)];
                      reg145 <= reg97;
                      reg146 <= forvar130;
                    end
                  else
                    begin
                      reg143 <= reg139;
                      reg144 <= (|reg116[(4'h8):(4'h8)]);
                      reg145 <= {{$signed(reg113)}};
                    end
                end
            end
        end
      reg147 <= reg100[(4'hc):(4'hc)];
      reg148 <= (((|(reg136 ? wire87 : reg140)) + $signed(forvar94)) ?
          $signed(reg109) : $unsigned(reg134[(3'h7):(1'h1)]));
    end
  always
    @(posedge clk) begin
      for (forvar149 = (1'h0); (forvar149 < (2'h2)); forvar149 = (forvar149 + (1'h1)))
        begin
          for (forvar150 = (1'h0); (forvar150 < (1'h1)); forvar150 = (forvar150 + (1'h1)))
            begin
              for (forvar151 = (1'h0); (forvar151 < (1'h0)); forvar151 = (forvar151 + (1'h1)))
                begin
                  for (forvar152 = (1'h0); (forvar152 < (2'h2)); forvar152 = (forvar152 + (1'h1)))
                    begin
                      reg153 <= reg107[(3'h5):(1'h0)];
                      reg154 <= (forvar149 <<< $unsigned($unsigned((reg104 || (8'haf)))));
                      reg155 <= ($signed(reg125[(3'h5):(1'h1)]) - reg125[(1'h1):(1'h1)]);
                      reg156 <= (((&(reg140 ?
                              forvar150 : forvar151)) ^~ ({reg114} ?
                              $unsigned((8'haa)) : wire90[(3'h4):(2'h2)])) ?
                          reg107 : (~|(!(reg118 && wire87))));
                    end
                  reg157 <= (8'ha9);
                  for (forvar158 = (1'h0); (forvar158 < (1'h0)); forvar158 = (forvar158 + (1'h1)))
                    begin
                      reg159 <= (~^(^~$unsigned((8'ha0))));
                      reg160 <= reg155;
                    end
                  for (forvar161 = (1'h0); (forvar161 < (2'h2)); forvar161 = (forvar161 + (1'h1)))
                    begin
                      reg162 <= ($signed(($signed(reg138) ?
                              reg114[(3'h5):(3'h4)] : reg109[(4'hd):(2'h3)])) ?
                          (8'ha6) : reg143);
                    end
                end
              for (forvar163 = (1'h0); (forvar163 < (1'h1)); forvar163 = (forvar163 + (1'h1)))
                begin
                  for (forvar164 = (1'h0); (forvar164 < (2'h2)); forvar164 = (forvar164 + (1'h1)))
                    begin
                      reg165 <= $unsigned({reg113});
                      reg166 <= $unsigned(((|{reg104}) ?
                          $signed((|(8'hb7))) : $signed(((8'ha1) ?
                              reg115 : forvar158))));
                    end
                  if (reg114[(4'h8):(3'h5)])
                    begin
                      reg167 <= ((((reg124 ? reg100 : reg118) ~^ (^~reg129)) ?
                              {reg124} : $unsigned(reg156)) ?
                          forvar152 : ({reg112} ^~ ($signed((8'ha7)) && $signed((8'ha3)))));
                      reg168 <= ($signed((8'hac)) ~^ ((^$unsigned((8'ha5))) | $unsigned($signed(reg98))));
                    end
                  else
                    begin
                      reg167 <= $unsigned(($signed(((8'ha6) ?
                              forvar163 : reg154)) ?
                          {(reg99 ? reg141 : reg117)} : (reg144 ?
                              $signed(reg127) : (reg128 < reg159))));
                    end
                  reg169 <= (({$signed(reg131)} <<< (&$signed(reg136))) ?
                      ((&$signed(reg101)) ?
                          reg113[(1'h0):(1'h0)] : (((8'ha3) > (8'hb6)) <<< reg118)) : $signed((reg100 - $unsigned(reg146))));
                  for (forvar170 = (1'h0); (forvar170 < (1'h1)); forvar170 = (forvar170 + (1'h1)))
                    begin
                      reg171 <= (~$unsigned(($unsigned(reg101) ?
                          $signed(reg136) : reg118[(2'h2):(1'h0)])));
                      reg172 <= (|(-($unsigned(reg112) ^~ $unsigned(reg126))));
                    end
                end
              for (forvar173 = (1'h0); (forvar173 < (2'h3)); forvar173 = (forvar173 + (1'h1)))
                begin
                  reg174 <= ((((^reg97) && (~forvar170)) << reg128) ?
                      reg112 : (((reg141 & reg131) ?
                              ((8'hb9) > reg99) : $signed(wire92)) ?
                          $unsigned((wire90 >>> reg146)) : $signed(wire87[(3'h5):(3'h5)])));
                  if (forvar149[(3'h6):(1'h0)])
                    begin
                      reg175 <= (+(reg101 ?
                          wire92[(3'h5):(1'h1)] : {((8'ha7) ?
                                  (8'had) : reg156)}));
                      reg176 <= $signed($unsigned($unsigned($unsigned(forvar151))));
                    end
                  else
                    begin
                      reg175 <= (8'h9c);
                      reg176 <= forvar158[(1'h1):(1'h1)];
                      reg177 <= $signed(reg111[(2'h2):(1'h1)]);
                      reg178 <= reg156[(4'h8):(3'h4)];
                    end
                end
              if (reg177)
                begin
                  for (forvar179 = (1'h0); (forvar179 < (1'h0)); forvar179 = (forvar179 + (1'h1)))
                    begin
                      reg180 <= ($unsigned((~{(8'h9e)})) > (|reg174));
                    end
                  for (forvar181 = (1'h0); (forvar181 < (1'h1)); forvar181 = (forvar181 + (1'h1)))
                    begin
                      reg182 <= wire87;
                      reg183 <= reg156;
                      reg184 <= ((|($unsigned(reg114) > (reg116 ?
                          reg172 : reg138))) <<< $signed($unsigned(reg180[(1'h1):(1'h0)])));
                    end
                  if ((+(reg145 ?
                      ((reg146 ^ (8'ha1)) >= $signed(reg155)) : {$unsigned(reg117)})))
                    begin
                      reg185 <= $signed($unsigned(reg143));
                      reg186 <= reg180;
                    end
                  else
                    begin
                      reg185 <= (8'ha0);
                      reg186 <= reg113[(2'h2):(1'h1)];
                      reg187 <= (-(|(reg116 >= (reg142 & (8'hba)))));
                    end
                end
              else
                begin
                  for (forvar179 = (1'h0); (forvar179 < (1'h1)); forvar179 = (forvar179 + (1'h1)))
                    begin
                      reg180 <= reg182[(1'h1):(1'h1)];
                    end
                  for (forvar181 = (1'h0); (forvar181 < (1'h1)); forvar181 = (forvar181 + (1'h1)))
                    begin
                      reg182 <= (({$unsigned(wire91)} ?
                          $signed((8'hb7)) : (reg110 ^~ $signed(reg136))) | ($unsigned(reg121[(2'h3):(1'h1)]) ?
                          reg168[(1'h1):(1'h0)] : ((forvar173 ?
                              reg169 : (8'h9d)) != $unsigned(reg171))));
                      reg183 <= ($signed(reg138) ^ ((reg180[(2'h3):(1'h1)] ~^ (~&forvar181)) << (reg144[(1'h0):(1'h0)] ?
                          forvar150 : $signed((8'hb6)))));
                      reg184 <= reg153;
                      reg185 <= wire91[(2'h2):(1'h0)];
                    end
                end
            end
          for (forvar188 = (1'h0); (forvar188 < (2'h2)); forvar188 = (forvar188 + (1'h1)))
            begin
              for (forvar189 = (1'h0); (forvar189 < (1'h0)); forvar189 = (forvar189 + (1'h1)))
                begin
                  for (forvar190 = (1'h0); (forvar190 < (2'h2)); forvar190 = (forvar190 + (1'h1)))
                    begin
                      reg191 <= reg116[(3'h5):(2'h3)];
                      reg192 <= $signed(($unsigned((!reg169)) ?
                          reg172[(1'h1):(1'h1)] : $unsigned($unsigned(reg186))));
                      reg193 <= reg176;
                    end
                  if (reg104)
                    begin
                      reg194 <= $signed(reg171);
                    end
                  else
                    begin
                      reg194 <= ((reg111 * ((|forvar152) ^ {reg178})) ?
                          $signed((^(~reg126))) : $signed((~|(wire91 < reg129))));
                      reg195 <= (^~(((reg184 ?
                          forvar181 : (8'ha1)) ~^ reg127[(5'h10):(3'h4)]) ^~ (~|forvar188)));
                      reg196 <= (~&(~&$unsigned((^reg169))));
                      reg197 <= $unsigned(($unsigned($signed(reg162)) >> ({(8'hb1)} ?
                          $unsigned(reg104) : $signed((8'h9e)))));
                    end
                  if (((((reg175 < forvar181) != $signed(reg113)) > ({(8'ha2)} ?
                          (forvar189 < reg99) : $signed(reg192))) ?
                      $unsigned((~&reg174[(3'h5):(3'h5)])) : {forvar163}))
                    begin
                      reg198 <= reg172[(4'hb):(3'h4)];
                      reg199 <= $signed($unsigned($signed($unsigned(wire92))));
                      reg200 <= forvar163;
                    end
                  else
                    begin
                      reg198 <= $unsigned($unsigned($signed(reg142)));
                      reg199 <= (~|reg136);
                    end
                end
              reg201 <= ((reg175 << {(|reg107)}) ?
                  reg196[(2'h2):(2'h2)] : reg200[(1'h0):(1'h0)]);
              reg202 <= reg97[(3'h5):(3'h4)];
              if ((reg117[(3'h4):(1'h0)] ? forvar151 : reg111[(3'h7):(3'h4)]))
                begin
                  if ($unsigned($signed(reg144[(4'h8):(3'h5)])))
                    begin
                      reg203 <= (((reg187 - (&(8'ha1))) ?
                          $unsigned(wire91[(1'h1):(1'h0)]) : reg104) + ((|(reg109 ?
                              reg121 : reg191)) ?
                          $signed(reg136[(4'hb):(1'h1)]) : (~^{reg140})));
                      reg204 <= (!$unsigned($unsigned((reg169 ^~ (8'haf)))));
                      reg205 <= (+$unsigned(wire91));
                    end
                  else
                    begin
                      reg203 <= forvar179;
                      reg204 <= {(8'hab)};
                      reg205 <= (~^({(reg178 ? reg144 : reg141)} ?
                          $signed(wire93[(2'h3):(2'h3)]) : ((^reg100) ^~ (reg141 | reg198))));
                    end
                  for (forvar206 = (1'h0); (forvar206 < (2'h3)); forvar206 = (forvar206 + (1'h1)))
                    begin
                      reg207 <= ((-(+(8'hb2))) - forvar188);
                      reg208 <= (($unsigned((reg186 ? wire89 : reg197)) ?
                              (^~{(8'ha2)}) : (reg113 ^~ {reg160})) ?
                          forvar188[(2'h2):(2'h2)] : (!reg136));
                      reg209 <= $signed($signed(forvar181[(3'h7):(3'h4)]));
                    end
                  for (forvar210 = (1'h0); (forvar210 < (1'h1)); forvar210 = (forvar210 + (1'h1)))
                    begin
                      reg211 <= $signed(reg187[(2'h2):(1'h1)]);
                      reg212 <= reg174;
                      reg213 <= forvar181[(4'h9):(3'h6)];
                    end
                end
              else
                begin
                  if ($signed({(~^forvar170)}))
                    begin
                      reg203 <= reg154[(4'h8):(1'h0)];
                      reg204 <= $unsigned(reg178);
                      reg205 <= forvar181[(3'h7):(3'h6)];
                    end
                  else
                    begin
                      reg203 <= (!((-$signed(reg104)) ?
                          reg126[(3'h6):(2'h2)] : ((reg138 ?
                                  reg156 : forvar188) ?
                              $unsigned((8'hae)) : reg153[(3'h4):(2'h2)])));
                      reg204 <= ({(((8'ha0) <<< wire87) << (reg123 + forvar170))} ?
                          ($unsigned((reg207 ?
                              (8'hb2) : (8'ha5))) + $unsigned($unsigned((8'hb6)))) : ({(reg103 <<< forvar206)} ?
                              wire93 : $signed(reg162[(2'h2):(2'h2)])));
                    end
                end
            end
          for (forvar214 = (1'h0); (forvar214 < (2'h2)); forvar214 = (forvar214 + (1'h1)))
            begin
              if ((+(((reg114 - reg134) ^ (reg143 ? wire92 : (8'h9d))) ?
                  ($unsigned(reg100) ?
                      (~reg110) : $unsigned(reg165)) : $signed(reg148[(1'h1):(1'h1)]))))
                begin
                  if ((forvar158[(2'h2):(1'h0)] ^~ $unsigned(reg211[(4'hc):(1'h0)])))
                    begin
                      reg215 <= wire93;
                      reg216 <= reg202[(3'h6):(3'h6)];
                      reg217 <= $unsigned($signed((8'ha0)));
                      reg218 <= (~reg198[(3'h6):(2'h3)]);
                    end
                  else
                    begin
                      reg215 <= {reg213};
                      reg216 <= reg177[(2'h3):(1'h0)];
                    end
                  for (forvar219 = (1'h0); (forvar219 < (2'h3)); forvar219 = (forvar219 + (1'h1)))
                    begin
                      reg220 <= ($unsigned((wire92[(3'h4):(1'h1)] ^ $unsigned((8'ha5)))) << (~forvar170));
                      reg221 <= $unsigned(reg139);
                      reg222 <= ($unsigned($signed((forvar158 <<< reg172))) ^ (8'h9c));
                      reg223 <= (+{reg159});
                    end
                  for (forvar224 = (1'h0); (forvar224 < (1'h1)); forvar224 = (forvar224 + (1'h1)))
                    begin
                      reg225 <= ($unsigned($signed($unsigned(forvar188))) ?
                          $unsigned(reg118) : $signed($unsigned($signed((8'hab)))));
                      reg226 <= reg176[(3'h4):(2'h2)];
                      reg227 <= {reg123};
                    end
                  for (forvar228 = (1'h0); (forvar228 < (2'h3)); forvar228 = (forvar228 + (1'h1)))
                    begin
                      reg229 <= $signed({$unsigned((+reg104))});
                    end
                end
              else
                begin
                  if (reg180)
                    begin
                      reg215 <= (((reg192 ^ (&reg125)) - $unsigned(reg97)) && $signed($unsigned(reg192[(3'h6):(2'h2)])));
                      reg216 <= $unsigned($signed((wire93 && (reg167 ?
                          reg221 : reg153))));
                    end
                  else
                    begin
                      reg215 <= reg107;
                    end
                  for (forvar217 = (1'h0); (forvar217 < (1'h0)); forvar217 = (forvar217 + (1'h1)))
                    begin
                      reg218 <= reg135;
                      reg219 <= ($unsigned($unsigned({reg125})) <<< (~^reg144));
                    end
                end
              if (reg193)
                begin
                  for (forvar230 = (1'h0); (forvar230 < (1'h0)); forvar230 = (forvar230 + (1'h1)))
                    begin
                      reg231 <= $unsigned(reg159[(3'h7):(3'h7)]);
                      reg232 <= $signed($signed(reg113[(1'h1):(1'h1)]));
                      reg233 <= (~|$signed(((-reg140) << (forvar161 >>> reg101))));
                      reg234 <= (reg204[(3'h7):(1'h1)] ?
                          ((8'hba) + ((~&reg98) == {wire88})) : (-$unsigned($signed(reg183))));
                    end
                end
              else
                begin
                  for (forvar230 = (1'h0); (forvar230 < (1'h1)); forvar230 = (forvar230 + (1'h1)))
                    begin
                      reg231 <= forvar224;
                      reg232 <= ({{(8'haf)}} != ($signed((~reg187)) ?
                          {{forvar189}} : $unsigned(((8'haf) ^ reg216))));
                      reg233 <= ((8'ha0) ?
                          (!{reg139[(2'h2):(2'h2)]}) : (+((&wire90) <<< (^reg115))));
                      reg234 <= reg199;
                    end
                  for (forvar235 = (1'h0); (forvar235 < (1'h0)); forvar235 = (forvar235 + (1'h1)))
                    begin
                      reg236 <= (8'ha9);
                      reg237 <= (!$signed((~&(reg160 && forvar170))));
                    end
                  if ({(~^reg131[(1'h0):(1'h0)])})
                    begin
                      reg238 <= $signed(wire91[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg238 <= (8'h9e);
                    end
                end
              if ($unsigned((forvar188 ?
                  $signed($unsigned(reg101)) : (^(reg155 ? (8'ha9) : reg160)))))
                begin
                  if ($signed(($signed((wire88 <<< reg113)) ?
                      ((-reg186) ?
                          $unsigned(reg155) : $signed(reg196)) : ((~|reg99) ?
                          $unsigned((8'ha9)) : (reg201 * forvar181)))))
                    begin
                      reg239 <= $unsigned((|(reg116[(4'h9):(4'h9)] ?
                          $unsigned(reg127) : reg236[(3'h7):(3'h4)])));
                      reg240 <= $unsigned({reg233});
                    end
                  else
                    begin
                      reg239 <= (reg202[(4'h8):(1'h0)] + (8'ha8));
                      reg240 <= forvar210;
                      reg241 <= ({reg166} != $unsigned((!{wire92})));
                      reg242 <= forvar173;
                    end
                  if (reg182)
                    begin
                      reg243 <= reg207[(3'h7):(3'h7)];
                    end
                  else
                    begin
                      reg243 <= $signed($unsigned($unsigned((~|forvar152))));
                      reg244 <= reg209;
                    end
                end
              else
                begin
                  if (reg114)
                    begin
                      reg239 <= $unsigned(reg156[(4'hd):(2'h2)]);
                      reg240 <= reg135[(2'h2):(2'h2)];
                      reg241 <= ({(^$unsigned((8'ha3)))} && ($signed(((8'hb2) == (8'hb4))) ?
                          $signed((reg138 <= reg174)) : (^~((8'hb6) ?
                              reg197 : reg141))));
                    end
                  else
                    begin
                      reg239 <= $unsigned(($unsigned((reg129 <= (8'hb8))) ~^ (reg160[(4'h9):(4'h9)] ?
                          $signed(reg177) : $unsigned((8'ha0)))));
                      reg240 <= (|reg138[(3'h6):(1'h1)]);
                      reg241 <= (((|reg155) <= $signed((reg147 || (8'hae)))) ?
                          (reg222[(1'h0):(1'h0)] ?
                              $signed($signed(forvar181)) : {{reg242}}) : $unsigned($unsigned({forvar188})));
                    end
                  for (forvar242 = (1'h0); (forvar242 < (1'h0)); forvar242 = (forvar242 + (1'h1)))
                    begin
                      reg243 <= ($signed(reg244) || $signed({reg147}));
                    end
                  reg244 <= reg199[(4'h8):(3'h7)];
                  for (forvar245 = (1'h0); (forvar245 < (2'h2)); forvar245 = (forvar245 + (1'h1)))
                    begin
                      reg246 <= ((^{((8'had) * reg234)}) > $unsigned(reg146[(2'h2):(2'h2)]));
                    end
                end
              if (reg244[(2'h2):(1'h0)])
                begin
                  reg247 <= (reg174[(3'h6):(3'h6)] ?
                      $signed((~|(reg105 ?
                          forvar179 : reg194))) : $unsigned((^~(reg185 ?
                          reg156 : reg231))));
                  if (((^~(&(&(8'hb8)))) & $unsigned(forvar164)))
                    begin
                      reg248 <= (~&$signed((8'hb6)));
                      reg249 <= (+(&({reg110} > (reg97 ? reg177 : reg220))));
                      reg250 <= (reg136[(4'ha):(3'h7)] ?
                          forvar161 : (-$signed(((8'hb0) ?
                              (8'h9f) : forvar235))));
                    end
                  else
                    begin
                      reg248 <= reg215;
                      reg249 <= (((8'ha8) ?
                          $unsigned(((8'h9d) || (8'h9c))) : (~$unsigned(forvar224))) >= (|reg121));
                      reg250 <= $signed($unsigned(((&(8'ha6)) <= reg139[(3'h7):(3'h5)])));
                      reg251 <= $signed(($signed(reg177[(4'h8):(3'h5)]) ?
                          reg154[(4'h8):(1'h1)] : forvar149[(1'h0):(1'h0)]));
                    end
                  if ($unsigned(reg251[(2'h2):(1'h0)]))
                    begin
                      reg252 <= reg168;
                      reg253 <= $signed(reg169[(4'h8):(1'h0)]);
                      reg254 <= (~|$unsigned(({reg136} ~^ reg155[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg252 <= $signed($signed($signed($unsigned((8'ha4)))));
                      reg253 <= ({reg229[(2'h3):(2'h3)]} < forvar181[(3'h4):(2'h3)]);
                      reg254 <= (~|(8'haf));
                      reg255 <= (+reg194[(1'h1):(1'h1)]);
                    end
                  if (forvar190[(4'hb):(3'h6)])
                    begin
                      reg256 <= ((reg145[(1'h0):(1'h0)] ?
                          $unsigned((~^reg101)) : $signed((reg134 >= reg169))) * $signed((+$unsigned(reg199))));
                    end
                  else
                    begin
                      reg256 <= (~|((reg180[(3'h5):(3'h5)] >= $signed(reg208)) <<< $unsigned($signed(reg183))));
                    end
                end
              else
                begin
                  reg247 <= $unsigned($signed(reg146[(4'hc):(4'h9)]));
                  reg248 <= reg109;
                end
            end
          for (forvar257 = (1'h0); (forvar257 < (1'h0)); forvar257 = (forvar257 + (1'h1)))
            begin
              reg258 <= reg105;
              for (forvar259 = (1'h0); (forvar259 < (1'h0)); forvar259 = (forvar259 + (1'h1)))
                begin
                  if (reg155)
                    begin
                      reg260 <= {forvar210};
                      reg261 <= $unsigned($unsigned((~&{reg125})));
                      reg262 <= reg261[(2'h3):(2'h2)];
                      reg263 <= (reg198[(3'h6):(3'h4)] ?
                          (|reg162[(1'h1):(1'h0)]) : $signed((~reg171[(4'h9):(3'h6)])));
                    end
                  else
                    begin
                      reg260 <= ($unsigned((reg99 < (!reg212))) | forvar245);
                    end
                  if (reg185)
                    begin
                      reg264 <= forvar228;
                    end
                  else
                    begin
                      reg264 <= ($signed((~&reg221[(4'h9):(1'h0)])) || {((8'hae) ?
                              $signed(reg240) : reg142)});
                    end
                end
              for (forvar265 = (1'h0); (forvar265 < (1'h1)); forvar265 = (forvar265 + (1'h1)))
                begin
                  for (forvar266 = (1'h0); (forvar266 < (1'h1)); forvar266 = (forvar266 + (1'h1)))
                    begin
                      reg267 <= (+(+(8'hac)));
                      reg268 <= reg171[(3'h6):(2'h3)];
                      reg269 <= reg237[(1'h1):(1'h1)];
                      reg270 <= ($signed(forvar152) ?
                          ({reg217} != $signed($unsigned(reg212))) : ((!(reg191 ?
                                  (8'ha2) : reg128)) ?
                              (8'hb6) : {((8'hb5) || (8'hb5))}));
                    end
                end
            end
        end
      if ($signed((($signed((8'ha1)) ? $signed(forvar214) : reg178) ?
          reg182[(4'hb):(1'h1)] : $signed(forvar228))))
        begin
          if ((reg226[(3'h6):(3'h6)] ?
              ((-(~(8'ha5))) - {(&reg269)}) : ((+forvar257[(3'h4):(1'h1)]) ?
                  $unsigned((8'hb6)) : ((8'hb2) >= $unsigned(reg131)))))
            begin
              if ((^~((((8'ha3) ? reg156 : reg110) ?
                  $signed(reg135) : (reg270 ? (8'h9e) : forvar164)) >= reg253)))
                begin
                  reg271 <= reg250[(3'h7):(1'h0)];
                  for (forvar272 = (1'h0); (forvar272 < (1'h0)); forvar272 = (forvar272 + (1'h1)))
                    begin
                      reg273 <= $signed(($signed($signed(reg144)) ?
                          reg191 : forvar228[(2'h3):(1'h1)]));
                    end
                  for (forvar274 = (1'h0); (forvar274 < (2'h3)); forvar274 = (forvar274 + (1'h1)))
                    begin
                      reg275 <= $signed($signed(((reg109 ?
                          reg126 : reg226) >>> $signed(reg123))));
                      reg276 <= reg263;
                      reg277 <= reg107[(3'h7):(3'h5)];
                    end
                  for (forvar278 = (1'h0); (forvar278 < (1'h0)); forvar278 = (forvar278 + (1'h1)))
                    begin
                      reg279 <= reg139[(4'hc):(3'h7)];
                      reg280 <= (+($unsigned((reg168 ? reg240 : forvar163)) ?
                          ($unsigned(reg246) && (reg269 | reg128)) : (~^reg222[(1'h0):(1'h0)])));
                      reg281 <= (8'hb2);
                      reg282 <= ({(^~reg98[(4'h8):(1'h0)])} ?
                          $signed($signed(((8'ha2) * reg280))) : $signed((|(wire91 ?
                              reg144 : reg231))));
                    end
                end
              else
                begin
                  for (forvar271 = (1'h0); (forvar271 < (1'h0)); forvar271 = (forvar271 + (1'h1)))
                    begin
                      reg272 <= reg223;
                      reg273 <= $unsigned((($signed((8'ha2)) & $signed(reg110)) ?
                          {reg242} : ((reg234 ? reg199 : forvar257) ?
                              $unsigned(forvar150) : $unsigned(reg111))));
                      reg274 <= $signed(reg209[(3'h5):(3'h4)]);
                      reg275 <= reg194[(2'h2):(2'h2)];
                    end
                  for (forvar276 = (1'h0); (forvar276 < (2'h3)); forvar276 = (forvar276 + (1'h1)))
                    begin
                      reg277 <= ((((8'hb1) && $unsigned(reg213)) <<< $signed((reg216 || reg264))) ?
                          $unsigned((8'ha2)) : $unsigned((forvar151[(1'h0):(1'h0)] - reg231[(3'h6):(3'h6)])));
                      reg278 <= reg115[(2'h2):(2'h2)];
                    end
                end
              for (forvar283 = (1'h0); (forvar283 < (1'h1)); forvar283 = (forvar283 + (1'h1)))
                begin
                  for (forvar284 = (1'h0); (forvar284 < (1'h0)); forvar284 = (forvar284 + (1'h1)))
                    begin
                      reg285 <= $signed(reg121);
                      reg286 <= ((&(|forvar242)) ?
                          $unsigned({reg129}) : $unsigned(((reg156 - reg123) > reg281)));
                    end
                  for (forvar287 = (1'h0); (forvar287 < (2'h3)); forvar287 = (forvar287 + (1'h1)))
                    begin
                      reg288 <= {$unsigned(forvar158[(2'h3):(2'h2)])};
                      reg289 <= ((({(8'hb9)} >= (reg169 ~^ reg180)) < (reg261[(4'hb):(3'h7)] != $unsigned(reg103))) ?
                          $unsigned(($unsigned((8'ha1)) | (reg260 | (8'ha2)))) : $signed(((reg134 ?
                              reg241 : (8'ha1)) < $signed(forvar150))));
                      reg290 <= (+(($signed(reg285) < {reg286}) ?
                          ({reg241} ?
                              {wire93} : reg121) : ((reg268 * forvar276) ?
                              reg212 : (reg180 ? reg280 : reg226))));
                      reg291 <= ($signed(reg229[(3'h5):(3'h4)]) && reg177);
                    end
                  for (forvar292 = (1'h0); (forvar292 < (2'h2)); forvar292 = (forvar292 + (1'h1)))
                    begin
                      reg293 <= (^(forvar272 >> reg128[(3'h5):(1'h1)]));
                      reg294 <= {$signed({(reg278 ? (8'ha9) : forvar274)})};
                      reg295 <= (forvar271[(4'h9):(2'h3)] | {reg219[(1'h1):(1'h1)]});
                      reg296 <= (((~|$signed(reg169)) ?
                              $unsigned(reg154[(2'h3):(2'h3)]) : $signed($unsigned(reg229))) ?
                          (~&((~&(8'hb6)) - $unsigned(reg101))) : (forvar190 ?
                              wire93 : (reg277 ?
                                  (+wire91) : ((8'haa) >>> reg272))));
                    end
                end
              for (forvar297 = (1'h0); (forvar297 < (2'h2)); forvar297 = (forvar297 + (1'h1)))
                begin
                  for (forvar298 = (1'h0); (forvar298 < (1'h1)); forvar298 = (forvar298 + (1'h1)))
                    begin
                      reg299 <= forvar181;
                      reg300 <= (~&($signed((~|wire88)) <<< $signed((&(8'hb1)))));
                    end
                  if (reg253)
                    begin
                      reg301 <= (!$unsigned((forvar150[(3'h7):(1'h1)] ^~ (reg281 ?
                          (8'ha1) : (8'haa)))));
                    end
                  else
                    begin
                      reg301 <= (8'h9f);
                      reg302 <= ($unsigned({reg208[(2'h3):(1'h1)]}) >> {((reg141 ~^ reg194) != reg237)});
                      reg303 <= reg109;
                    end
                end
            end
          else
            begin
              for (forvar271 = (1'h0); (forvar271 < (2'h2)); forvar271 = (forvar271 + (1'h1)))
                begin
                  for (forvar272 = (1'h0); (forvar272 < (1'h1)); forvar272 = (forvar272 + (1'h1)))
                    begin
                      reg273 <= ((!reg275[(4'he):(3'h5)]) <= (reg232[(4'hb):(4'ha)] ?
                          $unsigned(reg213) : ($signed(reg148) <<< reg300)));
                      reg274 <= (+$signed((~|$signed(reg193))));
                      reg275 <= reg169;
                    end
                  if (($unsigned($signed(wire93[(1'h0):(1'h0)])) >>> $signed((-(forvar161 & (8'ha7))))))
                    begin
                      reg276 <= (($unsigned((forvar219 ?
                          forvar161 : reg199)) ^~ reg121[(1'h1):(1'h1)]) > $signed(($signed(reg264) ^ (~&reg277))));
                    end
                  else
                    begin
                      reg276 <= (&($signed(reg155) != ($signed(reg140) >= $signed(reg212))));
                      reg277 <= $unsigned((~^$signed((reg301 ?
                          wire92 : reg126))));
                      reg278 <= reg117[(3'h4):(1'h1)];
                      reg279 <= $unsigned(($signed((~|forvar161)) <<< reg251[(3'h6):(2'h3)]));
                    end
                  reg280 <= wire87[(4'h8):(3'h7)];
                  for (forvar281 = (1'h0); (forvar281 < (1'h1)); forvar281 = (forvar281 + (1'h1)))
                    begin
                      reg282 <= (forvar257[(4'hb):(2'h2)] << (^{$unsigned(reg227)}));
                      reg283 <= ($signed((~(reg276 >> reg243))) ?
                          $signed($signed($signed(reg222))) : ($unsigned((forvar150 >= reg98)) != reg103));
                      reg284 <= (^{$signed({reg129})});
                    end
                end
              for (forvar285 = (1'h0); (forvar285 < (1'h1)); forvar285 = (forvar285 + (1'h1)))
                begin
                  if ($signed((reg284 >= reg105)))
                    begin
                      reg286 <= (&(8'hb4));
                      reg287 <= {(^~$signed({reg195}))};
                      reg288 <= (forvar266[(3'h5):(1'h1)] && reg268[(3'h5):(2'h2)]);
                    end
                  else
                    begin
                      reg286 <= $signed({((reg117 * reg107) ?
                              $unsigned(reg134) : reg157[(3'h5):(2'h2)])});
                      reg287 <= $signed(((((8'ha3) ?
                              reg216 : reg101) >>> (wire90 ?
                              (8'ha8) : reg287)) ?
                          $signed(forvar224) : $signed((+reg249))));
                      reg288 <= ((reg100 ?
                              $signed((reg258 & (8'haa))) : (~$signed(reg195))) ?
                          (+(^~reg241)) : $unsigned(reg272));
                    end
                  reg289 <= (($unsigned(reg107[(3'h7):(3'h7)]) == ($signed((8'ha9)) ?
                          (forvar181 && (8'hba)) : reg209[(2'h2):(1'h1)])) ?
                      (+(+{reg246})) : $signed($unsigned((forvar181 ?
                          forvar292 : wire89))));
                  if (($unsigned(reg269[(3'h7):(3'h4)]) ?
                      $unsigned({((8'ha6) ?
                              reg208 : reg256)}) : ($unsigned(((8'ha2) * reg246)) ?
                          (8'hb0) : wire90[(3'h7):(1'h0)])))
                    begin
                      reg290 <= $unsigned(reg187);
                      reg291 <= (wire92 ^~ (reg123[(4'h9):(1'h0)] ?
                          (^~(^~reg240)) : ($unsigned(forvar161) && $signed(reg115))));
                      reg292 <= reg238;
                    end
                  else
                    begin
                      reg290 <= forvar274[(2'h2):(1'h0)];
                      reg291 <= forvar149;
                    end
                  for (forvar293 = (1'h0); (forvar293 < (2'h2)); forvar293 = (forvar293 + (1'h1)))
                    begin
                      reg294 <= reg121[(4'hb):(4'h9)];
                    end
                end
            end
          reg304 <= {(((reg184 ^~ reg272) <<< ((8'haa) - reg212)) && $signed($signed(forvar188)))};
          for (forvar305 = (1'h0); (forvar305 < (2'h3)); forvar305 = (forvar305 + (1'h1)))
            begin
              for (forvar306 = (1'h0); (forvar306 < (2'h3)); forvar306 = (forvar306 + (1'h1)))
                begin
                  for (forvar307 = (1'h0); (forvar307 < (2'h3)); forvar307 = (forvar307 + (1'h1)))
                    begin
                      reg308 <= (($unsigned((~|reg215)) & ($unsigned(reg174) ^~ $unsigned(reg283))) ?
                          $unsigned(reg103[(4'hc):(1'h0)]) : (^~((forvar278 + reg121) * (~|wire89))));
                    end
                  for (forvar309 = (1'h0); (forvar309 < (1'h0)); forvar309 = (forvar309 + (1'h1)))
                    begin
                      reg310 <= ((8'hb7) ^ (&{$unsigned(reg197)}));
                      reg311 <= reg201[(3'h6):(3'h5)];
                    end
                  for (forvar312 = (1'h0); (forvar312 < (2'h3)); forvar312 = (forvar312 + (1'h1)))
                    begin
                      reg313 <= forvar235;
                    end
                  if ((-$signed(forvar163[(2'h3):(2'h3)])))
                    begin
                      reg314 <= {reg200[(2'h2):(1'h0)]};
                      reg315 <= (($unsigned($signed(reg276)) ?
                          ((reg239 >> reg128) >> reg231) : $unsigned($signed(reg199))) >>> $unsigned(($signed(reg278) >>> (wire87 ?
                          forvar271 : reg211))));
                      reg316 <= (~$unsigned($signed($signed(reg110))));
                      reg317 <= ($signed($unsigned((reg142 ?
                          reg223 : reg255))) | ((~|(reg143 >> forvar306)) < (forvar163[(1'h0):(1'h0)] | reg251[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg314 <= reg100;
                      reg315 <= reg129[(1'h1):(1'h1)];
                      reg316 <= (((&$signed(reg271)) ^ $unsigned((reg121 && (8'hb7)))) >= $unsigned((8'ha3)));
                      reg317 <= forvar228[(1'h0):(1'h0)];
                    end
                end
              if ((|(forvar214[(3'h4):(1'h0)] ?
                  $unsigned(((8'haf) ?
                      (8'hb9) : forvar217)) : {(reg315 >= reg186)})))
                begin
                  for (forvar318 = (1'h0); (forvar318 < (1'h0)); forvar318 = (forvar318 + (1'h1)))
                    begin
                      reg319 <= $signed((8'ha8));
                    end
                end
              else
                begin
                  if (reg269[(3'h4):(2'h2)])
                    begin
                      reg318 <= (($unsigned((wire87 ?
                              reg293 : (8'h9e))) && ($signed(reg242) ?
                              forvar210[(4'ha):(3'h5)] : {reg236})) ?
                          $signed(wire89[(1'h0):(1'h0)]) : (^((reg111 - reg142) ?
                              reg104 : forvar164[(3'h5):(3'h4)])));
                      reg319 <= forvar285[(1'h0):(1'h0)];
                      reg320 <= reg166;
                      reg321 <= ((~$unsigned((reg276 ? reg271 : reg261))) ?
                          reg142 : $unsigned((-$signed((8'ha9)))));
                    end
                  else
                    begin
                      reg318 <= reg283;
                    end
                  if ($unsigned(reg153))
                    begin
                      reg322 <= (reg213[(3'h4):(2'h3)] ?
                          $signed(reg143[(3'h5):(3'h5)]) : ((reg191[(1'h1):(1'h1)] >> (reg191 | reg100)) <= (~&$unsigned(reg153))));
                    end
                  else
                    begin
                      reg322 <= ((($unsigned(forvar265) >>> $unsigned(reg146)) ^ (!reg128[(1'h1):(1'h0)])) ?
                          ((reg237 ?
                              ((8'h9f) > forvar228) : {reg213}) * ((reg254 ?
                                  reg135 : forvar271) ?
                              (reg315 + reg290) : (~|reg169))) : ($signed(((8'hae) ?
                                  reg196 : reg166)) ?
                              (reg291[(1'h1):(1'h0)] ?
                                  {reg251} : $signed(reg186)) : $unsigned($signed(forvar228))));
                      reg323 <= reg254;
                      reg324 <= (forvar306 ? reg272 : reg284);
                    end
                end
              for (forvar325 = (1'h0); (forvar325 < (2'h3)); forvar325 = (forvar325 + (1'h1)))
                begin
                  for (forvar326 = (1'h0); (forvar326 < (2'h3)); forvar326 = (forvar326 + (1'h1)))
                    begin
                      reg327 <= $signed($unsigned((^~$unsigned(reg98))));
                      reg328 <= $signed(reg278[(4'h9):(2'h3)]);
                      reg329 <= $unsigned($unsigned((^(reg220 >= wire89))));
                      reg330 <= $signed({$unsigned({reg121})});
                    end
                  if ((~^(reg209[(4'hb):(4'h9)] ?
                      ($signed((8'hb8)) >> (|reg143)) : (-((8'ha3) ?
                          reg299 : reg277)))))
                    begin
                      reg331 <= reg268;
                      reg332 <= (^$signed(($signed(reg217) ^~ ((8'haf) && reg122))));
                    end
                  else
                    begin
                      reg331 <= $unsigned(reg308[(3'h6):(1'h1)]);
                      reg332 <= $signed(($unsigned($signed((8'hb2))) ?
                          reg258[(1'h0):(1'h0)] : $signed((reg311 && wire89))));
                      reg333 <= ((^((reg128 && reg231) >>> $signed(forvar278))) == (|(8'hab)));
                      reg334 <= $unsigned(({$signed(reg101)} ?
                          {$signed(reg153)} : reg302));
                    end
                  for (forvar335 = (1'h0); (forvar335 < (1'h1)); forvar335 = (forvar335 + (1'h1)))
                    begin
                      reg336 <= $signed(reg113[(1'h0):(1'h0)]);
                      reg337 <= (~&{reg321});
                      reg338 <= (($signed(forvar170[(2'h2):(1'h1)]) != reg268) ?
                          ({$unsigned((8'ha8))} <<< reg139[(3'h5):(2'h2)]) : $signed(reg105[(2'h3):(1'h0)]));
                    end
                  reg339 <= ((({reg97} + $signed(forvar293)) ?
                      ((^reg322) > (reg204 & forvar307)) : {$unsigned(wire88)}) && $signed(($unsigned(reg271) ~^ reg243)));
                end
            end
        end
      else
        begin
          for (forvar271 = (1'h0); (forvar271 < (2'h2)); forvar271 = (forvar271 + (1'h1)))
            begin
              if (((&reg295) ~^ ((~&(~^reg287)) >> $unsigned((&forvar214)))))
                begin
                  if ((+$unsigned(reg135[(1'h1):(1'h1)])))
                    begin
                      reg272 <= (~&$signed($unsigned($signed((8'h9d)))));
                      reg273 <= {$signed({reg104})};
                      reg274 <= $unsigned($unsigned({reg329[(1'h1):(1'h1)]}));
                      reg275 <= reg282[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg272 <= ({forvar163[(1'h1):(1'h0)]} ?
                          forvar150[(4'hb):(3'h5)] : $unsigned((reg229 ?
                              ((8'hb9) ?
                                  forvar297 : reg103) : $unsigned(forvar257))));
                      reg273 <= (!$unsigned(reg295[(3'h5):(2'h2)]));
                      reg274 <= $signed($unsigned(((~^reg308) < $signed(forvar292))));
                    end
                  for (forvar276 = (1'h0); (forvar276 < (2'h2)); forvar276 = (forvar276 + (1'h1)))
                    begin
                      reg277 <= (~|((reg157 ?
                          $unsigned(reg202) : reg184[(4'hc):(4'hc)]) ~^ $signed(reg264[(3'h5):(3'h4)])));
                    end
                end
              else
                begin
                  for (forvar272 = (1'h0); (forvar272 < (1'h1)); forvar272 = (forvar272 + (1'h1)))
                    begin
                      reg273 <= (($unsigned((forvar219 ? reg289 : (8'hb5))) ?
                          (-(8'ha7)) : {(reg223 - reg264)}) << (!(&reg276[(1'h1):(1'h1)])));
                      reg274 <= {($unsigned(forvar206) ?
                              (~&(reg192 ?
                                  forvar158 : reg146)) : $unsigned(forvar206))};
                      reg275 <= ($unsigned((((8'hb6) << reg244) ?
                              (forvar287 ?
                                  forvar217 : (8'haa)) : (reg319 <<< forvar285))) ?
                          $unsigned($unsigned($unsigned(reg146))) : ($unsigned(reg160) ~^ (!$signed(forvar164))));
                    end
                end
              if ((^~($unsigned(reg239) ?
                  reg185 : $unsigned($unsigned(forvar305)))))
                begin
                  if ($signed((((reg331 ? reg219 : reg314) ?
                      (reg112 ? reg117 : reg209) : forvar272) + reg112)))
                    begin
                      reg278 <= forvar325[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg278 <= ($signed(((reg278 ?
                          reg248 : reg248) | $unsigned(reg98))) >> ({(reg135 == (8'hb9))} < reg246[(1'h1):(1'h0)]));
                      reg279 <= reg313;
                    end
                end
              else
                begin
                  for (forvar278 = (1'h0); (forvar278 < (2'h2)); forvar278 = (forvar278 + (1'h1)))
                    begin
                      reg279 <= {reg327};
                      reg280 <= {(&(((8'hac) ? reg157 : (8'hb2)) ?
                              reg165 : (reg178 ? reg284 : forvar281)))};
                    end
                  for (forvar281 = (1'h0); (forvar281 < (1'h1)); forvar281 = (forvar281 + (1'h1)))
                    begin
                      reg282 <= $signed($signed((((8'ha7) ^~ reg321) ?
                          (8'ha2) : $signed(reg256))));
                      reg283 <= $signed((8'ha0));
                    end
                  for (forvar284 = (1'h0); (forvar284 < (2'h3)); forvar284 = (forvar284 + (1'h1)))
                    begin
                      reg285 <= $signed($signed($unsigned((^(8'h9e)))));
                      reg286 <= reg178;
                      reg287 <= $signed($signed($signed((reg146 >>> (8'ha7)))));
                      reg288 <= (&(reg303 ? (~^(^reg329)) : (~|reg241)));
                    end
                end
              if (reg231)
                begin
                  if ((~^((^~reg213) <<< (^reg191))))
                    begin
                      reg289 <= wire89;
                      reg290 <= $unsigned(reg154[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg289 <= $signed((!$signed(reg338)));
                      reg290 <= ($unsigned($unsigned($unsigned((8'ha0)))) <<< ($unsigned((reg100 ?
                          reg225 : reg268)) <<< $signed($unsigned(reg191))));
                    end
                end
              else
                begin
                  for (forvar289 = (1'h0); (forvar289 < (1'h1)); forvar289 = (forvar289 + (1'h1)))
                    begin
                      reg290 <= {(^~(|(~(8'hb9))))};
                      reg291 <= (((|(~forvar189)) ?
                              (-forvar283[(3'h4):(2'h3)]) : {(~^reg301)}) ?
                          ((reg171 ?
                              forvar312[(2'h2):(1'h0)] : reg247[(2'h2):(1'h1)]) <= (~^$unsigned((8'h9c)))) : $signed(((reg116 != reg247) ?
                              {reg202} : reg254)));
                    end
                  if ((({((8'ha3) ?
                              reg131 : reg218)} & $signed($unsigned((8'hb5)))) ?
                      reg208 : reg322[(1'h1):(1'h0)]))
                    begin
                      reg292 <= ((+(~{reg182})) ?
                          wire93[(3'h4):(1'h0)] : forvar242);
                      reg293 <= (-(!reg140[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg292 <= $signed(reg331);
                      reg293 <= (reg115 <<< (forvar214 ?
                          ((~^forvar170) ?
                              reg242 : $signed(reg339)) : $signed({reg232})));
                      reg294 <= (($unsigned(reg222) ?
                              $unsigned(reg177[(3'h5):(2'h3)]) : reg112) ?
                          forvar259 : forvar309[(4'he):(3'h6)]);
                      reg295 <= (~|$unsigned(reg251));
                    end
                end
            end
        end
      if ($unsigned(((~reg223[(3'h6):(2'h2)]) - ((forvar210 * forvar235) - (+wire88)))))
        begin
          for (forvar340 = (1'h0); (forvar340 < (2'h2)); forvar340 = (forvar340 + (1'h1)))
            begin
              if (forvar190)
                begin
                  if ($signed((reg198 ^ reg289[(2'h2):(2'h2)])))
                    begin
                      reg341 <= (forvar318[(1'h1):(1'h1)] ?
                          wire91[(3'h5):(1'h1)] : ({$signed(reg315)} >= (~(~&reg127))));
                      reg342 <= (reg270[(3'h4):(1'h0)] != reg195);
                      reg343 <= {$unsigned({reg166})};
                      reg344 <= (^(+((reg300 && (8'hb5)) | (~|reg177))));
                    end
                  else
                    begin
                      reg341 <= forvar266;
                      reg342 <= reg276[(2'h2):(2'h2)];
                      reg343 <= $signed((8'haf));
                      reg344 <= $signed({$signed((-forvar266))});
                    end
                  for (forvar345 = (1'h0); (forvar345 < (2'h2)); forvar345 = (forvar345 + (1'h1)))
                    begin
                      reg346 <= reg104;
                      reg347 <= $signed(forvar287);
                    end
                end
              else
                begin
                  if (reg252[(1'h0):(1'h0)])
                    begin
                      reg341 <= reg219;
                      reg342 <= $signed(forvar149);
                      reg343 <= ($unsigned(forvar266[(4'ha):(3'h6)]) ?
                          ((((8'hae) <= reg215) ?
                              reg227 : (reg169 | forvar285)) | reg203[(4'he):(4'h9)]) : {($unsigned(reg199) >>> (reg168 ?
                                  reg105 : reg221))});
                    end
                  else
                    begin
                      reg341 <= $unsigned($signed((8'hb1)));
                      reg342 <= reg220;
                    end
                  if ($unsigned($unsigned(reg186)))
                    begin
                      reg344 <= reg269[(2'h3):(2'h3)];
                      reg345 <= $signed(reg315);
                      reg346 <= reg171[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg344 <= $unsigned((^{(!reg321)}));
                      reg345 <= reg200[(2'h3):(1'h1)];
                      reg346 <= (reg241[(3'h5):(3'h5)] ?
                          reg273[(2'h2):(1'h0)] : reg308[(1'h0):(1'h0)]);
                      reg347 <= reg105[(1'h0):(1'h0)];
                    end
                  if ($unsigned(((reg128 ?
                          (reg155 < reg271) : reg168[(2'h2):(2'h2)]) ?
                      $unsigned($unsigned(reg205)) : $signed(reg345))))
                    begin
                      reg348 <= $unsigned($unsigned((+(8'hb4))));
                      reg349 <= ((forvar219[(1'h0):(1'h0)] < ($unsigned(reg271) ?
                              (^~reg323) : (~|reg242))) ?
                          forvar309[(3'h7):(1'h0)] : reg346);
                    end
                  else
                    begin
                      reg348 <= ($unsigned($signed((forvar228 < forvar173))) ?
                          reg103 : (($unsigned(forvar266) ?
                              (8'ha9) : $signed(reg204)) >= $signed(reg208)));
                      reg349 <= (((~$unsigned(forvar164)) ?
                              reg226[(2'h3):(2'h2)] : (+reg248)) ?
                          $unsigned($unsigned(((8'ha1) ?
                              reg191 : reg100))) : ($unsigned(reg285) ?
                              $signed((|reg118)) : $unsigned($signed(reg114))));
                      reg350 <= $signed(({$signed(forvar289)} ~^ {$signed((8'ha4))}));
                    end
                end
              for (forvar351 = (1'h0); (forvar351 < (2'h2)); forvar351 = (forvar351 + (1'h1)))
                begin
                  for (forvar352 = (1'h0); (forvar352 < (1'h0)); forvar352 = (forvar352 + (1'h1)))
                    begin
                      reg353 <= $unsigned($signed(((reg196 ?
                          reg101 : (8'hb4)) >= $unsigned(forvar274))));
                      reg354 <= (~&{(8'h9d)});
                      reg355 <= (($signed({reg320}) ?
                              $unsigned(reg260[(1'h1):(1'h1)]) : reg354[(3'h4):(2'h3)]) ?
                          ((^~((8'ha6) ? forvar340 : reg169)) ?
                              (^reg282[(3'h4):(2'h2)]) : ($unsigned(reg342) ^~ $unsigned(reg159))) : reg264);
                    end
                  for (forvar356 = (1'h0); (forvar356 < (1'h1)); forvar356 = (forvar356 + (1'h1)))
                    begin
                      reg357 <= $signed((|reg165[(1'h1):(1'h0)]));
                    end
                  for (forvar358 = (1'h0); (forvar358 < (1'h0)); forvar358 = (forvar358 + (1'h1)))
                    begin
                      reg359 <= (|$unsigned($signed((|reg165))));
                      reg360 <= (8'ha7);
                      reg361 <= ((-((~^reg191) < reg320[(1'h0):(1'h0)])) ?
                          ($signed(forvar259[(2'h3):(2'h2)]) & $signed(reg176[(1'h1):(1'h1)])) : {{(reg125 + reg98)}});
                    end
                end
              for (forvar362 = (1'h0); (forvar362 < (2'h2)); forvar362 = (forvar362 + (1'h1)))
                begin
                  for (forvar363 = (1'h0); (forvar363 < (1'h1)); forvar363 = (forvar363 + (1'h1)))
                    begin
                      reg364 <= reg278;
                      reg365 <= reg244;
                    end
                  if ($signed($unsigned(($unsigned(reg293) <= (reg247 ?
                      reg247 : reg128)))))
                    begin
                      reg366 <= (!({{reg127}} ~^ (8'ha0)));
                    end
                  else
                    begin
                      reg366 <= $signed($unsigned($unsigned((reg263 - reg213))));
                      reg367 <= (($unsigned(reg168) ? (8'hb1) : reg219) ?
                          ($signed($signed((8'had))) < {(reg314 >> reg311)}) : ({forvar326[(3'h4):(2'h2)]} > $signed((reg194 ?
                              (8'h9e) : forvar181))));
                      reg368 <= reg131[(1'h0):(1'h0)];
                      reg369 <= ($unsigned(reg274[(2'h2):(2'h2)]) ?
                          forvar271 : reg323);
                    end
                end
              reg370 <= $signed((({reg349} ?
                      forvar312 : reg212[(1'h0):(1'h0)]) ?
                  reg327[(3'h6):(3'h4)] : (reg159 * reg128)));
            end
          reg371 <= reg110[(4'h9):(1'h1)];
        end
      else
        begin
          for (forvar340 = (1'h0); (forvar340 < (1'h0)); forvar340 = (forvar340 + (1'h1)))
            begin
              if ($unsigned(((reg139[(1'h1):(1'h0)] + ((8'h9e) ?
                      reg268 : reg223)) ?
                  $signed(reg111) : reg243)))
                begin
                  for (forvar341 = (1'h0); (forvar341 < (1'h1)); forvar341 = (forvar341 + (1'h1)))
                    begin
                      reg342 <= $unsigned($unsigned((8'hb4)));
                      reg343 <= $unsigned(wire89);
                    end
                end
              else
                begin
                  reg341 <= $signed(((reg115 ~^ (reg99 ?
                      forvar235 : forvar326)) || reg286[(2'h2):(2'h2)]));
                end
              if ((($signed((~&forvar352)) ^ reg314) ?
                  $signed(reg361[(4'hc):(4'h9)]) : ({$signed(reg292)} && (8'ha8))))
                begin
                  if ((reg353[(2'h3):(1'h0)] ~^ ($unsigned((reg201 != reg284)) ?
                      (^~(reg225 == forvar363)) : (~reg274[(2'h2):(1'h0)]))))
                    begin
                      reg344 <= $unsigned($unsigned(({reg162} < (forvar341 ?
                          (8'hb5) : forvar325))));
                    end
                  else
                    begin
                      reg344 <= $signed((!reg283[(1'h0):(1'h0)]));
                      reg345 <= $signed(((((8'hb2) >> forvar230) ?
                          (reg279 ?
                              reg101 : reg110) : reg248) > ((reg262 * forvar158) - (reg112 ?
                          reg302 : reg357))));
                    end
                  if (reg281)
                    begin
                      reg346 <= $unsigned((~|($unsigned(reg209) & $unsigned(reg234))));
                      reg347 <= (~|(reg124[(3'h4):(2'h2)] != $signed((forvar272 >> reg271))));
                      reg348 <= $unsigned($unsigned($unsigned((8'ha4))));
                      reg349 <= $signed($signed((reg124[(3'h5):(2'h3)] ?
                          $signed((8'hb2)) : {forvar265})));
                    end
                  else
                    begin
                      reg346 <= {($unsigned((~(8'h9d))) & {(reg334 && reg128)})};
                      reg347 <= reg329[(2'h2):(1'h0)];
                      reg348 <= forvar297;
                      reg349 <= (8'ha0);
                    end
                end
              else
                begin
                  for (forvar344 = (1'h0); (forvar344 < (2'h3)); forvar344 = (forvar344 + (1'h1)))
                    begin
                      reg345 <= $unsigned($unsigned($signed(((8'hb8) << forvar150))));
                      reg346 <= ((reg341 ?
                          (~^$unsigned(reg234)) : (~&$signed((8'haa)))) * $signed(reg145[(2'h3):(1'h1)]));
                      reg347 <= {$signed($signed(reg216[(3'h7):(2'h2)]))};
                    end
                  reg348 <= reg338;
                end
              for (forvar350 = (1'h0); (forvar350 < (2'h3)); forvar350 = (forvar350 + (1'h1)))
                begin
                  reg351 <= reg300[(4'hb):(4'h8)];
                  for (forvar352 = (1'h0); (forvar352 < (2'h3)); forvar352 = (forvar352 + (1'h1)))
                    begin
                      reg353 <= {(~^reg201[(4'h9):(1'h0)])};
                      reg354 <= reg191[(3'h5):(3'h4)];
                      reg355 <= (forvar149[(3'h5):(3'h5)] != ((^~(forvar190 & reg280)) ?
                          reg168 : (^~(~|(8'ha9)))));
                      reg356 <= (~&(8'h9d));
                    end
                  if (((reg348[(1'h1):(1'h1)] > (8'h9d)) == wire89))
                    begin
                      reg357 <= (((8'ha5) <<< reg318[(2'h2):(1'h0)]) ?
                          reg282[(2'h2):(2'h2)] : reg136);
                      reg358 <= (((|$signed(forvar257)) <= ($unsigned(reg252) ?
                              {reg371} : (+reg115))) ?
                          $unsigned((|{(8'ha3)})) : $signed($signed($signed(reg234))));
                      reg359 <= ($unsigned({(reg129 << (8'ha3))}) <= reg333);
                    end
                  else
                    begin
                      reg357 <= $unsigned({(~&$unsigned(forvar271))});
                      reg358 <= $unsigned((8'h9e));
                    end
                  if (reg337)
                    begin
                      reg360 <= (-(reg165 ?
                          (reg177 ?
                              (|wire90) : reg324[(2'h3):(1'h1)]) : (reg147 ?
                              (8'ha8) : (forvar335 >= forvar217))));
                      reg361 <= $unsigned($signed($signed({reg215})));
                      reg362 <= ($unsigned($signed((reg177 ?
                              reg136 : reg308))) ?
                          $signed((reg226 ? (8'hba) : {reg184})) : ((((8'ha5) ?
                                      forvar358 : reg262) ?
                                  (~|reg268) : reg358) ?
                              (^~reg215) : $signed($signed(forvar335))));
                    end
                  else
                    begin
                      reg360 <= reg113[(1'h0):(1'h0)];
                      reg361 <= $unsigned(forvar318[(1'h0):(1'h0)]);
                      reg362 <= reg319[(3'h4):(1'h0)];
                      reg363 <= (~(~|$unsigned($unsigned(forvar189))));
                    end
                end
              for (forvar364 = (1'h0); (forvar364 < (2'h2)); forvar364 = (forvar364 + (1'h1)))
                begin
                  reg365 <= (!($signed((reg295 <= reg252)) ?
                      ($signed(reg331) <= {forvar189}) : (reg191 > (reg129 ?
                          forvar283 : reg339))));
                  if (($unsigned($unsigned(reg118)) ?
                      (8'hac) : ((8'ha8) + $signed(reg250[(1'h1):(1'h0)]))))
                    begin
                      reg366 <= reg126[(4'h8):(3'h5)];
                      reg367 <= (~&(&(^reg171)));
                      reg368 <= $unsigned((!(reg345 ?
                          (reg174 <= reg343) : reg287)));
                      reg369 <= reg105;
                    end
                  else
                    begin
                      reg366 <= $unsigned(({reg367[(1'h0):(1'h0)]} ?
                          reg239[(4'h9):(3'h4)] : (~{reg360})));
                      reg367 <= reg279[(1'h0):(1'h0)];
                    end
                end
            end
          for (forvar370 = (1'h0); (forvar370 < (2'h3)); forvar370 = (forvar370 + (1'h1)))
            begin
              for (forvar371 = (1'h0); (forvar371 < (1'h0)); forvar371 = (forvar371 + (1'h1)))
                begin
                  for (forvar372 = (1'h0); (forvar372 < (2'h2)); forvar372 = (forvar372 + (1'h1)))
                    begin
                      reg373 <= $unsigned((reg344[(1'h1):(1'h1)] | (reg315[(3'h4):(2'h3)] * (~^reg155))));
                      reg374 <= ({({reg143} ? reg360 : (~^reg280))} ?
                          (~^{(reg115 ? reg197 : reg332)}) : (~^(8'ha3)));
                    end
                  if (forvar272)
                    begin
                      reg375 <= ((reg129[(3'h4):(2'h2)] ?
                              ($unsigned(reg191) ?
                                  $signed(forvar292) : reg153) : $unsigned(reg233)) ?
                          (reg105 >= {$unsigned(forvar284)}) : reg315);
                    end
                  else
                    begin
                      reg375 <= (!({reg117[(2'h3):(2'h3)]} ?
                          {(reg225 ? forvar362 : reg209)} : ($signed((8'hb6)) ?
                              {forvar372} : reg285[(1'h0):(1'h0)])));
                      reg376 <= ((((reg310 & reg289) >> $unsigned(reg140)) <<< (reg339 ?
                              reg243 : reg183)) ?
                          (reg320[(4'h8):(3'h7)] ^~ (~(reg192 ?
                              reg285 : reg289))) : (((reg198 ?
                                  forvar335 : reg160) ?
                              $signed(reg320) : (forvar214 ?
                                  forvar257 : reg112)) != (reg226[(2'h2):(1'h1)] ?
                              reg211[(4'hd):(4'h8)] : forvar281[(3'h7):(2'h2)])));
                      reg377 <= (8'ha6);
                    end
                  if ((8'hac))
                    begin
                      reg378 <= reg293;
                      reg379 <= reg322;
                    end
                  else
                    begin
                      reg378 <= (~|((reg217[(1'h0):(1'h0)] <= forvar370[(3'h7):(3'h4)]) ?
                          $unsigned({forvar297}) : $unsigned((reg118 >> reg211))));
                      reg379 <= forvar364;
                      reg380 <= (~forvar276[(1'h1):(1'h0)]);
                    end
                end
              for (forvar381 = (1'h0); (forvar381 < (2'h2)); forvar381 = (forvar381 + (1'h1)))
                begin
                  for (forvar382 = (1'h0); (forvar382 < (1'h0)); forvar382 = (forvar382 + (1'h1)))
                    begin
                      reg383 <= $unsigned($signed($signed((&reg295))));
                    end
                  if ({((!forvar266) < $unsigned($signed(forvar224)))})
                    begin
                      reg384 <= ($unsigned($unsigned((reg162 >>> forvar309))) ?
                          $signed((~&$unsigned(reg194))) : (wire88 < (^~reg282)));
                      reg385 <= reg148[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg384 <= $signed($unsigned({(reg240 ?
                              forvar259 : reg218)}));
                      reg385 <= (8'h9d);
                      reg386 <= forvar245;
                    end
                  for (forvar387 = (1'h0); (forvar387 < (1'h1)); forvar387 = (forvar387 + (1'h1)))
                    begin
                      reg388 <= reg344;
                    end
                end
              if (reg104)
                begin
                  if ((forvar382 != (|forvar224[(1'h0):(1'h0)])))
                    begin
                      reg389 <= reg356[(2'h2):(2'h2)];
                      reg390 <= ($signed((~|$unsigned(reg369))) ?
                          $signed(reg250) : (^{reg321}));
                    end
                  else
                    begin
                      reg389 <= ((&reg250[(3'h4):(2'h3)]) ?
                          reg184 : (((forvar340 ? forvar362 : reg331) ?
                                  reg220[(1'h1):(1'h1)] : $unsigned(reg217)) ?
                              $signed(reg229[(3'h4):(2'h2)]) : (reg374 ?
                                  $unsigned((8'h9c)) : $signed(reg110))));
                    end
                  reg391 <= (((reg209 ?
                          reg356[(3'h4):(2'h3)] : reg262) ^ {(~|reg282)}) ?
                      ($unsigned(reg302) ?
                          $unsigned(((8'h9f) ?
                              reg244 : reg267)) : ($signed((8'hb5)) ?
                              $unsigned(reg184) : reg109)) : $unsigned($unsigned((|reg145))));
                end
              else
                begin
                  for (forvar389 = (1'h0); (forvar389 < (2'h3)); forvar389 = (forvar389 + (1'h1)))
                    begin
                      reg390 <= reg97;
                      reg391 <= $unsigned($unsigned(((reg177 ?
                          forvar309 : reg194) ^ (^~reg252))));
                      reg392 <= ($signed((reg274[(2'h2):(1'h1)] + {forvar206})) ?
                          {(8'ha1)} : reg314);
                      reg393 <= ($unsigned($signed($unsigned(reg321))) * reg184);
                    end
                end
              for (forvar394 = (1'h0); (forvar394 < (2'h3)); forvar394 = (forvar394 + (1'h1)))
                begin
                  for (forvar395 = (1'h0); (forvar395 < (2'h2)); forvar395 = (forvar395 + (1'h1)))
                    begin
                      reg396 <= ((~^(^(reg363 & forvar170))) & forvar289);
                      reg397 <= $signed((|({(8'had)} ?
                          (wire90 != (8'hb3)) : $unsigned(reg168))));
                    end
                  for (forvar398 = (1'h0); (forvar398 < (2'h2)); forvar398 = (forvar398 + (1'h1)))
                    begin
                      reg399 <= {reg122[(3'h4):(1'h0)]};
                      reg400 <= (&(~^($unsigned((8'h9c)) * (reg185 ?
                          forvar312 : reg282))));
                      reg401 <= reg136;
                      reg402 <= (~|$unsigned((reg215 ~^ ((8'hb2) & reg148))));
                    end
                  for (forvar403 = (1'h0); (forvar403 < (2'h2)); forvar403 = (forvar403 + (1'h1)))
                    begin
                      reg404 <= (~^(reg136 - reg177[(3'h5):(2'h2)]));
                    end
                end
            end
          for (forvar405 = (1'h0); (forvar405 < (1'h1)); forvar405 = (forvar405 + (1'h1)))
            begin
              if ($unsigned((~((forvar309 ? forvar206 : (8'hb5)) ?
                  reg243 : (reg109 - forvar293)))))
                begin
                  if ((|reg303))
                    begin
                      reg406 <= reg402;
                      reg407 <= (8'ha7);
                      reg408 <= ($unsigned(({wire89} ?
                          reg109 : reg244[(2'h3):(1'h0)])) > ($unsigned((reg113 * reg337)) ?
                          ($signed(reg361) ?
                              (~^(8'hb8)) : $unsigned((8'hb0))) : forvar363));
                    end
                  else
                    begin
                      reg406 <= $unsigned($unsigned(wire90));
                      reg407 <= (|$signed(reg290));
                      reg408 <= reg223[(3'h5):(3'h4)];
                      reg409 <= ((8'hac) ?
                          ($signed(reg105) ?
                              $signed({reg112}) : $signed(reg127)) : (^~((reg172 ?
                                  reg162 : wire89) ?
                              $signed(reg291) : $signed(reg341))));
                    end
                end
              else
                begin
                  if ({{$unsigned($unsigned(forvar363))}})
                    begin
                      reg406 <= (~|(wire90 ?
                          (&(forvar210 || reg146)) : $signed((8'hb4))));
                      reg407 <= (~^{$unsigned(reg205)});
                    end
                  else
                    begin
                      reg406 <= reg286[(3'h4):(3'h4)];
                      reg407 <= wire93;
                    end
                end
              for (forvar410 = (1'h0); (forvar410 < (2'h3)); forvar410 = (forvar410 + (1'h1)))
                begin
                  for (forvar411 = (1'h0); (forvar411 < (2'h2)); forvar411 = (forvar411 + (1'h1)))
                    begin
                      reg412 <= ({{{reg156}}} ?
                          $signed((reg392[(3'h5):(1'h0)] ?
                              (forvar245 ?
                                  reg180 : reg357) : reg404)) : (8'ha3));
                      reg413 <= $unsigned($unsigned(reg268[(4'h9):(3'h6)]));
                      reg414 <= ((8'haf) ^~ (~^(reg250[(1'h0):(1'h0)] ^ (reg324 ?
                          reg236 : (8'hb1)))));
                    end
                  for (forvar415 = (1'h0); (forvar415 < (1'h1)); forvar415 = (forvar415 + (1'h1)))
                    begin
                      reg416 <= {$unsigned(reg154[(3'h7):(3'h5)])};
                      reg417 <= ((&$unsigned(reg183)) ?
                          $signed(((&reg367) ~^ forvar179)) : {reg349[(1'h0):(1'h0)]});
                      reg418 <= $signed($signed((forvar389[(1'h1):(1'h0)] ^ $signed(reg167))));
                      reg419 <= forvar362[(2'h3):(1'h0)];
                    end
                  if ((^$unsigned((!(reg211 >>> reg322)))))
                    begin
                      reg420 <= ($signed(reg218) || forvar297[(3'h4):(1'h1)]);
                      reg421 <= reg302;
                      reg422 <= (({(~forvar307)} ?
                              (reg162[(1'h0):(1'h0)] == (8'ha5)) : ({reg258} || forvar356)) ?
                          reg244[(3'h5):(2'h2)] : (8'hb5));
                    end
                  else
                    begin
                      reg420 <= ($signed(($signed(reg363) ?
                          (^~reg376) : reg348)) <= $signed(reg237));
                      reg421 <= (forvar152 ?
                          $signed((!(forvar350 >>> reg330))) : reg229[(2'h3):(2'h2)]);
                      reg422 <= $signed(reg355);
                    end
                  for (forvar423 = (1'h0); (forvar423 < (1'h1)); forvar423 = (forvar423 + (1'h1)))
                    begin
                      reg424 <= reg337[(3'h5):(3'h4)];
                      reg425 <= forvar284[(3'h4):(3'h4)];
                      reg426 <= $signed($unsigned((~^reg363)));
                    end
                end
              reg427 <= reg397;
              for (forvar428 = (1'h0); (forvar428 < (1'h0)); forvar428 = (forvar428 + (1'h1)))
                begin
                  for (forvar429 = (1'h0); (forvar429 < (1'h1)); forvar429 = (forvar429 + (1'h1)))
                    begin
                      reg430 <= (-(|$unsigned(((8'hb5) ? forvar389 : reg315))));
                    end
                end
            end
        end
      for (forvar431 = (1'h0); (forvar431 < (2'h2)); forvar431 = (forvar431 + (1'h1)))
        begin
          for (forvar432 = (1'h0); (forvar432 < (1'h0)); forvar432 = (forvar432 + (1'h1)))
            begin
              for (forvar433 = (1'h0); (forvar433 < (1'h1)); forvar433 = (forvar433 + (1'h1)))
                begin
                  if ($signed(reg255))
                    begin
                      reg434 <= $signed(({reg360[(3'h5):(1'h1)]} ~^ $signed(((8'h9c) ?
                          reg199 : forvar271))));
                    end
                  else
                    begin
                      reg434 <= {reg258[(1'h1):(1'h0)]};
                      reg435 <= {$signed(reg300)};
                      reg436 <= $signed(({((8'ha8) ?
                              reg299 : reg243)} <= (!(reg341 < (8'haa)))));
                      reg437 <= ({($signed(reg318) ?
                              (reg215 ?
                                  (8'ha7) : (8'hb8)) : reg316[(4'hb):(4'hb)])} ^ reg142);
                    end
                  if ($signed(reg107[(2'h2):(2'h2)]))
                    begin
                      reg438 <= ({$signed(((8'ha2) ^~ reg374))} ?
                          ($unsigned($unsigned(reg194)) > $signed((reg413 || wire90))) : $unsigned((&(reg308 ?
                              reg223 : reg200))));
                      reg439 <= reg349;
                      reg440 <= $unsigned($unsigned(((reg302 ?
                          reg162 : reg283) >>> reg208)));
                      reg441 <= (^$unsigned($signed($unsigned(reg269))));
                    end
                  else
                    begin
                      reg438 <= $unsigned((^~forvar287[(4'h9):(3'h4)]));
                      reg439 <= (^~reg331[(2'h2):(1'h0)]);
                      reg440 <= reg417[(2'h3):(1'h1)];
                      reg441 <= (reg253[(3'h4):(1'h0)] ?
                          {$signed($signed(reg147))} : (~^(&(reg296 && forvar245))));
                    end
                  for (forvar442 = (1'h0); (forvar442 < (2'h2)); forvar442 = (forvar442 + (1'h1)))
                    begin
                      reg443 <= ($unsigned((~&wire91[(3'h5):(2'h2)])) ?
                          forvar210 : reg313);
                      reg444 <= {reg244};
                    end
                end
              if (reg287[(3'h5):(2'h3)])
                begin
                  if ($signed({($unsigned(reg439) == wire87)}))
                    begin
                      reg445 <= (-($unsigned(reg267) | reg260[(3'h4):(2'h2)]));
                      reg446 <= (^~(&($unsigned(reg437) != (reg288 < reg343))));
                    end
                  else
                    begin
                      reg445 <= reg143;
                      reg446 <= reg323[(2'h2):(1'h1)];
                      reg447 <= $signed($unsigned((reg328 || reg353)));
                    end
                  for (forvar448 = (1'h0); (forvar448 < (1'h1)); forvar448 = (forvar448 + (1'h1)))
                    begin
                      reg449 <= wire93[(3'h4):(1'h0)];
                      reg450 <= ({((reg357 | reg363) ?
                                  (forvar432 <<< forvar356) : {reg330})} ?
                          reg243 : ($unsigned(reg246) ~^ ($unsigned((8'hac)) ?
                              (~|forvar442) : {reg162})));
                      reg451 <= ((~&(+(8'hb5))) ?
                          (reg182 ?
                              ((forvar281 && (8'ha5)) ?
                                  (reg263 * (8'ha0)) : reg162) : $unsigned((^reg393))) : $unsigned(reg339[(3'h7):(1'h0)]));
                      reg452 <= $signed((((8'hae) ?
                          {(8'ha5)} : (wire90 <= reg413)) ^~ (^~((8'hb0) ?
                          forvar431 : reg248))));
                    end
                end
              else
                begin
                  for (forvar445 = (1'h0); (forvar445 < (1'h1)); forvar445 = (forvar445 + (1'h1)))
                    begin
                      reg446 <= {(~^($unsigned(reg350) >> (reg180 ?
                              reg376 : reg233)))};
                    end
                end
              for (forvar453 = (1'h0); (forvar453 < (1'h1)); forvar453 = (forvar453 + (1'h1)))
                begin
                  reg454 <= $unsigned(reg366[(4'hb):(1'h1)]);
                  for (forvar455 = (1'h0); (forvar455 < (2'h2)); forvar455 = (forvar455 + (1'h1)))
                    begin
                      reg456 <= (reg243[(1'h0):(1'h0)] ?
                          (reg353[(3'h7):(3'h7)] ?
                              reg215[(4'h9):(2'h2)] : ((forvar242 ?
                                      reg159 : reg341) ?
                                  $unsigned(reg426) : (forvar448 ^~ (8'ha5)))) : $signed(reg275));
                    end
                  if ((((~|(forvar394 ? reg285 : forvar309)) ?
                          (forvar242[(4'hf):(3'h4)] > reg279[(1'h1):(1'h1)]) : ((~&reg348) ?
                              (reg146 ? reg196 : reg142) : reg362)) ?
                      {(~^(reg174 ? reg225 : reg388))} : reg399))
                    begin
                      reg457 <= $unsigned({forvar306[(2'h3):(1'h0)]});
                      reg458 <= (reg97[(1'h0):(1'h0)] ?
                          (($signed(reg447) ?
                              (reg346 ?
                                  forvar272 : reg142) : forvar281) ~^ forvar372[(3'h5):(2'h3)]) : (((reg346 != (8'ha7)) ?
                                  $unsigned(reg273) : {reg396}) ?
                              forvar297 : $signed(((8'hac) <= reg113))));
                      reg459 <= reg338[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg457 <= {$unsigned(($signed(reg263) ^ {reg358}))};
                    end
                  for (forvar460 = (1'h0); (forvar460 < (2'h3)); forvar460 = (forvar460 + (1'h1)))
                    begin
                      reg461 <= (^reg195);
                    end
                end
              if (reg167)
                begin
                  for (forvar462 = (1'h0); (forvar462 < (2'h3)); forvar462 = (forvar462 + (1'h1)))
                    begin
                      reg463 <= ({($signed(forvar352) ?
                                  (-reg361) : (!reg194))} ?
                          (~|reg334) : $signed(reg195[(2'h3):(1'h0)]));
                      reg464 <= forvar228;
                      reg465 <= $signed(($signed({reg360}) > $signed((|reg263))));
                    end
                  for (forvar466 = (1'h0); (forvar466 < (1'h1)); forvar466 = (forvar466 + (1'h1)))
                    begin
                      reg467 <= reg416[(1'h0):(1'h0)];
                      reg468 <= reg390[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  if ((~($unsigned($unsigned((8'h9f))) ?
                      (~(forvar297 ^~ forvar428)) : forvar210[(2'h3):(2'h3)])))
                    begin
                      reg462 <= $unsigned((forvar206[(4'he):(1'h0)] == ((-forvar455) ?
                          (reg213 <<< reg148) : (^reg127))));
                      reg463 <= (reg247 - ((8'h9e) | (|$unsigned(reg238))));
                      reg464 <= reg221;
                    end
                  else
                    begin
                      reg462 <= $unsigned((~|(|$signed(reg97))));
                      reg463 <= reg371[(1'h0):(1'h0)];
                      reg464 <= (reg282[(2'h3):(2'h2)] ?
                          $signed({{reg222}}) : ({((8'hb7) ? reg391 : reg147)} ?
                              (&$signed(reg445)) : ($signed(reg370) << (reg393 * (8'h9c)))));
                    end
                  for (forvar465 = (1'h0); (forvar465 < (2'h3)); forvar465 = (forvar465 + (1'h1)))
                    begin
                      reg466 <= $unsigned({$signed({reg232})});
                    end
                  for (forvar467 = (1'h0); (forvar467 < (1'h1)); forvar467 = (forvar467 + (1'h1)))
                    begin
                      reg468 <= (^$unsigned(reg165));
                      reg469 <= $unsigned((&(|reg273)));
                    end
                  reg470 <= (!reg280);
                end
            end
          for (forvar471 = (1'h0); (forvar471 < (2'h3)); forvar471 = (forvar471 + (1'h1)))
            begin
              if ($signed({(~&$unsigned(reg109))}))
                begin
                  for (forvar472 = (1'h0); (forvar472 < (1'h0)); forvar472 = (forvar472 + (1'h1)))
                    begin
                      reg473 <= forvar257[(4'ha):(4'ha)];
                      reg474 <= $signed({((+reg269) ?
                              (reg294 == reg421) : (reg241 >>> reg247))});
                      reg475 <= (((~^{(8'h9d)}) ^~ reg145) ?
                          reg361 : reg359[(1'h1):(1'h1)]);
                    end
                  for (forvar476 = (1'h0); (forvar476 < (1'h0)); forvar476 = (forvar476 + (1'h1)))
                    begin
                      reg477 <= {reg456};
                      reg478 <= $unsigned(reg113[(1'h0):(1'h0)]);
                      reg479 <= forvar271;
                    end
                  if ((($unsigned((reg280 ? reg353 : forvar465)) ?
                      $unsigned(forvar152) : reg451) ^ reg110[(4'ha):(4'ha)]))
                    begin
                      reg480 <= (forvar432 >>> reg333[(4'hb):(1'h0)]);
                    end
                  else
                    begin
                      reg480 <= {($unsigned(((8'ha7) * reg351)) ?
                              ((reg207 > reg314) ?
                                  $unsigned(reg414) : (!reg182)) : reg384)};
                    end
                end
              else
                begin
                  for (forvar472 = (1'h0); (forvar472 < (2'h2)); forvar472 = (forvar472 + (1'h1)))
                    begin
                      reg473 <= $unsigned((forvar293 ?
                          ({reg379} ? {reg186} : (~&(8'ha1))) : forvar284));
                      reg474 <= reg371;
                      reg475 <= (((~^(-forvar297)) ?
                          (reg258[(2'h2):(2'h2)] ?
                              (-forvar307) : $signed(reg329)) : reg261[(3'h7):(2'h2)]) >> reg193[(1'h0):(1'h0)]);
                    end
                  for (forvar476 = (1'h0); (forvar476 < (2'h3)); forvar476 = (forvar476 + (1'h1)))
                    begin
                      reg477 <= $unsigned(({(~^forvar181)} ?
                          forvar455 : (~&reg231)));
                    end
                end
              for (forvar481 = (1'h0); (forvar481 < (2'h2)); forvar481 = (forvar481 + (1'h1)))
                begin
                  if ({(-(reg114 ?
                          $signed(forvar281) : forvar158[(2'h3):(2'h3)]))})
                    begin
                      reg482 <= reg186[(2'h3):(1'h1)];
                      reg483 <= (8'h9d);
                      reg484 <= $unsigned({$unsigned((~reg320))});
                      reg485 <= ((reg365 ?
                          wire90 : $unsigned($signed(reg300))) + $unsigned(((8'h9f) ^ $signed(forvar281))));
                    end
                  else
                    begin
                      reg482 <= forvar170;
                      reg483 <= (~(~&$signed((reg418 ^ reg304))));
                    end
                  reg486 <= ($signed($signed($unsigned(reg117))) << $signed($signed(((8'h9d) ?
                      reg271 : reg434))));
                end
            end
          for (forvar487 = (1'h0); (forvar487 < (1'h1)); forvar487 = (forvar487 + (1'h1)))
            begin
              if ($unsigned(wire89))
                begin
                  for (forvar488 = (1'h0); (forvar488 < (2'h2)); forvar488 = (forvar488 + (1'h1)))
                    begin
                      reg489 <= ((^~{$unsigned(reg383)}) ?
                          $signed($signed(reg241[(4'hd):(3'h4)])) : (~((-forvar245) ?
                              $signed((8'ha8)) : reg279[(2'h2):(1'h1)])));
                      reg490 <= reg344[(2'h2):(2'h2)];
                      reg491 <= (reg308[(3'h7):(3'h5)] ? reg409 : reg144);
                      reg492 <= ({(-(reg175 + (8'ha8)))} ?
                          ($signed($unsigned(reg316)) ?
                              $signed((forvar466 ?
                                  reg218 : forvar292)) : ((8'hb0) ^ (forvar265 ?
                                  (8'h9f) : reg180))) : reg466);
                    end
                end
              else
                begin
                  reg488 <= (~^$unsigned(reg254[(3'h4):(2'h3)]));
                  if ($unsigned({$signed(reg184[(2'h3):(2'h3)])}))
                    begin
                      reg489 <= wire91;
                      reg490 <= reg176[(1'h1):(1'h1)];
                      reg491 <= reg318;
                    end
                  else
                    begin
                      reg489 <= ((-reg295) * {(~&(forvar188 < reg196))});
                      reg490 <= reg478[(4'h8):(2'h2)];
                      reg491 <= $unsigned($unsigned(($signed(forvar465) ?
                          (reg319 ? reg365 : forvar242) : (forvar214 ?
                              forvar476 : reg392))));
                    end
                  if (reg386[(1'h1):(1'h0)])
                    begin
                      reg492 <= ($signed(reg166[(2'h2):(1'h1)]) ?
                          reg241[(2'h3):(2'h3)] : reg198[(3'h5):(3'h5)]);
                      reg493 <= $signed($signed((forvar364[(3'h7):(2'h2)] ?
                          reg274 : forvar344[(3'h4):(3'h4)])));
                      reg494 <= (|reg375);
                    end
                  else
                    begin
                      reg492 <= {reg358};
                      reg493 <= (((!reg391) ?
                          reg322[(3'h7):(3'h5)] : ((~^reg345) <= {reg292})) ~^ reg172);
                    end
                end
              reg495 <= {{(~|(reg360 - reg350))}};
              if ((reg401[(4'h9):(3'h6)] ?
                  $signed((&reg483)) : $unsigned($signed($unsigned((8'ha2))))))
                begin
                  reg496 <= ((&(((8'ha5) >> (8'hb1)) ~^ (~|forvar179))) >>> ((~&(reg478 & forvar206)) >> (8'hb5)));
                end
              else
                begin
                  for (forvar496 = (1'h0); (forvar496 < (2'h2)); forvar496 = (forvar496 + (1'h1)))
                    begin
                      reg497 <= ($signed(reg111[(4'ha):(1'h0)]) ?
                          reg462 : $signed($signed($signed(reg494))));
                      reg498 <= $unsigned((((reg191 <= reg107) ?
                              (8'hb1) : (~&reg169)) ?
                          $signed(forvar312) : reg129[(2'h3):(1'h0)]));
                      reg499 <= ((-(!reg116[(3'h6):(2'h3)])) > reg290);
                    end
                  if (reg140[(2'h2):(1'h1)])
                    begin
                      reg500 <= ({$signed((forvar460 + forvar433))} ?
                          ($signed((reg457 ?
                              reg389 : reg342)) || $signed(reg480)) : (forvar245 <= reg167));
                    end
                  else
                    begin
                      reg500 <= ({(-reg294[(2'h2):(1'h1)])} > (8'hb8));
                      reg501 <= (forvar259[(4'he):(3'h5)] ?
                          (^~forvar335) : reg187[(1'h0):(1'h0)]);
                      reg502 <= reg426[(1'h0):(1'h0)];
                    end
                  if (($signed(reg319) ?
                      ({(reg168 | reg454)} >>> $signed(forvar188)) : forvar423[(2'h2):(1'h0)]))
                    begin
                      reg503 <= $unsigned((reg211 && ($signed((8'hb3)) ?
                          $unsigned(reg209) : $unsigned(reg322))));
                    end
                  else
                    begin
                      reg503 <= ((-((~reg488) ?
                          {reg183} : (-forvar455))) | reg314[(1'h0):(1'h0)]);
                      reg504 <= reg413;
                      reg505 <= reg178;
                    end
                end
              if ({(~$unsigned($signed(reg327)))})
                begin
                  if ((^~$signed(reg144)))
                    begin
                      reg506 <= reg277;
                      reg507 <= $signed(reg420[(3'h4):(1'h1)]);
                      reg508 <= ((8'hb0) == $unsigned(($signed(reg299) << (&reg366))));
                    end
                  else
                    begin
                      reg506 <= ({(forvar462 ?
                              (~|reg370) : forvar462[(4'h9):(1'h1)])} || $signed($signed((~|(8'ha9)))));
                    end
                end
              else
                begin
                  for (forvar506 = (1'h0); (forvar506 < (1'h1)); forvar506 = (forvar506 + (1'h1)))
                    begin
                      reg507 <= (~|forvar467[(2'h2):(1'h0)]);
                    end
                end
            end
          reg509 <= (((reg222 ? reg148 : (8'ha5)) ?
                  reg110[(2'h2):(1'h0)] : ((~(8'hb0)) - (!reg464))) ?
              $signed(reg357) : $signed($signed(reg304[(2'h3):(2'h2)])));
        end
    end
  assign wire510 = {reg425[(2'h2):(1'h0)]};
  assign wire511 = (+(reg333 ?
                       (|(reg322 ? reg240 : reg195)) : reg293[(2'h3):(1'h0)]));
  assign wire512 = reg240[(3'h7):(1'h1)];
  module513 #() modinst719 (.wire514(reg446), .wire517(reg250), .wire518(reg491), .wire515(reg286), .y(wire718), .clk(clk), .wire516(reg140));
  assign wire720 = $unsigned($signed((8'hb5)));
  assign wire721 = $unsigned(reg497);
  module722 #() modinst3630 (wire3629, clk, reg379, reg342, reg438, reg242, reg364);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module722
#(parameter param3628 = (~&((&{(8'had)}) || {((8'ha1) >>> (8'ha2))})))
(y, clk, wire727, wire726, wire725, wire724, wire723);
  output wire [(32'hf40):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire727;
  input wire [(3'h5):(1'h0)] wire726;
  input wire [(2'h3):(1'h0)] wire725;
  input wire signed [(4'hf):(1'h0)] wire724;
  input wire [(2'h2):(1'h0)] wire723;
  wire signed [(3'h7):(1'h0)] wire3425;
  wire signed [(3'h6):(1'h0)] wire2033;
  wire [(2'h3):(1'h0)] wire2031;
  reg signed [(4'hb):(1'h0)] reg3627 = (1'h0);
  reg [(4'h8):(1'h0)] reg3626 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3625 = (1'h0);
  reg [(3'h6):(1'h0)] reg3624 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3623 = (1'h0);
  reg [(4'hc):(1'h0)] reg3621 = (1'h0);
  reg [(2'h2):(1'h0)] reg3620 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3619 = (1'h0);
  reg [(2'h2):(1'h0)] reg3618 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3617 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3616 = (1'h0);
  reg [(4'h8):(1'h0)] reg3615 = (1'h0);
  reg [(4'hc):(1'h0)] reg3614 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3612 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3611 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3610 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3608 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3607 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3606 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3605 = (1'h0);
  reg [(3'h7):(1'h0)] reg3602 = (1'h0);
  reg [(2'h2):(1'h0)] reg3601 = (1'h0);
  reg [(3'h4):(1'h0)] reg3600 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3599 = (1'h0);
  reg [(3'h5):(1'h0)] reg3598 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3597 = (1'h0);
  reg [(2'h2):(1'h0)] reg3595 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3594 = (1'h0);
  reg [(4'hf):(1'h0)] reg3593 = (1'h0);
  reg [(4'hd):(1'h0)] reg3592 = (1'h0);
  reg [(3'h4):(1'h0)] reg3591 = (1'h0);
  reg [(4'he):(1'h0)] reg3590 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3589 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3588 = (1'h0);
  reg [(3'h4):(1'h0)] reg3587 = (1'h0);
  reg [(4'h9):(1'h0)] reg3586 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3585 = (1'h0);
  reg [(4'hd):(1'h0)] reg3584 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3583 = (1'h0);
  reg [(4'h8):(1'h0)] reg3582 = (1'h0);
  reg [(5'h10):(1'h0)] reg3580 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3579 = (1'h0);
  reg [(3'h4):(1'h0)] reg3578 = (1'h0);
  reg [(4'h9):(1'h0)] reg3573 = (1'h0);
  reg [(4'hb):(1'h0)] reg3576 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3575 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3574 = (1'h0);
  reg [(3'h7):(1'h0)] reg3570 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3572 = (1'h0);
  reg [(4'he):(1'h0)] reg3571 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3561 = (1'h0);
  reg [(4'he):(1'h0)] reg3560 = (1'h0);
  reg [(2'h3):(1'h0)] reg3552 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3538 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3569 = (1'h0);
  reg [(4'h9):(1'h0)] reg3568 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3567 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3566 = (1'h0);
  reg [(2'h3):(1'h0)] reg3565 = (1'h0);
  reg [(2'h3):(1'h0)] reg3564 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3563 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3562 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3559 = (1'h0);
  reg [(4'hd):(1'h0)] reg3558 = (1'h0);
  reg [(3'h6):(1'h0)] reg3557 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3556 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3555 = (1'h0);
  reg [(4'h8):(1'h0)] reg3554 = (1'h0);
  reg [(4'h9):(1'h0)] reg3553 = (1'h0);
  reg [(2'h3):(1'h0)] reg3551 = (1'h0);
  reg [(4'h9):(1'h0)] reg3550 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3549 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3548 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3547 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3546 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3545 = (1'h0);
  reg [(3'h5):(1'h0)] reg3544 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3543 = (1'h0);
  reg [(3'h7):(1'h0)] reg3542 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3541 = (1'h0);
  reg [(4'hd):(1'h0)] reg3540 = (1'h0);
  reg [(4'hc):(1'h0)] reg3539 = (1'h0);
  reg [(3'h4):(1'h0)] reg3537 = (1'h0);
  reg [(4'h9):(1'h0)] reg3536 = (1'h0);
  reg [(3'h6):(1'h0)] reg3535 = (1'h0);
  reg [(5'h10):(1'h0)] reg3534 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3532 = (1'h0);
  reg [(3'h6):(1'h0)] reg3531 = (1'h0);
  reg [(2'h2):(1'h0)] reg3530 = (1'h0);
  reg [(3'h6):(1'h0)] reg3529 = (1'h0);
  reg [(4'hd):(1'h0)] reg3528 = (1'h0);
  reg [(4'hb):(1'h0)] reg3527 = (1'h0);
  reg [(4'ha):(1'h0)] reg3526 = (1'h0);
  reg [(4'hc):(1'h0)] reg3522 = (1'h0);
  reg [(4'hc):(1'h0)] reg3517 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3525 = (1'h0);
  reg [(5'h10):(1'h0)] reg3524 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3523 = (1'h0);
  reg [(3'h6):(1'h0)] reg3521 = (1'h0);
  reg [(4'h9):(1'h0)] reg3520 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3519 = (1'h0);
  reg [(4'hd):(1'h0)] reg3518 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3516 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3515 = (1'h0);
  reg [(4'ha):(1'h0)] reg3514 = (1'h0);
  reg [(5'h10):(1'h0)] reg3513 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3512 = (1'h0);
  reg [(3'h6):(1'h0)] reg3511 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3510 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3509 = (1'h0);
  reg [(2'h2):(1'h0)] reg3508 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3507 = (1'h0);
  reg [(2'h3):(1'h0)] reg3506 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3505 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3504 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3503 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3502 = (1'h0);
  reg [(2'h3):(1'h0)] reg3501 = (1'h0);
  reg [(2'h2):(1'h0)] reg3500 = (1'h0);
  reg [(4'hf):(1'h0)] reg3499 = (1'h0);
  reg [(4'ha):(1'h0)] reg3498 = (1'h0);
  reg [(4'h9):(1'h0)] reg3497 = (1'h0);
  reg [(4'hc):(1'h0)] reg3494 = (1'h0);
  reg [(3'h6):(1'h0)] reg3493 = (1'h0);
  reg [(3'h7):(1'h0)] reg3492 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3491 = (1'h0);
  reg [(4'h9):(1'h0)] reg3490 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3489 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3488 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3487 = (1'h0);
  reg [(4'hd):(1'h0)] reg3486 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3482 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3476 = (1'h0);
  reg [(3'h5):(1'h0)] reg3485 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3484 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3483 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3481 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3480 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3479 = (1'h0);
  reg [(3'h6):(1'h0)] reg3478 = (1'h0);
  reg [(4'ha):(1'h0)] reg3477 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3474 = (1'h0);
  reg [(5'h10):(1'h0)] reg3471 = (1'h0);
  reg [(4'hf):(1'h0)] reg3467 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3458 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3447 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3473 = (1'h0);
  reg [(4'hf):(1'h0)] reg3472 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3470 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3469 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3468 = (1'h0);
  reg [(3'h7):(1'h0)] reg3466 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3465 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3464 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3461 = (1'h0);
  reg [(4'hd):(1'h0)] reg3456 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3452 = (1'h0);
  reg [(4'h8):(1'h0)] reg3463 = (1'h0);
  reg [(3'h7):(1'h0)] reg3462 = (1'h0);
  reg [(3'h5):(1'h0)] reg3460 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3459 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3457 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3455 = (1'h0);
  reg [(3'h7):(1'h0)] reg3454 = (1'h0);
  reg [(4'ha):(1'h0)] reg3453 = (1'h0);
  reg [(4'hd):(1'h0)] reg3451 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3450 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3449 = (1'h0);
  reg [(4'hb):(1'h0)] reg3448 = (1'h0);
  reg [(2'h3):(1'h0)] reg3445 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3444 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3443 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3442 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3439 = (1'h0);
  reg [(3'h6):(1'h0)] reg3438 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3437 = (1'h0);
  reg [(2'h3):(1'h0)] reg3436 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3435 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3434 = (1'h0);
  reg [(4'hc):(1'h0)] reg3433 = (1'h0);
  reg [(4'hf):(1'h0)] reg3432 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3431 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3430 = (1'h0);
  reg [(4'hc):(1'h0)] reg3429 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg866 = (1'h0);
  reg signed [(4'he):(1'h0)] reg865 = (1'h0);
  reg [(3'h4):(1'h0)] reg864 = (1'h0);
  reg [(2'h3):(1'h0)] reg863 = (1'h0);
  reg [(4'hc):(1'h0)] reg861 = (1'h0);
  reg [(4'hf):(1'h0)] reg860 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg859 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg848 = (1'h0);
  reg [(3'h6):(1'h0)] reg856 = (1'h0);
  reg [(3'h5):(1'h0)] reg855 = (1'h0);
  reg signed [(4'he):(1'h0)] reg854 = (1'h0);
  reg [(4'hf):(1'h0)] reg853 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg852 = (1'h0);
  reg [(4'he):(1'h0)] reg851 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg850 = (1'h0);
  reg [(5'h10):(1'h0)] reg849 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg838 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg837 = (1'h0);
  reg [(4'he):(1'h0)] reg835 = (1'h0);
  reg [(4'ha):(1'h0)] reg830 = (1'h0);
  reg [(4'he):(1'h0)] reg846 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg845 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg844 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg843 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg841 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg840 = (1'h0);
  reg [(2'h2):(1'h0)] reg839 = (1'h0);
  reg [(2'h3):(1'h0)] reg836 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg834 = (1'h0);
  reg [(3'h6):(1'h0)] reg833 = (1'h0);
  reg [(4'hf):(1'h0)] reg832 = (1'h0);
  reg [(3'h6):(1'h0)] reg831 = (1'h0);
  reg signed [(4'he):(1'h0)] reg829 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg828 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg827 = (1'h0);
  reg signed [(4'he):(1'h0)] reg825 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg824 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg823 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg822 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg821 = (1'h0);
  reg [(4'hb):(1'h0)] reg820 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg819 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg818 = (1'h0);
  reg [(4'he):(1'h0)] reg812 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg817 = (1'h0);
  reg [(4'hc):(1'h0)] reg816 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg815 = (1'h0);
  reg [(2'h2):(1'h0)] reg814 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg813 = (1'h0);
  reg [(2'h2):(1'h0)] reg758 = (1'h0);
  reg [(3'h5):(1'h0)] reg752 = (1'h0);
  reg [(5'h10):(1'h0)] reg742 = (1'h0);
  reg [(4'hc):(1'h0)] reg810 = (1'h0);
  reg [(3'h6):(1'h0)] reg805 = (1'h0);
  reg [(5'h10):(1'h0)] reg796 = (1'h0);
  reg [(2'h2):(1'h0)] reg794 = (1'h0);
  reg [(3'h6):(1'h0)] reg809 = (1'h0);
  reg signed [(4'he):(1'h0)] reg808 = (1'h0);
  reg [(2'h3):(1'h0)] reg807 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg806 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg803 = (1'h0);
  reg [(5'h10):(1'h0)] reg802 = (1'h0);
  reg signed [(4'he):(1'h0)] reg801 = (1'h0);
  reg [(5'h10):(1'h0)] reg800 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg799 = (1'h0);
  reg [(3'h7):(1'h0)] reg798 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg797 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg795 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg793 = (1'h0);
  reg [(4'he):(1'h0)] reg792 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg791 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg790 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg788 = (1'h0);
  reg [(4'he):(1'h0)] reg787 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg786 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg785 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg784 = (1'h0);
  reg [(4'hc):(1'h0)] reg783 = (1'h0);
  reg [(4'ha):(1'h0)] reg782 = (1'h0);
  reg [(3'h4):(1'h0)] reg781 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg780 = (1'h0);
  reg [(4'hd):(1'h0)] reg779 = (1'h0);
  reg [(4'he):(1'h0)] reg777 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg776 = (1'h0);
  reg [(4'hc):(1'h0)] reg775 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg774 = (1'h0);
  reg [(4'h8):(1'h0)] reg773 = (1'h0);
  reg [(3'h6):(1'h0)] reg772 = (1'h0);
  reg [(5'h10):(1'h0)] reg771 = (1'h0);
  reg [(3'h4):(1'h0)] reg770 = (1'h0);
  reg [(3'h5):(1'h0)] reg769 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg768 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg765 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg764 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg763 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg762 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg761 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg760 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg759 = (1'h0);
  reg [(4'hd):(1'h0)] reg757 = (1'h0);
  reg [(3'h5):(1'h0)] reg747 = (1'h0);
  reg [(4'ha):(1'h0)] reg756 = (1'h0);
  reg [(4'hc):(1'h0)] reg755 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg754 = (1'h0);
  reg [(4'ha):(1'h0)] reg753 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg751 = (1'h0);
  reg [(3'h4):(1'h0)] reg750 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg749 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg748 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg746 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg745 = (1'h0);
  reg [(4'h8):(1'h0)] reg744 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg743 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg741 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg740 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg739 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg738 = (1'h0);
  reg [(4'hb):(1'h0)] reg737 = (1'h0);
  reg [(4'ha):(1'h0)] reg736 = (1'h0);
  reg [(4'hc):(1'h0)] reg735 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg734 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg733 = (1'h0);
  reg signed [(4'he):(1'h0)] reg732 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg731 = (1'h0);
  reg [(5'h10):(1'h0)] reg730 = (1'h0);
  reg signed [(4'he):(1'h0)] reg729 = (1'h0);
  reg [(3'h7):(1'h0)] reg728 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3622 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3613 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3609 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3604 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3603 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3590 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3591 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3596 = (1'h0);
  reg [(4'he):(1'h0)] forvar3581 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3577 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3576 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3573 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3570 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3559 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3558 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3553 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3549 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3545 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3530 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3527 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3526 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3561 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3560 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3548 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3552 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3531 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3538 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3533 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3518 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3512 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3522 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3517 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3513 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3496 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3495 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3486 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3482 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3476 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3475 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3464 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3468 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3465 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3449 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3471 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3467 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3453 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3450 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3461 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3458 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3456 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3452 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3447 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3446 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3441 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3440 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3428 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3427 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar862 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar858 = (1'h0);
  reg [(5'h10):(1'h0)] forvar857 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar848 = (1'h0);
  reg [(3'h5):(1'h0)] forvar847 = (1'h0);
  reg [(2'h2):(1'h0)] forvar840 = (1'h0);
  reg [(4'he):(1'h0)] forvar836 = (1'h0);
  reg [(4'hb):(1'h0)] forvar834 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar831 = (1'h0);
  reg [(3'h7):(1'h0)] forvar842 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar838 = (1'h0);
  reg [(4'hc):(1'h0)] forvar837 = (1'h0);
  reg [(5'h10):(1'h0)] forvar835 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar830 = (1'h0);
  reg [(4'ha):(1'h0)] forvar822 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar826 = (1'h0);
  reg [(4'h9):(1'h0)] forvar814 = (1'h0);
  reg [(4'hd):(1'h0)] forvar812 = (1'h0);
  reg [(2'h2):(1'h0)] forvar811 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar764 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar761 = (1'h0);
  reg [(3'h6):(1'h0)] forvar760 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar753 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar751 = (1'h0);
  reg [(3'h7):(1'h0)] forvar749 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar748 = (1'h0);
  reg [(4'h9):(1'h0)] forvar743 = (1'h0);
  reg [(4'hc):(1'h0)] forvar739 = (1'h0);
  reg [(3'h4):(1'h0)] forvar730 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar808 = (1'h0);
  reg [(4'h8):(1'h0)] forvar800 = (1'h0);
  reg [(2'h2):(1'h0)] forvar795 = (1'h0);
  reg [(4'h8):(1'h0)] forvar790 = (1'h0);
  reg [(4'ha):(1'h0)] forvar805 = (1'h0);
  reg [(4'ha):(1'h0)] forvar804 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar796 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar794 = (1'h0);
  reg [(4'hc):(1'h0)] forvar789 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar778 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar773 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar767 = (1'h0);
  reg [(5'h10):(1'h0)] forvar766 = (1'h0);
  reg [(4'he):(1'h0)] forvar759 = (1'h0);
  reg [(5'h10):(1'h0)] forvar758 = (1'h0);
  reg [(5'h10):(1'h0)] forvar746 = (1'h0);
  reg [(5'h10):(1'h0)] forvar752 = (1'h0);
  reg [(3'h4):(1'h0)] forvar747 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar742 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar735 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar732 = (1'h0);
  assign y = {wire3425,
                 wire2033,
                 wire2031,
                 reg3627,
                 reg3626,
                 reg3625,
                 reg3624,
                 reg3623,
                 reg3621,
                 reg3620,
                 reg3619,
                 reg3618,
                 reg3617,
                 reg3616,
                 reg3615,
                 reg3614,
                 reg3612,
                 reg3611,
                 reg3610,
                 reg3608,
                 reg3607,
                 reg3606,
                 reg3605,
                 reg3602,
                 reg3601,
                 reg3600,
                 reg3599,
                 reg3598,
                 reg3597,
                 reg3595,
                 reg3594,
                 reg3593,
                 reg3592,
                 reg3591,
                 reg3590,
                 reg3589,
                 reg3588,
                 reg3587,
                 reg3586,
                 reg3585,
                 reg3584,
                 reg3583,
                 reg3582,
                 reg3580,
                 reg3579,
                 reg3578,
                 reg3573,
                 reg3576,
                 reg3575,
                 reg3574,
                 reg3570,
                 reg3572,
                 reg3571,
                 reg3561,
                 reg3560,
                 reg3552,
                 reg3538,
                 reg3569,
                 reg3568,
                 reg3567,
                 reg3566,
                 reg3565,
                 reg3564,
                 reg3563,
                 reg3562,
                 reg3559,
                 reg3558,
                 reg3557,
                 reg3556,
                 reg3555,
                 reg3554,
                 reg3553,
                 reg3551,
                 reg3550,
                 reg3549,
                 reg3548,
                 reg3547,
                 reg3546,
                 reg3545,
                 reg3544,
                 reg3543,
                 reg3542,
                 reg3541,
                 reg3540,
                 reg3539,
                 reg3537,
                 reg3536,
                 reg3535,
                 reg3534,
                 reg3532,
                 reg3531,
                 reg3530,
                 reg3529,
                 reg3528,
                 reg3527,
                 reg3526,
                 reg3522,
                 reg3517,
                 reg3525,
                 reg3524,
                 reg3523,
                 reg3521,
                 reg3520,
                 reg3519,
                 reg3518,
                 reg3516,
                 reg3515,
                 reg3514,
                 reg3513,
                 reg3512,
                 reg3511,
                 reg3510,
                 reg3509,
                 reg3508,
                 reg3507,
                 reg3506,
                 reg3505,
                 reg3504,
                 reg3503,
                 reg3502,
                 reg3501,
                 reg3500,
                 reg3499,
                 reg3498,
                 reg3497,
                 reg3494,
                 reg3493,
                 reg3492,
                 reg3491,
                 reg3490,
                 reg3489,
                 reg3488,
                 reg3487,
                 reg3486,
                 reg3482,
                 reg3476,
                 reg3485,
                 reg3484,
                 reg3483,
                 reg3481,
                 reg3480,
                 reg3479,
                 reg3478,
                 reg3477,
                 reg3474,
                 reg3471,
                 reg3467,
                 reg3458,
                 reg3447,
                 reg3473,
                 reg3472,
                 reg3470,
                 reg3469,
                 reg3468,
                 reg3466,
                 reg3465,
                 reg3464,
                 reg3461,
                 reg3456,
                 reg3452,
                 reg3463,
                 reg3462,
                 reg3460,
                 reg3459,
                 reg3457,
                 reg3455,
                 reg3454,
                 reg3453,
                 reg3451,
                 reg3450,
                 reg3449,
                 reg3448,
                 reg3445,
                 reg3444,
                 reg3443,
                 reg3442,
                 reg3439,
                 reg3438,
                 reg3437,
                 reg3436,
                 reg3435,
                 reg3434,
                 reg3433,
                 reg3432,
                 reg3431,
                 reg3430,
                 reg3429,
                 reg866,
                 reg865,
                 reg864,
                 reg863,
                 reg861,
                 reg860,
                 reg859,
                 reg848,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 reg852,
                 reg851,
                 reg850,
                 reg849,
                 reg838,
                 reg837,
                 reg835,
                 reg830,
                 reg846,
                 reg845,
                 reg844,
                 reg843,
                 reg841,
                 reg840,
                 reg839,
                 reg836,
                 reg834,
                 reg833,
                 reg832,
                 reg831,
                 reg829,
                 reg828,
                 reg827,
                 reg825,
                 reg824,
                 reg823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 reg818,
                 reg812,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 reg758,
                 reg752,
                 reg742,
                 reg810,
                 reg805,
                 reg796,
                 reg794,
                 reg809,
                 reg808,
                 reg807,
                 reg806,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 reg798,
                 reg797,
                 reg795,
                 reg793,
                 reg792,
                 reg791,
                 reg790,
                 reg788,
                 reg787,
                 reg786,
                 reg785,
                 reg784,
                 reg783,
                 reg782,
                 reg781,
                 reg780,
                 reg779,
                 reg777,
                 reg776,
                 reg775,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 reg769,
                 reg768,
                 reg765,
                 reg764,
                 reg763,
                 reg762,
                 reg761,
                 reg760,
                 reg759,
                 reg757,
                 reg747,
                 reg756,
                 reg755,
                 reg754,
                 reg753,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg746,
                 reg745,
                 reg744,
                 reg743,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 reg730,
                 reg729,
                 reg728,
                 forvar3622,
                 forvar3613,
                 forvar3609,
                 forvar3604,
                 forvar3603,
                 forvar3590,
                 forvar3591,
                 forvar3596,
                 forvar3581,
                 forvar3577,
                 forvar3576,
                 forvar3573,
                 forvar3570,
                 forvar3559,
                 forvar3558,
                 forvar3553,
                 forvar3549,
                 forvar3545,
                 forvar3530,
                 forvar3527,
                 forvar3526,
                 forvar3561,
                 forvar3560,
                 forvar3548,
                 forvar3552,
                 forvar3531,
                 forvar3538,
                 forvar3533,
                 forvar3518,
                 forvar3512,
                 forvar3522,
                 forvar3517,
                 forvar3513,
                 forvar3496,
                 forvar3495,
                 forvar3486,
                 forvar3482,
                 forvar3476,
                 forvar3475,
                 forvar3464,
                 forvar3468,
                 forvar3465,
                 forvar3449,
                 forvar3471,
                 forvar3467,
                 forvar3453,
                 forvar3450,
                 forvar3461,
                 forvar3458,
                 forvar3456,
                 forvar3452,
                 forvar3447,
                 forvar3446,
                 forvar3441,
                 forvar3440,
                 forvar3428,
                 forvar3427,
                 forvar862,
                 forvar858,
                 forvar857,
                 forvar848,
                 forvar847,
                 forvar840,
                 forvar836,
                 forvar834,
                 forvar831,
                 forvar842,
                 forvar838,
                 forvar837,
                 forvar835,
                 forvar830,
                 forvar822,
                 forvar826,
                 forvar814,
                 forvar812,
                 forvar811,
                 forvar764,
                 forvar761,
                 forvar760,
                 forvar753,
                 forvar751,
                 forvar749,
                 forvar748,
                 forvar743,
                 forvar739,
                 forvar730,
                 forvar808,
                 forvar800,
                 forvar795,
                 forvar790,
                 forvar805,
                 forvar804,
                 forvar796,
                 forvar794,
                 forvar789,
                 forvar778,
                 forvar773,
                 forvar767,
                 forvar766,
                 forvar759,
                 forvar758,
                 forvar746,
                 forvar752,
                 forvar747,
                 forvar742,
                 forvar735,
                 forvar732,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg728 <= {wire725};
      reg729 <= ((wire723[(2'h2):(1'h1)] & (8'ha3)) ?
          wire723[(1'h0):(1'h0)] : wire726[(2'h2):(1'h1)]);
      if (wire725)
        begin
          reg730 <= $unsigned($signed(wire727[(4'hd):(2'h2)]));
          if (((reg730[(4'hf):(3'h5)] ? (8'hab) : {((8'hb0) | reg729)}) ?
              wire727 : ($unsigned({wire727}) > ($unsigned(wire726) ?
                  wire723[(2'h2):(2'h2)] : (reg728 ? wire725 : reg730)))))
            begin
              reg731 <= (!($unsigned($unsigned(reg730)) == wire724));
              if ((wire727[(1'h0):(1'h0)] & ({$signed(wire726)} >>> (8'ha9))))
                begin
                  if ({(wire723 & (~(wire725 >> (8'ha1))))})
                    begin
                      reg732 <= $unsigned((((~reg731) ?
                          $unsigned(reg728) : reg728[(3'h5):(1'h0)]) | reg728[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg732 <= wire727;
                    end
                  if (wire723[(2'h2):(2'h2)])
                    begin
                      reg733 <= (!(!(((8'ha7) ? reg732 : reg732) >>> reg732)));
                      reg734 <= $unsigned($signed(reg730));
                    end
                  else
                    begin
                      reg733 <= (wire723[(2'h2):(1'h0)] ?
                          $signed((wire723[(1'h0):(1'h0)] ^~ reg730)) : $signed($unsigned($signed((8'hb1)))));
                    end
                  reg735 <= $unsigned(reg732[(2'h3):(2'h2)]);
                end
              else
                begin
                  for (forvar732 = (1'h0); (forvar732 < (1'h0)); forvar732 = (forvar732 + (1'h1)))
                    begin
                      reg733 <= ($unsigned(reg733) ?
                          (&($signed(forvar732) ?
                              ((8'ha3) ?
                                  (8'ha8) : (8'ha1)) : $unsigned(reg733))) : $unsigned($signed((reg730 ?
                              wire727 : wire724))));
                      reg734 <= wire724[(4'h9):(3'h6)];
                    end
                  for (forvar735 = (1'h0); (forvar735 < (1'h1)); forvar735 = (forvar735 + (1'h1)))
                    begin
                      reg736 <= {reg732};
                      reg737 <= reg736[(1'h0):(1'h0)];
                      reg738 <= {$signed($signed(wire723))};
                    end
                  if ($unsigned((8'ha8)))
                    begin
                      reg739 <= {($signed(wire723) ?
                              $unsigned((^reg729)) : ((~^reg729) ?
                                  $signed(reg738) : wire726))};
                      reg740 <= (~^({wire726} <<< $unsigned($signed(forvar732))));
                      reg741 <= $unsigned(reg732[(3'h6):(2'h3)]);
                    end
                  else
                    begin
                      reg739 <= {reg733[(1'h0):(1'h0)]};
                    end
                  for (forvar742 = (1'h0); (forvar742 < (1'h0)); forvar742 = (forvar742 + (1'h1)))
                    begin
                      reg743 <= (($signed(reg739[(1'h1):(1'h0)]) >= reg738) ?
                          $signed({reg736}) : $unsigned(({(8'h9e)} ?
                              (8'hb3) : $signed(forvar735))));
                      reg744 <= reg739[(1'h1):(1'h0)];
                      reg745 <= {(|(8'ha0))};
                    end
                end
              if ((!wire723))
                begin
                  reg746 <= wire724;
                  for (forvar747 = (1'h0); (forvar747 < (1'h1)); forvar747 = (forvar747 + (1'h1)))
                    begin
                      reg748 <= $signed((8'hb2));
                      reg749 <= (reg741[(4'h9):(3'h4)] <<< (~&(-(reg743 >>> (8'h9e)))));
                      reg750 <= (({(~reg748)} ^~ ((reg740 & reg748) ?
                          reg748 : $signed(forvar742))) == $unsigned(reg735[(4'hc):(2'h2)]));
                      reg751 <= wire726[(1'h1):(1'h1)];
                    end
                  for (forvar752 = (1'h0); (forvar752 < (2'h3)); forvar752 = (forvar752 + (1'h1)))
                    begin
                      reg753 <= reg732[(4'ha):(4'ha)];
                      reg754 <= reg750;
                      reg755 <= $unsigned(reg737[(1'h0):(1'h0)]);
                      reg756 <= {$signed(reg745)};
                    end
                end
              else
                begin
                  for (forvar746 = (1'h0); (forvar746 < (1'h1)); forvar746 = (forvar746 + (1'h1)))
                    begin
                      reg747 <= reg750;
                      reg748 <= (|$unsigned((!wire724[(1'h0):(1'h0)])));
                    end
                end
              reg757 <= $signed(reg756[(3'h5):(3'h5)]);
            end
          else
            begin
              reg731 <= ((^~(8'ha0)) - (8'haf));
            end
          for (forvar758 = (1'h0); (forvar758 < (1'h1)); forvar758 = (forvar758 + (1'h1)))
            begin
              if ((reg740 + {$unsigned((reg729 ? reg749 : forvar747))}))
                begin
                  reg759 <= forvar747;
                end
              else
                begin
                  for (forvar759 = (1'h0); (forvar759 < (1'h1)); forvar759 = (forvar759 + (1'h1)))
                    begin
                      reg760 <= reg733;
                      reg761 <= $signed($signed((&((8'ha4) ^ reg754))));
                    end
                  if (((reg741[(2'h2):(1'h1)] ?
                          ((forvar747 < reg756) <<< $unsigned((8'h9c))) : wire723) ?
                      $signed($signed($unsigned(reg748))) : $signed(reg761[(4'hb):(4'h8)])))
                    begin
                      reg762 <= reg755[(1'h0):(1'h0)];
                      reg763 <= ({(reg730[(4'hf):(4'hd)] || $signed(reg757))} ?
                          reg732 : reg738[(4'h8):(3'h6)]);
                      reg764 <= reg730;
                      reg765 <= reg755[(4'h8):(1'h0)];
                    end
                  else
                    begin
                      reg762 <= forvar735;
                      reg763 <= (reg741[(3'h6):(2'h3)] == $signed((reg730 ?
                          (reg745 >= reg737) : reg761)));
                    end
                end
              for (forvar766 = (1'h0); (forvar766 < (1'h1)); forvar766 = (forvar766 + (1'h1)))
                begin
                  for (forvar767 = (1'h0); (forvar767 < (1'h0)); forvar767 = (forvar767 + (1'h1)))
                    begin
                      reg768 <= forvar747[(2'h3):(1'h0)];
                      reg769 <= forvar735[(1'h0):(1'h0)];
                      reg770 <= wire723[(1'h1):(1'h0)];
                      reg771 <= (((~forvar735[(1'h1):(1'h1)]) <<< forvar767) ^ ($signed($unsigned((8'hb0))) >>> ((wire724 + reg770) ?
                          (reg759 >>> (8'ha6)) : reg750[(3'h4):(1'h0)])));
                    end
                end
              reg772 <= (|{$unsigned($unsigned(forvar767))});
              if ((~reg737))
                begin
                  reg773 <= $unsigned(reg768);
                  if ((8'hb8))
                    begin
                      reg774 <= forvar759;
                      reg775 <= reg757;
                      reg776 <= reg749;
                      reg777 <= $signed($signed(forvar758[(3'h4):(2'h3)]));
                    end
                  else
                    begin
                      reg774 <= $unsigned(reg751[(3'h7):(1'h0)]);
                      reg775 <= ($signed((|(reg756 + (8'haf)))) ?
                          reg744[(4'h8):(3'h7)] : $unsigned((~(reg750 ~^ (8'hb3)))));
                      reg776 <= forvar758;
                      reg777 <= reg768[(2'h3):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar773 = (1'h0); (forvar773 < (1'h1)); forvar773 = (forvar773 + (1'h1)))
                    begin
                      reg774 <= (^~(reg770[(1'h0):(1'h0)] ?
                          ({reg759} ?
                              (forvar732 ^ reg745) : (|reg765)) : forvar767));
                      reg775 <= ($unsigned(reg755[(4'hc):(3'h4)]) ?
                          $unsigned((8'hac)) : (((wire726 + (8'hba)) & reg732) ?
                              $unsigned((-(8'h9c))) : $signed({reg735})));
                      reg776 <= $unsigned(($signed(reg763[(4'h8):(2'h3)]) ?
                          ((reg731 * reg751) || $unsigned(reg765)) : $signed($unsigned(reg768))));
                      reg777 <= ($signed($signed(reg733[(2'h3):(2'h3)])) == ($signed((~&reg740)) * $signed(reg775[(4'hc):(3'h5)])));
                    end
                  for (forvar778 = (1'h0); (forvar778 < (1'h0)); forvar778 = (forvar778 + (1'h1)))
                    begin
                      reg779 <= $signed((~^$unsigned((reg753 ?
                          reg777 : (8'h9e)))));
                      reg780 <= reg740;
                      reg781 <= $signed((-forvar752));
                    end
                  if ({((+{reg754}) - (-$unsigned(reg750)))})
                    begin
                      reg782 <= reg761;
                    end
                  else
                    begin
                      reg782 <= (8'ha4);
                      reg783 <= $signed(reg757);
                      reg784 <= $signed(($unsigned((reg749 == wire727)) >> ((8'hb2) && reg745)));
                    end
                  if ($signed((~|forvar747)))
                    begin
                      reg785 <= reg736[(3'h4):(2'h2)];
                      reg786 <= ($unsigned(((reg731 <= wire725) ?
                          reg764[(1'h1):(1'h1)] : reg744)) | {(forvar746[(4'h8):(3'h6)] ?
                              reg771[(3'h4):(1'h1)] : (reg761 ?
                                  reg743 : reg747))});
                      reg787 <= reg774[(2'h2):(1'h1)];
                      reg788 <= (|$signed((8'hb5)));
                    end
                  else
                    begin
                      reg785 <= $unsigned($unsigned(((reg734 ?
                              wire723 : forvar766) ?
                          $unsigned(reg735) : (!reg745))));
                    end
                end
            end
          if ((~^(|($unsigned(reg747) ^~ $unsigned(reg737)))))
            begin
              for (forvar789 = (1'h0); (forvar789 < (1'h1)); forvar789 = (forvar789 + (1'h1)))
                begin
                  if ($signed(reg740[(3'h6):(2'h3)]))
                    begin
                      reg790 <= forvar742;
                      reg791 <= (|$unsigned(((wire724 ?
                          reg785 : reg753) + reg780)));
                      reg792 <= (((|$signed(reg776)) ?
                              $unsigned($unsigned(reg741)) : reg785) ?
                          (~|reg751[(3'h5):(2'h3)]) : reg772);
                      reg793 <= ($unsigned($unsigned($signed((8'h9f)))) << reg762[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg790 <= ($unsigned(((reg786 ? reg756 : reg748) ?
                          (&forvar747) : (reg790 << reg740))) + $unsigned((((8'hb7) - (8'hb6)) || $unsigned((8'ha4)))));
                      reg791 <= (reg741 ?
                          $signed(({reg793} & $unsigned(reg729))) : (-(8'hb4)));
                    end
                  for (forvar794 = (1'h0); (forvar794 < (1'h0)); forvar794 = (forvar794 + (1'h1)))
                    begin
                      reg795 <= ((reg731 ?
                              reg776[(3'h6):(3'h6)] : (reg730 ?
                                  (reg732 ? (8'ha4) : (8'ha6)) : (~&(8'h9e)))) ?
                          (8'h9f) : ((8'hb8) && ((~^reg783) ~^ forvar752)));
                    end
                  for (forvar796 = (1'h0); (forvar796 < (2'h2)); forvar796 = (forvar796 + (1'h1)))
                    begin
                      reg797 <= {reg772[(2'h3):(2'h3)]};
                      reg798 <= ((8'hb2) ? reg773 : wire726);
                      reg799 <= reg750;
                    end
                end
              if (((8'hab) | $signed(wire726)))
                begin
                  reg800 <= (8'hb6);
                  if ((($signed((forvar742 ?
                      (8'ha0) : reg772)) & $unsigned(reg779[(1'h1):(1'h0)])) > (reg797[(3'h5):(1'h0)] ?
                      reg732[(4'ha):(1'h0)] : (reg773[(1'h0):(1'h0)] ^~ $unsigned(reg762)))))
                    begin
                      reg801 <= $unsigned(($unsigned(reg792[(4'ha):(2'h2)]) >>> forvar742));
                      reg802 <= forvar747;
                      reg803 <= $signed($signed($unsigned((reg744 ?
                          (8'ha1) : reg768))));
                    end
                  else
                    begin
                      reg801 <= ($signed($signed(reg739[(3'h5):(1'h1)])) + {(8'had)});
                      reg802 <= reg731;
                    end
                end
              else
                begin
                  if ($signed(reg747[(3'h4):(3'h4)]))
                    begin
                      reg800 <= reg728;
                      reg801 <= (forvar732 ?
                          wire727[(4'hb):(4'h8)] : ((&(reg740 == reg801)) * (^~(reg743 ~^ reg734))));
                      reg802 <= ((reg772[(1'h1):(1'h1)] == ((reg761 ?
                          reg747 : (8'hb0)) && (forvar767 <<< reg731))) >> (^($signed((8'haf)) ?
                          reg749[(2'h3):(1'h1)] : forvar752[(1'h0):(1'h0)])));
                      reg803 <= reg799;
                    end
                  else
                    begin
                      reg800 <= (~^$unsigned(reg768[(2'h3):(2'h2)]));
                    end
                end
              for (forvar804 = (1'h0); (forvar804 < (2'h3)); forvar804 = (forvar804 + (1'h1)))
                begin
                  for (forvar805 = (1'h0); (forvar805 < (2'h2)); forvar805 = (forvar805 + (1'h1)))
                    begin
                      reg806 <= $unsigned(forvar758);
                      reg807 <= (^((8'hb1) ? (^~$unsigned(reg765)) : (8'ha0)));
                      reg808 <= (reg768[(2'h2):(2'h2)] ^~ (reg768[(4'hb):(3'h6)] ?
                          $unsigned((-reg751)) : $signed($unsigned(reg749))));
                      reg809 <= ((8'hb9) ^ forvar759);
                    end
                end
            end
          else
            begin
              for (forvar789 = (1'h0); (forvar789 < (2'h2)); forvar789 = (forvar789 + (1'h1)))
                begin
                  for (forvar790 = (1'h0); (forvar790 < (1'h1)); forvar790 = (forvar790 + (1'h1)))
                    begin
                      reg791 <= (~^$signed($signed($signed(forvar805))));
                    end
                  if (reg798[(2'h2):(1'h1)])
                    begin
                      reg792 <= reg757[(3'h7):(3'h7)];
                    end
                  else
                    begin
                      reg792 <= reg768;
                      reg793 <= $unsigned({{$unsigned(forvar767)}});
                      reg794 <= $signed(reg774[(2'h3):(1'h0)]);
                    end
                end
              for (forvar795 = (1'h0); (forvar795 < (2'h3)); forvar795 = (forvar795 + (1'h1)))
                begin
                  if (forvar796[(3'h4):(1'h1)])
                    begin
                      reg796 <= forvar767[(3'h4):(1'h1)];
                      reg797 <= (((~|reg739) && $signed((reg754 <= (8'hb9)))) ?
                          ({forvar778[(4'hd):(4'hb)]} ?
                              (^$unsigned(reg754)) : reg774) : (reg771 ?
                              ((~^reg734) * (~^forvar742)) : {(reg787 ~^ reg760)}));
                      reg798 <= reg772;
                    end
                  else
                    begin
                      reg796 <= reg748;
                      reg797 <= (($signed(reg807[(2'h3):(1'h1)]) ?
                          (forvar732[(1'h1):(1'h1)] & (forvar752 >= reg780)) : (&(8'hae))) * $unsigned(reg728[(3'h5):(3'h5)]));
                      reg798 <= $signed($signed(((!reg731) ?
                          $unsigned((8'hb8)) : reg792)));
                      reg799 <= {$unsigned($unsigned($signed(reg762)))};
                    end
                end
              for (forvar800 = (1'h0); (forvar800 < (1'h1)); forvar800 = (forvar800 + (1'h1)))
                begin
                  if ({((+reg793[(4'hb):(3'h6)]) ? (^~{reg775}) : (8'ha2))})
                    begin
                      reg801 <= (forvar735[(2'h2):(2'h2)] >= reg763);
                      reg802 <= (reg728[(1'h1):(1'h0)] + $signed(($signed(forvar794) ?
                          reg808 : forvar767[(3'h4):(2'h3)])));
                    end
                  else
                    begin
                      reg801 <= (((&$signed(reg809)) ?
                          reg744 : reg744) - reg744[(3'h7):(2'h3)]);
                      reg802 <= ((8'hb0) ?
                          (($unsigned((8'hba)) < $unsigned(reg729)) ?
                              (8'ha6) : $unsigned((forvar732 != reg775))) : (((reg806 ?
                              forvar794 : reg802) <= reg735) ^~ (forvar805 ^ $signed(reg768))));
                      reg803 <= (reg738 != {(forvar747[(3'h4):(2'h3)] * ((8'ha0) > (8'hb5)))});
                    end
                  for (forvar804 = (1'h0); (forvar804 < (2'h2)); forvar804 = (forvar804 + (1'h1)))
                    begin
                      reg805 <= reg799[(4'ha):(1'h1)];
                      reg806 <= $unsigned($unsigned(reg803));
                    end
                  reg807 <= $unsigned($signed($signed((|reg794))));
                  for (forvar808 = (1'h0); (forvar808 < (1'h0)); forvar808 = (forvar808 + (1'h1)))
                    begin
                      reg809 <= ($signed(((reg794 > reg808) ?
                              $unsigned(reg788) : reg748)) ?
                          (8'ha6) : (~&(|reg763)));
                      reg810 <= $signed($unsigned(reg772[(1'h1):(1'h0)]));
                    end
                end
            end
        end
      else
        begin
          if ((8'hb7))
            begin
              reg730 <= (reg776[(2'h3):(1'h0)] > (8'ha1));
              reg731 <= forvar778[(4'ha):(4'h9)];
            end
          else
            begin
              if ({$signed({(~^reg780)})})
                begin
                  for (forvar730 = (1'h0); (forvar730 < (1'h1)); forvar730 = (forvar730 + (1'h1)))
                    begin
                      reg731 <= $unsigned(forvar795);
                    end
                  for (forvar732 = (1'h0); (forvar732 < (2'h2)); forvar732 = (forvar732 + (1'h1)))
                    begin
                      reg733 <= $signed(reg785[(2'h2):(1'h0)]);
                      reg734 <= {$unsigned(reg756)};
                      reg735 <= reg799;
                    end
                  reg736 <= $signed((-forvar773[(1'h0):(1'h0)]));
                end
              else
                begin
                  for (forvar730 = (1'h0); (forvar730 < (1'h1)); forvar730 = (forvar730 + (1'h1)))
                    begin
                      reg731 <= $signed($unsigned((~^(forvar758 | forvar730))));
                      reg732 <= ($signed(forvar732) < wire725[(2'h2):(2'h2)]);
                      reg733 <= reg798[(3'h4):(2'h3)];
                      reg734 <= wire726[(3'h4):(2'h2)];
                    end
                  reg735 <= reg757;
                  if ((+((8'haf) ?
                      forvar747[(1'h1):(1'h0)] : $unsigned(reg755))))
                    begin
                      reg736 <= wire727[(3'h4):(2'h2)];
                      reg737 <= (~|(reg777 ^ ((~|(8'hab)) && $signed(reg802))));
                      reg738 <= reg806;
                    end
                  else
                    begin
                      reg736 <= ((-((forvar796 >> (8'ha7)) >> $unsigned(reg785))) < reg787[(3'h5):(3'h5)]);
                    end
                  for (forvar739 = (1'h0); (forvar739 < (2'h3)); forvar739 = (forvar739 + (1'h1)))
                    begin
                      reg740 <= {reg751[(2'h2):(2'h2)]};
                      reg741 <= reg793[(1'h0):(1'h0)];
                      reg742 <= (reg770[(1'h0):(1'h0)] ?
                          reg754 : reg799[(3'h4):(3'h4)]);
                    end
                end
              if (reg802[(5'h10):(3'h5)])
                begin
                  for (forvar743 = (1'h0); (forvar743 < (1'h1)); forvar743 = (forvar743 + (1'h1)))
                    begin
                      reg744 <= ($signed(reg802) == (reg743 ?
                          $signed(reg743[(3'h6):(1'h0)]) : (reg785[(3'h6):(2'h3)] ?
                              reg809 : (reg774 ^ wire725))));
                      reg745 <= ((wire725[(1'h1):(1'h0)] ?
                          reg743[(3'h7):(3'h7)] : reg765) > $signed($unsigned({reg736})));
                      reg746 <= (&reg787[(3'h7):(3'h5)]);
                    end
                  reg747 <= ($signed($signed({reg753})) ?
                      $signed($signed($signed(reg796))) : $signed(((reg773 ?
                              reg739 : reg793) ?
                          wire724[(4'hb):(3'h5)] : $unsigned(reg802))));
                end
              else
                begin
                  for (forvar743 = (1'h0); (forvar743 < (1'h0)); forvar743 = (forvar743 + (1'h1)))
                    begin
                      reg744 <= reg810[(4'h9):(4'h8)];
                    end
                end
            end
          for (forvar748 = (1'h0); (forvar748 < (1'h1)); forvar748 = (forvar748 + (1'h1)))
            begin
              if (reg786)
                begin
                  for (forvar749 = (1'h0); (forvar749 < (2'h2)); forvar749 = (forvar749 + (1'h1)))
                    begin
                      reg750 <= reg749;
                    end
                  for (forvar751 = (1'h0); (forvar751 < (1'h0)); forvar751 = (forvar751 + (1'h1)))
                    begin
                      reg752 <= $signed(reg808[(3'h6):(3'h5)]);
                      reg753 <= reg744[(3'h7):(2'h3)];
                    end
                  reg754 <= $unsigned(wire723);
                  if ($signed((((~|reg729) ?
                      (!(8'ha7)) : (forvar766 >= forvar795)) >= (8'h9e))))
                    begin
                      reg755 <= (!reg740);
                      reg756 <= $signed($unsigned(((~|(8'hb3)) < $unsigned(reg754))));
                      reg757 <= reg756;
                      reg758 <= reg748[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg755 <= $signed((($signed(reg748) ?
                              $unsigned(reg809) : $signed(reg772)) ?
                          (wire723[(1'h1):(1'h1)] ?
                              (^reg736) : (wire723 > reg807)) : $unsigned(reg759)));
                      reg756 <= ({(reg776[(1'h0):(1'h0)] ?
                                  $signed(reg765) : (reg772 - reg734))} ?
                          {forvar748} : (~$unsigned(reg754[(4'ha):(3'h7)])));
                    end
                end
              else
                begin
                  for (forvar749 = (1'h0); (forvar749 < (1'h1)); forvar749 = (forvar749 + (1'h1)))
                    begin
                      reg750 <= $unsigned((((forvar794 ? forvar759 : reg740) ?
                              $unsigned(reg793) : (forvar749 ?
                                  reg794 : reg791)) ?
                          reg763 : $unsigned((reg790 ?
                              forvar796 : forvar805))));
                      reg751 <= $unsigned(((-reg738[(4'ha):(4'ha)]) < wire724));
                      reg752 <= (($signed($signed(reg797)) ?
                              ($signed(reg735) >> reg783[(4'h8):(3'h5)]) : {(wire725 - reg732)}) ?
                          (({reg734} >> reg754[(4'hc):(2'h3)]) ?
                              ($signed(forvar735) ?
                                  (forvar808 ?
                                      reg757 : reg741) : {(8'ha8)}) : $signed((reg779 ^~ forvar751))) : $signed((^forvar767[(2'h3):(2'h2)])));
                    end
                  for (forvar753 = (1'h0); (forvar753 < (2'h3)); forvar753 = (forvar753 + (1'h1)))
                    begin
                      reg754 <= ((($signed(forvar742) ~^ $signed(forvar747)) >= (~|(|reg750))) < (!(~&forvar747[(2'h2):(1'h0)])));
                      reg755 <= ($unsigned(((reg770 >= (8'hb1)) & (reg791 ^~ (8'ha4)))) ?
                          $signed(forvar739) : ((^~reg802[(3'h4):(1'h0)]) ?
                              ($signed(reg790) ?
                                  $signed(reg748) : $unsigned(reg790)) : (reg796[(4'hb):(3'h6)] ?
                                  $signed(reg748) : $signed(forvar805))));
                      reg756 <= forvar804[(1'h0):(1'h0)];
                      reg757 <= ($signed((^$unsigned(reg808))) == ((reg737 * $signed(reg750)) != reg755));
                    end
                  if ($unsigned({reg780[(1'h1):(1'h1)]}))
                    begin
                      reg758 <= ((~|forvar752) ?
                          $unsigned($unsigned($unsigned(reg773))) : {(reg730[(4'he):(4'hb)] ?
                                  (reg749 ?
                                      reg751 : (8'ha6)) : $signed(reg736))});
                      reg759 <= (!$signed(reg747[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg758 <= (^$unsigned($unsigned(wire727[(4'h8):(1'h0)])));
                      reg759 <= (|{({reg795} ?
                              (forvar773 ? reg741 : reg729) : (^reg765))});
                    end
                end
              for (forvar760 = (1'h0); (forvar760 < (2'h2)); forvar760 = (forvar760 + (1'h1)))
                begin
                  for (forvar761 = (1'h0); (forvar761 < (2'h3)); forvar761 = (forvar761 + (1'h1)))
                    begin
                      reg762 <= forvar730[(1'h1):(1'h1)];
                      reg763 <= $signed(reg729[(4'h8):(2'h2)]);
                    end
                  for (forvar764 = (1'h0); (forvar764 < (2'h2)); forvar764 = (forvar764 + (1'h1)))
                    begin
                      reg765 <= $signed((-(reg746[(2'h2):(2'h2)] != $unsigned((8'h9e)))));
                    end
                end
            end
        end
      for (forvar811 = (1'h0); (forvar811 < (1'h0)); forvar811 = (forvar811 + (1'h1)))
        begin
          if (reg730)
            begin
              for (forvar812 = (1'h0); (forvar812 < (2'h3)); forvar812 = (forvar812 + (1'h1)))
                begin
                  reg813 <= (!($signed($signed(forvar804)) >= $signed({(8'hae)})));
                end
              if (reg793)
                begin
                  if ($unsigned((!({reg746} | forvar735))))
                    begin
                      reg814 <= reg786[(1'h1):(1'h0)];
                      reg815 <= reg809[(3'h6):(1'h0)];
                    end
                  else
                    begin
                      reg814 <= reg728[(2'h2):(1'h0)];
                    end
                  reg816 <= forvar752[(2'h3):(2'h2)];
                end
              else
                begin
                  for (forvar814 = (1'h0); (forvar814 < (1'h1)); forvar814 = (forvar814 + (1'h1)))
                    begin
                      reg815 <= $signed(((~(^~reg760)) >= ({forvar749} == (forvar747 << reg770))));
                      reg816 <= (((~&(forvar761 ?
                              forvar739 : forvar742)) & reg744[(2'h2):(1'h0)]) ?
                          {$signed({(8'hb5)})} : (forvar749 ?
                              reg783[(2'h2):(1'h0)] : reg760));
                    end
                end
              reg817 <= (((|(reg796 ?
                  wire724 : forvar758)) ^ $unsigned({reg810})) + forvar735);
            end
          else
            begin
              if ((((^(^forvar805)) ~^ {{reg786}}) >= forvar796[(2'h3):(1'h0)]))
                begin
                  reg812 <= $signed($unsigned(forvar808));
                end
              else
                begin
                  if (reg738[(4'hc):(3'h7)])
                    begin
                      reg812 <= ($unsigned($signed((~|reg732))) == (forvar778[(3'h6):(2'h2)] == (8'haa)));
                    end
                  else
                    begin
                      reg812 <= $unsigned($signed(reg786));
                      reg813 <= reg765;
                    end
                  if (forvar758)
                    begin
                      reg814 <= $signed((~|(|$signed(reg785))));
                    end
                  else
                    begin
                      reg814 <= $unsigned(($unsigned(((8'hb2) <<< reg803)) ?
                          reg798[(3'h4):(2'h2)] : reg785));
                      reg815 <= (~|(^~(8'hba)));
                      reg816 <= reg762[(3'h4):(1'h1)];
                      reg817 <= (($signed($unsigned(forvar790)) ?
                          (reg799 ?
                              {(8'h9c)} : forvar730[(1'h1):(1'h1)]) : ({reg768} << (reg749 ^~ forvar747))) <= reg729[(4'hc):(2'h3)]);
                    end
                end
              if ($signed((~forvar760[(3'h6):(3'h6)])))
                begin
                  if ($unsigned(reg815[(3'h6):(1'h0)]))
                    begin
                      reg818 <= {$signed(($unsigned(reg762) || (reg796 == reg752)))};
                      reg819 <= {(($signed(reg745) ?
                              $unsigned(reg768) : $unsigned(reg793)) > (reg739[(3'h6):(2'h3)] != reg774[(2'h3):(1'h1)]))};
                      reg820 <= (reg771 + reg781[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg818 <= $signed($signed($unsigned($unsigned(reg736))));
                      reg819 <= (|$signed($unsigned(reg790)));
                    end
                  reg821 <= (!$signed((^{reg786})));
                  if ($signed($unsigned(reg770[(1'h1):(1'h1)])))
                    begin
                      reg822 <= ($unsigned((forvar759 ?
                              (forvar749 ^ reg733) : (reg786 ^~ reg749))) ?
                          (^~reg749) : forvar804);
                      reg823 <= ({$unsigned((reg791 + forvar794))} ?
                          (reg744 ?
                              (-$unsigned(reg765)) : {(reg749 < forvar814)}) : ((~&(~reg796)) ?
                              (!(reg764 ?
                                  forvar732 : (8'hae))) : ((reg756 == wire726) ^~ reg793)));
                    end
                  else
                    begin
                      reg822 <= ((reg793[(4'hb):(4'ha)] ~^ reg819[(3'h5):(3'h4)]) >> {reg802});
                      reg823 <= $signed(($unsigned(forvar766[(4'h9):(3'h6)]) | (&reg810)));
                      reg824 <= (&$signed({$signed(reg729)}));
                      reg825 <= reg729[(1'h0):(1'h0)];
                    end
                  for (forvar826 = (1'h0); (forvar826 < (1'h0)); forvar826 = (forvar826 + (1'h1)))
                    begin
                      reg827 <= (($signed((forvar804 | reg821)) == (reg739[(1'h0):(1'h0)] ?
                              reg749 : reg814[(1'h0):(1'h0)])) ?
                          (reg741 ?
                              $signed(reg812[(4'h8):(2'h3)]) : {((8'hb4) ?
                                      reg758 : reg755)}) : reg750[(1'h0):(1'h0)]);
                      reg828 <= wire723;
                    end
                end
              else
                begin
                  if ((~$unsigned({(forvar811 ? (8'ha6) : reg791)})))
                    begin
                      reg818 <= reg802;
                      reg819 <= $signed(forvar758);
                      reg820 <= $signed({forvar804});
                      reg821 <= reg805;
                    end
                  else
                    begin
                      reg818 <= $unsigned(((~&(reg762 ?
                          (8'had) : (8'hb1))) <= (~|(reg815 ?
                          (8'hb3) : (8'ha5)))));
                      reg819 <= $unsigned(reg772[(3'h4):(3'h4)]);
                      reg820 <= (+(^~(~|reg746)));
                    end
                  for (forvar822 = (1'h0); (forvar822 < (2'h2)); forvar822 = (forvar822 + (1'h1)))
                    begin
                      reg823 <= ($unsigned(reg742[(4'hf):(4'h9)]) || ((^wire723[(1'h0):(1'h0)]) ?
                          (reg805 << (reg820 >= reg736)) : ({(8'hb3)} ?
                              {reg802} : reg798)));
                      reg824 <= ((((forvar800 ?
                              (8'hb3) : forvar795) && $signed((8'ha0))) > ($signed((8'ha0)) && {reg728})) ?
                          (&reg817[(2'h3):(1'h1)]) : ($unsigned($signed((8'ha6))) <= reg773[(1'h1):(1'h0)]));
                      reg825 <= forvar751;
                    end
                  for (forvar826 = (1'h0); (forvar826 < (2'h2)); forvar826 = (forvar826 + (1'h1)))
                    begin
                      reg827 <= reg749[(4'ha):(4'h8)];
                      reg828 <= (~&{forvar746[(4'h8):(3'h7)]});
                    end
                end
              reg829 <= {({reg824} != ((~^wire726) ?
                      (|(8'hae)) : ((8'hab) ? forvar751 : reg786)))};
            end
          if ($signed(reg809[(2'h3):(1'h0)]))
            begin
              for (forvar830 = (1'h0); (forvar830 < (2'h3)); forvar830 = (forvar830 + (1'h1)))
                begin
                  if (((^({reg799} == (forvar759 >>> (8'hb7)))) & (&({reg746} <= (reg783 ?
                      reg732 : (8'hb3))))))
                    begin
                      reg831 <= $signed($signed(((-(8'ha4)) <<< reg787[(3'h4):(1'h1)])));
                      reg832 <= $unsigned(reg765[(4'h8):(2'h2)]);
                      reg833 <= forvar767;
                      reg834 <= wire724[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg831 <= ($unsigned(reg760) != (8'hab));
                    end
                  for (forvar835 = (1'h0); (forvar835 < (1'h1)); forvar835 = (forvar835 + (1'h1)))
                    begin
                      reg836 <= ($signed((!wire725)) ?
                          $signed(((forvar732 * forvar794) >= $signed(reg781))) : $signed(($unsigned((8'hb9)) <= {reg756})));
                    end
                end
              for (forvar837 = (1'h0); (forvar837 < (2'h2)); forvar837 = (forvar837 + (1'h1)))
                begin
                  for (forvar838 = (1'h0); (forvar838 < (1'h0)); forvar838 = (forvar838 + (1'h1)))
                    begin
                      reg839 <= forvar735[(1'h0):(1'h0)];
                      reg840 <= (^~$signed($signed($signed(reg831))));
                      reg841 <= (({(8'hac)} ?
                              {(~^reg732)} : $unsigned((reg822 < (8'h9e)))) ?
                          $signed(reg735) : forvar778);
                    end
                  for (forvar842 = (1'h0); (forvar842 < (1'h0)); forvar842 = (forvar842 + (1'h1)))
                    begin
                      reg843 <= $unsigned($unsigned((!reg745)));
                      reg844 <= reg829[(3'h5):(2'h3)];
                      reg845 <= {$unsigned(reg823[(3'h4):(2'h3)])};
                      reg846 <= ((|reg829) ^ $unsigned((((8'hb4) | forvar838) ?
                          $signed(forvar830) : (reg758 >> reg772))));
                    end
                end
            end
          else
            begin
              reg830 <= ($unsigned((reg821 != ((8'hb0) ? reg841 : reg798))) ?
                  (~$unsigned($signed(reg821))) : $signed(reg820));
              if ((8'hb1))
                begin
                  for (forvar831 = (1'h0); (forvar831 < (2'h3)); forvar831 = (forvar831 + (1'h1)))
                    begin
                      reg832 <= (8'hb5);
                      reg833 <= ($signed(reg762) ?
                          ({$unsigned((8'hb1))} ?
                              forvar794[(2'h3):(1'h0)] : (reg825[(4'ha):(3'h6)] ?
                                  forvar761 : reg765)) : (((8'ha5) ?
                              reg738[(4'hf):(1'h1)] : (wire723 ?
                                  (8'hb0) : reg751)) <= $unsigned($signed(reg772))));
                      reg834 <= $signed(((-reg791[(3'h5):(2'h2)]) - $signed({forvar766})));
                    end
                end
              else
                begin
                  if ($signed(reg795[(1'h0):(1'h0)]))
                    begin
                      reg831 <= $unsigned({reg815});
                    end
                  else
                    begin
                      reg831 <= ((!{(reg769 ? (8'hb8) : reg771)}) || reg738);
                      reg832 <= forvar842[(3'h6):(3'h4)];
                      reg833 <= $signed(reg772[(3'h5):(2'h3)]);
                    end
                  for (forvar834 = (1'h0); (forvar834 < (1'h0)); forvar834 = (forvar834 + (1'h1)))
                    begin
                      reg835 <= reg783[(3'h7):(2'h2)];
                    end
                end
              for (forvar836 = (1'h0); (forvar836 < (1'h1)); forvar836 = (forvar836 + (1'h1)))
                begin
                  if (reg753)
                    begin
                      reg837 <= $signed(({forvar739[(2'h3):(1'h0)]} ^ ($unsigned(reg750) ?
                          $signed((8'haa)) : forvar742)));
                    end
                  else
                    begin
                      reg837 <= $signed($unsigned($signed(((8'hb6) ?
                          forvar773 : (8'hb1)))));
                      reg838 <= ($unsigned(forvar794[(2'h3):(2'h2)]) - reg746[(3'h4):(1'h0)]);
                      reg839 <= ((($unsigned(forvar730) < (-forvar837)) ?
                              ({reg831} & (reg756 << (8'haa))) : (8'ha8)) ?
                          $signed(reg747[(2'h3):(1'h0)]) : {reg739});
                    end
                  for (forvar840 = (1'h0); (forvar840 < (2'h3)); forvar840 = (forvar840 + (1'h1)))
                    begin
                      reg841 <= (|($unsigned(((8'haf) ? reg754 : reg770)) ?
                          ({forvar812} || {reg796}) : (forvar752 ?
                              (reg738 ?
                                  reg756 : (8'ha6)) : reg753[(3'h6):(3'h5)])));
                    end
                end
            end
          for (forvar847 = (1'h0); (forvar847 < (2'h3)); forvar847 = (forvar847 + (1'h1)))
            begin
              if ((~^(~reg793)))
                begin
                  for (forvar848 = (1'h0); (forvar848 < (2'h3)); forvar848 = (forvar848 + (1'h1)))
                    begin
                      reg849 <= reg829[(3'h4):(1'h1)];
                      reg850 <= {(($unsigned(reg835) ?
                              (8'haf) : $unsigned(reg768)) ^ reg732[(4'hc):(1'h0)])};
                      reg851 <= (^~reg764);
                      reg852 <= (~reg812);
                    end
                  if (reg769)
                    begin
                      reg853 <= $unsigned((!forvar764));
                      reg854 <= {(-((!(8'ha4)) ?
                              (forvar778 > reg790) : wire727[(4'h9):(1'h1)]))};
                    end
                  else
                    begin
                      reg853 <= (($signed((~^reg734)) ?
                          ($unsigned((8'hb2)) ?
                              (forvar759 >> (8'ha9)) : (|forvar748)) : ({(8'hb1)} && $signed(forvar842))) && {forvar830});
                      reg854 <= (reg827[(4'h8):(3'h6)] < forvar835);
                      reg855 <= reg794[(1'h1):(1'h0)];
                      reg856 <= (|(!(|reg810[(1'h1):(1'h1)])));
                    end
                end
              else
                begin
                  if ($unsigned(reg833))
                    begin
                      reg848 <= $unsigned(($signed(reg770[(2'h3):(2'h2)]) ?
                          $signed(((8'ha4) ?
                              (8'hab) : (8'had))) : (^~(~reg751))));
                      reg849 <= $unsigned($unsigned(reg751[(3'h6):(3'h4)]));
                      reg850 <= reg773;
                    end
                  else
                    begin
                      reg848 <= (reg753[(3'h6):(2'h3)] + (-(reg805[(2'h2):(1'h1)] ?
                          (reg831 ?
                              forvar847 : forvar840) : (reg831 ^~ forvar795))));
                      reg849 <= reg797[(4'h8):(2'h3)];
                    end
                end
              for (forvar857 = (1'h0); (forvar857 < (2'h2)); forvar857 = (forvar857 + (1'h1)))
                begin
                  for (forvar858 = (1'h0); (forvar858 < (2'h2)); forvar858 = (forvar858 + (1'h1)))
                    begin
                      reg859 <= $signed((((forvar808 * reg788) ?
                          {forvar842} : {reg836}) || wire727));
                      reg860 <= ($signed((forvar773[(2'h3):(1'h1)] ?
                          reg854 : ((8'hac) ^ reg821))) || forvar746);
                      reg861 <= (($unsigned({reg757}) ~^ $unsigned(forvar808[(1'h0):(1'h0)])) * $unsigned($signed((8'ha7))));
                    end
                  for (forvar862 = (1'h0); (forvar862 < (1'h1)); forvar862 = (forvar862 + (1'h1)))
                    begin
                      reg863 <= $signed((((forvar826 ?
                          reg787 : (8'ha9)) - (~&reg737)) && (reg836 <<< $signed(reg833))));
                      reg864 <= {{$signed((~reg788))}};
                      reg865 <= ({$unsigned($signed((8'ha7)))} >>> $signed(forvar746[(2'h3):(2'h3)]));
                    end
                end
              reg866 <= ($signed((~&(~&wire725))) | ({reg797} - {$signed((8'hac))}));
            end
        end
    end
  module867 #() modinst2032 (.wire868(reg820), .wire871(reg832), .wire869(reg849), .y(wire2031), .clk(clk), .wire870(reg765));
  assign wire2033 = $unsigned(reg799[(1'h0):(1'h0)]);
  module2034 #() modinst3426 (.wire2038(reg822), .wire2035(reg785), .clk(clk), .wire2036(reg853), .y(wire3425), .wire2037(reg773));
  always
    @(posedge clk) begin
      for (forvar3427 = (1'h0); (forvar3427 < (2'h2)); forvar3427 = (forvar3427 + (1'h1)))
        begin
          for (forvar3428 = (1'h0); (forvar3428 < (2'h3)); forvar3428 = (forvar3428 + (1'h1)))
            begin
              if (reg846)
                begin
                  if ($signed($signed(($unsigned(reg731) ?
                      ((8'hae) ? reg743 : reg788) : reg853))))
                    begin
                      reg3429 <= $signed((~|{reg791}));
                      reg3430 <= $signed(reg753);
                    end
                  else
                    begin
                      reg3429 <= reg849[(3'h7):(2'h3)];
                      reg3430 <= ((((~|(8'hba)) ?
                                  (~^reg741) : (reg796 <<< reg784)) ?
                              (reg761[(3'h7):(3'h4)] ?
                                  (8'h9f) : reg770) : reg852) ?
                          $unsigned((8'haa)) : ((|reg741) && $signed($unsigned(reg839))));
                      reg3431 <= reg805[(3'h6):(2'h2)];
                      reg3432 <= reg844[(3'h5):(1'h1)];
                    end
                  if ((($signed(reg822) ?
                          ((reg742 && reg807) * (reg735 ?
                              reg758 : reg784)) : reg733) ?
                      ($signed((reg787 | reg807)) ?
                          reg805[(1'h0):(1'h0)] : (-(8'hb3))) : ((~|(reg797 ?
                          reg827 : reg854)) >>> (~|(reg796 <= reg787)))))
                    begin
                      reg3433 <= $unsigned($signed($signed($signed(reg819))));
                    end
                  else
                    begin
                      reg3433 <= (~|$signed($signed(reg757)));
                      reg3434 <= ((^~$signed($unsigned(reg853))) ?
                          {((reg820 & reg728) ?
                                  (reg799 ?
                                      reg752 : reg770) : reg833)} : reg808[(4'hc):(2'h3)]);
                      reg3435 <= reg853;
                    end
                  if (reg806[(2'h2):(2'h2)])
                    begin
                      reg3436 <= ($unsigned($unsigned({reg757})) ?
                          reg866[(2'h2):(2'h2)] : $signed($unsigned($unsigned((8'ha1)))));
                      reg3437 <= reg764;
                      reg3438 <= (&reg859[(4'ha):(1'h0)]);
                      reg3439 <= ($signed(((~reg837) ?
                              ((8'hb3) || reg775) : reg863)) ?
                          reg790[(4'hf):(3'h7)] : $signed(reg780));
                    end
                  else
                    begin
                      reg3436 <= $signed($unsigned((~reg853)));
                      reg3437 <= $unsigned($unsigned(reg802[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  reg3429 <= reg820;
                end
              for (forvar3440 = (1'h0); (forvar3440 < (2'h3)); forvar3440 = (forvar3440 + (1'h1)))
                begin
                  for (forvar3441 = (1'h0); (forvar3441 < (1'h1)); forvar3441 = (forvar3441 + (1'h1)))
                    begin
                      reg3442 <= reg856[(3'h4):(2'h3)];
                    end
                  reg3443 <= $signed((((reg809 ? reg866 : (8'hb2)) ?
                      {forvar3427} : reg810[(3'h5):(1'h0)]) | ({reg821} << (~|(8'hb6)))));
                  reg3444 <= {$unsigned(reg831[(1'h1):(1'h1)])};
                end
            end
          reg3445 <= ((reg802[(1'h1):(1'h1)] && (~$unsigned(reg775))) >>> $signed(($signed(reg741) < reg787)));
        end
      if (($unsigned($unsigned($signed((8'ha9)))) <<< $unsigned(($signed(reg859) ?
          ((8'ha8) >>> reg742) : (~reg809)))))
        begin
          for (forvar3446 = (1'h0); (forvar3446 < (1'h0)); forvar3446 = (forvar3446 + (1'h1)))
            begin
              if ((^(reg787 ?
                  ((&reg863) >>> (reg732 < reg809)) : $unsigned({(8'ha9)}))))
                begin
                  for (forvar3447 = (1'h0); (forvar3447 < (2'h3)); forvar3447 = (forvar3447 + (1'h1)))
                    begin
                      reg3448 <= $signed((&(forvar3427[(2'h2):(1'h1)] ?
                          forvar3446 : (reg756 ? reg864 : (8'h9f)))));
                      reg3449 <= reg843[(1'h1):(1'h1)];
                      reg3450 <= reg786;
                    end
                end
              else
                begin
                  for (forvar3447 = (1'h0); (forvar3447 < (2'h3)); forvar3447 = (forvar3447 + (1'h1)))
                    begin
                      reg3448 <= reg822[(4'ha):(3'h6)];
                      reg3449 <= ((reg856 ? $unsigned(reg3430) : reg781) ?
                          (-(8'h9e)) : ((8'had) ?
                              (forvar3427[(1'h1):(1'h1)] ?
                                  $unsigned(reg3437) : (8'ha4)) : reg851[(3'h5):(3'h5)]));
                      reg3450 <= reg834;
                      reg3451 <= $unsigned(reg3429[(3'h5):(2'h3)]);
                    end
                  for (forvar3452 = (1'h0); (forvar3452 < (1'h0)); forvar3452 = (forvar3452 + (1'h1)))
                    begin
                      reg3453 <= reg796;
                      reg3454 <= ((~|(forvar3427 ?
                          $signed((8'ha1)) : $signed(reg794))) < ((^~(reg777 > reg3451)) ?
                          reg772[(1'h1):(1'h1)] : (wire2033[(1'h1):(1'h1)] ?
                              $signed((8'hb4)) : (reg817 + reg785))));
                      reg3455 <= $signed($signed(reg3449));
                    end
                end
              for (forvar3456 = (1'h0); (forvar3456 < (1'h1)); forvar3456 = (forvar3456 + (1'h1)))
                begin
                  reg3457 <= (~&reg737[(3'h5):(1'h1)]);
                  for (forvar3458 = (1'h0); (forvar3458 < (1'h0)); forvar3458 = (forvar3458 + (1'h1)))
                    begin
                      reg3459 <= reg3429[(3'h7):(2'h2)];
                      reg3460 <= (8'hb7);
                    end
                  for (forvar3461 = (1'h0); (forvar3461 < (1'h1)); forvar3461 = (forvar3461 + (1'h1)))
                    begin
                      reg3462 <= $unsigned(reg764);
                      reg3463 <= reg735;
                    end
                end
            end
        end
      else
        begin
          if ($signed((~(~&reg763[(3'h5):(3'h4)]))))
            begin
              for (forvar3446 = (1'h0); (forvar3446 < (2'h2)); forvar3446 = (forvar3446 + (1'h1)))
                begin
                  for (forvar3447 = (1'h0); (forvar3447 < (2'h2)); forvar3447 = (forvar3447 + (1'h1)))
                    begin
                      reg3448 <= wire724;
                      reg3449 <= ({(reg3459[(1'h1):(1'h1)] == (reg839 > reg777))} ?
                          (reg806 & (-$signed(reg3439))) : $unsigned($unsigned((&reg732))));
                    end
                end
              if ($signed((($signed(reg752) + (&forvar3447)) ?
                  ((reg774 | reg3463) ?
                      (reg853 ? reg820 : (8'h9f)) : (^reg757)) : reg779)))
                begin
                  for (forvar3450 = (1'h0); (forvar3450 < (1'h1)); forvar3450 = (forvar3450 + (1'h1)))
                    begin
                      reg3451 <= $unsigned(reg799[(1'h0):(1'h0)]);
                      reg3452 <= reg751[(3'h6):(2'h2)];
                      reg3453 <= (~&$unsigned({{(8'h9e)}}));
                      reg3454 <= $signed($unsigned(reg765));
                    end
                  reg3455 <= reg861;
                  for (forvar3456 = (1'h0); (forvar3456 < (2'h3)); forvar3456 = (forvar3456 + (1'h1)))
                    begin
                      reg3457 <= ($unsigned((((8'hb9) ?
                              reg3435 : reg791) <= (reg755 ?
                              reg813 : (8'ha7)))) ?
                          reg3429 : (-$unsigned($unsigned(reg782))));
                    end
                end
              else
                begin
                  for (forvar3450 = (1'h0); (forvar3450 < (1'h0)); forvar3450 = (forvar3450 + (1'h1)))
                    begin
                      reg3451 <= reg739[(3'h7):(3'h7)];
                    end
                  reg3452 <= reg743[(3'h4):(2'h3)];
                  for (forvar3453 = (1'h0); (forvar3453 < (1'h1)); forvar3453 = (forvar3453 + (1'h1)))
                    begin
                      reg3454 <= $unsigned({wire724});
                      reg3455 <= $unsigned((~&((forvar3428 ?
                          reg760 : reg760) >>> (reg852 ^ reg3443))));
                      reg3456 <= $unsigned(($unsigned({reg850}) >> (~|(reg852 || reg781))));
                    end
                end
              if (reg728[(2'h3):(2'h2)])
                begin
                  for (forvar3458 = (1'h0); (forvar3458 < (1'h0)); forvar3458 = (forvar3458 + (1'h1)))
                    begin
                      reg3459 <= ((~^(~|forvar3427[(1'h0):(1'h0)])) || reg3450[(4'h8):(4'h8)]);
                    end
                end
              else
                begin
                  for (forvar3458 = (1'h0); (forvar3458 < (2'h2)); forvar3458 = (forvar3458 + (1'h1)))
                    begin
                      reg3459 <= reg805[(2'h3):(1'h0)];
                      reg3460 <= (8'h9d);
                      reg3461 <= ((({reg796} ?
                              (reg850 ? (8'hab) : reg3452) : (^~(8'had))) ?
                          $signed($signed(reg737)) : (reg3450[(4'h8):(3'h4)] > $unsigned(reg821))) && reg3432[(3'h7):(3'h7)]);
                      reg3462 <= $signed($signed({(~^reg834)}));
                    end
                  if (($signed({$signed((8'hb1))}) ?
                      $unsigned((reg3453[(4'h8):(3'h4)] != $unsigned(reg3450))) : wire3425))
                    begin
                      reg3463 <= $unsigned({($signed(reg791) ?
                              $unsigned((8'ha3)) : reg800[(2'h3):(2'h3)])});
                      reg3464 <= $unsigned(reg850);
                      reg3465 <= $unsigned((($unsigned(reg865) >= reg830[(2'h3):(1'h1)]) > (|$signed(reg861))));
                      reg3466 <= (($unsigned(reg823) - (8'h9e)) < reg3450[(3'h7):(3'h7)]);
                    end
                  else
                    begin
                      reg3463 <= $signed(($unsigned((-reg850)) ?
                          wire2033[(3'h6):(2'h2)] : $signed(reg820)));
                    end
                  for (forvar3467 = (1'h0); (forvar3467 < (2'h3)); forvar3467 = (forvar3467 + (1'h1)))
                    begin
                      reg3468 <= reg828[(4'h8):(3'h7)];
                      reg3469 <= (reg783[(1'h0):(1'h0)] >> reg735[(3'h6):(3'h4)]);
                      reg3470 <= (~&$unsigned($signed(reg3435[(2'h2):(1'h0)])));
                    end
                end
              for (forvar3471 = (1'h0); (forvar3471 < (2'h3)); forvar3471 = (forvar3471 + (1'h1)))
                begin
                  if (reg3455)
                    begin
                      reg3472 <= $unsigned((reg757[(2'h3):(1'h0)] ~^ {{reg749}}));
                    end
                  else
                    begin
                      reg3472 <= (reg865[(3'h4):(2'h2)] ?
                          reg753[(3'h4):(1'h0)] : ($unsigned((reg838 - reg801)) ?
                              {$unsigned(reg771)} : (8'hb2)));
                      reg3473 <= $unsigned(reg3469[(2'h2):(1'h1)]);
                    end
                end
            end
          else
            begin
              if ((~({$unsigned(reg828)} ?
                  $signed(reg832) : $unsigned((reg859 ? reg840 : reg861)))))
                begin
                  for (forvar3446 = (1'h0); (forvar3446 < (2'h2)); forvar3446 = (forvar3446 + (1'h1)))
                    begin
                      reg3447 <= reg831[(2'h3):(2'h2)];
                      reg3448 <= $unsigned((^reg733[(2'h3):(2'h2)]));
                    end
                  for (forvar3449 = (1'h0); (forvar3449 < (1'h0)); forvar3449 = (forvar3449 + (1'h1)))
                    begin
                      reg3450 <= reg3462;
                      reg3451 <= reg843[(3'h4):(2'h3)];
                      reg3452 <= forvar3456[(1'h0):(1'h0)];
                    end
                  if ($unsigned((reg731 ?
                      wire726 : $unsigned((reg765 ? reg757 : reg837)))))
                    begin
                      reg3453 <= (^~reg3466[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg3453 <= $signed({$signed((reg764 && (8'h9f)))});
                      reg3454 <= $signed(((8'ha5) ?
                          (wire2033 && reg740) : ((reg768 ?
                                  (8'hb6) : wire2031) ?
                              $unsigned(forvar3450) : $unsigned((8'hb3)))));
                    end
                  reg3455 <= (8'h9c);
                end
              else
                begin
                  for (forvar3446 = (1'h0); (forvar3446 < (2'h3)); forvar3446 = (forvar3446 + (1'h1)))
                    begin
                      reg3447 <= (|forvar3446);
                    end
                end
              for (forvar3456 = (1'h0); (forvar3456 < (1'h1)); forvar3456 = (forvar3456 + (1'h1)))
                begin
                  if ($signed(reg3462))
                    begin
                      reg3457 <= (((reg3452[(4'hb):(2'h2)] << (~|reg865)) ?
                          (8'ha1) : reg729[(3'h5):(2'h2)]) ^~ (~^reg790));
                      reg3458 <= $signed(($unsigned({reg850}) ?
                          ((8'haa) ?
                              ((8'hac) <<< (8'hb7)) : {reg740}) : $unsigned((!forvar3458))));
                    end
                  else
                    begin
                      reg3457 <= (8'ha5);
                      reg3458 <= (~|(reg748 <<< (-reg796)));
                      reg3459 <= $signed(((8'hb3) ~^ ((~&reg827) ^ (+reg3473))));
                      reg3460 <= (($signed($unsigned(reg3452)) ^ reg823[(3'h5):(3'h4)]) ?
                          $unsigned((~&$signed(reg772))) : reg733);
                    end
                end
              if (((8'ha1) ?
                  $unsigned($signed($unsigned((8'hb6)))) : $signed($unsigned(reg742[(4'hf):(4'ha)]))))
                begin
                  if ($signed((reg846[(3'h4):(2'h2)] >>> reg3447[(4'ha):(2'h3)])))
                    begin
                      reg3461 <= reg841;
                      reg3462 <= (reg836[(1'h0):(1'h0)] ?
                          (!reg729) : $unsigned((!(reg752 ? reg743 : reg846))));
                      reg3463 <= ((^{$unsigned(reg3451)}) < $unsigned((!$unsigned(reg854))));
                    end
                  else
                    begin
                      reg3461 <= ($unsigned(forvar3461[(2'h3):(2'h3)]) >> reg3450[(4'hc):(4'h8)]);
                      reg3462 <= (~|{(reg820[(2'h2):(1'h1)] * (reg837 || reg773))});
                    end
                  reg3464 <= (~^$unsigned(reg852[(3'h5):(3'h4)]));
                  for (forvar3465 = (1'h0); (forvar3465 < (1'h1)); forvar3465 = (forvar3465 + (1'h1)))
                    begin
                      reg3466 <= reg736;
                      reg3467 <= $signed(forvar3446[(3'h5):(1'h0)]);
                    end
                  for (forvar3468 = (1'h0); (forvar3468 < (1'h1)); forvar3468 = (forvar3468 + (1'h1)))
                    begin
                      reg3469 <= $unsigned($unsigned((forvar3447 ?
                          reg854 : (+reg859))));
                      reg3470 <= ({(|((8'hb2) ? reg792 : reg838))} ?
                          reg822 : (((~|reg733) + (&reg793)) > (reg3437[(3'h4):(1'h0)] ?
                              $signed(forvar3458) : reg793)));
                      reg3471 <= ((^reg3466[(1'h0):(1'h0)]) ?
                          (reg779[(3'h7):(1'h0)] << reg737[(3'h7):(3'h6)]) : $unsigned(reg814));
                      reg3472 <= ((forvar3450 ?
                          reg840 : $signed($signed(reg3431))) >= reg838);
                    end
                end
              else
                begin
                  for (forvar3461 = (1'h0); (forvar3461 < (2'h3)); forvar3461 = (forvar3461 + (1'h1)))
                    begin
                      reg3462 <= {reg3436};
                      reg3463 <= ({reg752} < $signed(({reg848} - $signed(reg753))));
                    end
                  for (forvar3464 = (1'h0); (forvar3464 < (2'h3)); forvar3464 = (forvar3464 + (1'h1)))
                    begin
                      reg3465 <= $signed($signed($signed((^~reg821))));
                      reg3466 <= $unsigned($signed($unsigned(reg832[(3'h4):(1'h1)])));
                      reg3467 <= (reg3465 ?
                          (reg3466[(1'h0):(1'h0)] && (!reg846)) : (($unsigned(forvar3452) >>> (reg835 << reg3430)) == (reg3439[(3'h7):(3'h7)] ?
                              (reg753 >> reg790) : {reg808})));
                      reg3468 <= reg741[(3'h5):(1'h1)];
                    end
                end
              reg3473 <= ($unsigned($unsigned((&(8'haa)))) << {(reg3432 ?
                      reg3451[(3'h7):(3'h5)] : $unsigned((8'ha5)))});
            end
          reg3474 <= $signed(reg749);
          for (forvar3475 = (1'h0); (forvar3475 < (2'h3)); forvar3475 = (forvar3475 + (1'h1)))
            begin
              if ((($signed($signed(reg747)) ?
                  (reg781[(1'h0):(1'h0)] >>> (wire727 || reg772)) : (reg866[(1'h0):(1'h0)] <<< $signed(reg806))) >= reg806[(3'h5):(2'h2)]))
                begin
                  for (forvar3476 = (1'h0); (forvar3476 < (2'h3)); forvar3476 = (forvar3476 + (1'h1)))
                    begin
                      reg3477 <= $signed(($signed($signed(reg3444)) ?
                          $unsigned(reg812[(3'h5):(1'h1)]) : reg824[(3'h4):(2'h2)]));
                      reg3478 <= ((((8'h9f) ?
                              ((8'hb1) ?
                                  reg824 : reg734) : reg860[(3'h5):(3'h5)]) <= (~&reg3455[(4'he):(2'h2)])) ?
                          (reg807 ~^ $signed($signed(forvar3471))) : reg746[(3'h5):(1'h0)]);
                      reg3479 <= ((((reg3473 + reg855) ?
                              $unsigned(reg3454) : reg802) <<< ($signed(reg753) ?
                              $unsigned(reg810) : $signed(reg797))) ?
                          forvar3449[(2'h3):(2'h2)] : ((((8'hb4) < reg849) << (|(8'ha1))) >> forvar3467[(3'h5):(3'h4)]));
                    end
                  reg3480 <= (reg761[(2'h3):(1'h1)] | reg812);
                  reg3481 <= reg843;
                  for (forvar3482 = (1'h0); (forvar3482 < (1'h1)); forvar3482 = (forvar3482 + (1'h1)))
                    begin
                      reg3483 <= ((($unsigned(reg3471) > reg3451) >>> (~&reg741)) | reg855[(2'h3):(2'h3)]);
                      reg3484 <= $signed($unsigned($signed($signed(reg835))));
                      reg3485 <= (8'ha0);
                    end
                end
              else
                begin
                  if ((~((~{reg856}) ? reg806 : reg728)))
                    begin
                      reg3476 <= $unsigned($signed(reg802[(2'h2):(2'h2)]));
                      reg3477 <= reg769[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg3476 <= reg782[(4'h9):(2'h3)];
                      reg3477 <= ((8'h9e) ?
                          (~^{(reg819 > (8'ha9))}) : (!$unsigned((&reg792))));
                      reg3478 <= $unsigned((reg846[(1'h1):(1'h1)] * $unsigned($signed(reg776))));
                      reg3479 <= {($signed((!forvar3453)) ?
                              {reg3454[(3'h5):(3'h5)]} : ((~reg775) ?
                                  (forvar3446 ?
                                      (8'hb0) : (8'ha2)) : (reg3429 > reg3433)))};
                    end
                  reg3480 <= reg3474;
                  reg3481 <= forvar3464;
                  reg3482 <= ($signed((~&$unsigned((8'hb4)))) ?
                      $unsigned({{reg769}}) : (wire724[(4'hf):(4'hd)] ?
                          $signed($signed(reg794)) : (reg3448 && (8'h9d))));
                end
              if (reg827)
                begin
                  if (((~|reg764[(3'h6):(3'h4)]) ?
                      reg848[(3'h7):(3'h5)] : reg758[(2'h2):(2'h2)]))
                    begin
                      reg3486 <= {$unsigned(($unsigned((8'ha5)) ?
                              ((8'hb1) ? reg756 : reg771) : (|reg783)))};
                    end
                  else
                    begin
                      reg3486 <= $signed((~|$unsigned((reg864 <<< reg3478))));
                      reg3487 <= (|$unsigned($signed((reg830 | reg3466))));
                      reg3488 <= ($unsigned(wire725) ?
                          reg777 : reg780[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar3486 = (1'h0); (forvar3486 < (2'h3)); forvar3486 = (forvar3486 + (1'h1)))
                    begin
                      reg3487 <= (8'ha3);
                      reg3488 <= ((^~(^(+reg815))) ?
                          ($signed((forvar3446 - (8'hae))) ?
                              $signed($signed((8'ha3))) : reg3461[(2'h2):(1'h1)]) : $signed($signed($unsigned(reg832))));
                      reg3489 <= $signed($signed($signed($unsigned(reg814))));
                      reg3490 <= ((reg829 ?
                          {reg762} : reg3457[(4'hf):(4'ha)]) * (8'hb3));
                    end
                  if (reg832)
                    begin
                      reg3491 <= {(~^($signed(reg853) ?
                              reg817[(1'h0):(1'h0)] : $unsigned(reg784)))};
                      reg3492 <= reg848;
                      reg3493 <= (reg741[(3'h5):(3'h5)] ?
                          $signed($signed((reg754 ?
                              reg856 : reg812))) : reg798[(2'h2):(1'h0)]);
                      reg3494 <= reg731[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg3491 <= {reg825[(4'h9):(1'h0)]};
                      reg3492 <= (((8'h9e) || $unsigned({reg3436})) ?
                          (^~{reg3437[(3'h5):(3'h4)]}) : (($unsigned(forvar3482) >>> (reg747 ?
                                  reg846 : reg3478)) ?
                              reg757[(4'hc):(4'hb)] : reg814));
                      reg3493 <= reg3486[(4'ha):(4'ha)];
                    end
                end
              for (forvar3495 = (1'h0); (forvar3495 < (2'h2)); forvar3495 = (forvar3495 + (1'h1)))
                begin
                  for (forvar3496 = (1'h0); (forvar3496 < (1'h0)); forvar3496 = (forvar3496 + (1'h1)))
                    begin
                      reg3497 <= $signed((!$signed({reg3471})));
                      reg3498 <= $signed(reg3432[(4'h8):(3'h6)]);
                      reg3499 <= (8'hba);
                      reg3500 <= (~&(8'ha7));
                    end
                  if (reg812[(3'h7):(2'h2)])
                    begin
                      reg3501 <= ((^~reg3497) + $signed(reg773));
                      reg3502 <= $unsigned(($signed((reg3486 * reg846)) ?
                          (!$unsigned(reg822)) : reg3457[(4'h8):(3'h5)]));
                      reg3503 <= (~{(((8'h9f) ~^ reg836) < (reg3453 * reg810))});
                    end
                  else
                    begin
                      reg3501 <= reg735;
                      reg3502 <= (~&((((8'ha3) ^ (8'h9e)) != (reg3478 & reg763)) ?
                          (8'hb2) : (reg3453 ?
                              (reg3456 <= reg742) : (reg779 >> (8'hb7)))));
                      reg3503 <= (^~((&reg3481) ? reg3467 : $unsigned(reg787)));
                    end
                end
              if (reg3456)
                begin
                  if ({(8'hb6)})
                    begin
                      reg3504 <= ((^~reg843[(2'h3):(2'h3)]) >>> ((^~(reg799 ^~ reg3443)) ?
                          ((reg812 ? reg3457 : reg791) ?
                              $signed(forvar3464) : $signed(reg813)) : {$signed(reg822)}));
                      reg3505 <= reg852;
                      reg3506 <= $unsigned((^~$unsigned($unsigned((8'hb9)))));
                    end
                  else
                    begin
                      reg3504 <= reg3490[(2'h2):(2'h2)];
                      reg3505 <= reg801[(1'h1):(1'h1)];
                      reg3506 <= reg3447;
                    end
                end
              else
                begin
                  if ({(&$unsigned($signed(reg3453)))})
                    begin
                      reg3504 <= (reg779[(3'h6):(1'h1)] ?
                          reg834 : $unsigned($unsigned((reg824 ?
                              reg3498 : wire724))));
                    end
                  else
                    begin
                      reg3504 <= (($unsigned((reg785 ? reg731 : (8'ha9))) ?
                              {reg735[(1'h1):(1'h1)]} : reg3473) ?
                          reg798 : ($signed((&reg771)) ^ reg748));
                    end
                  if ($signed(($signed((~|reg865)) ^ reg798)))
                    begin
                      reg3505 <= ($unsigned((-reg838)) ?
                          (8'h9c) : $signed(reg3478));
                      reg3506 <= (!(reg777 ? (8'ha7) : reg3481[(3'h6):(2'h3)]));
                    end
                  else
                    begin
                      reg3505 <= reg779;
                    end
                  if ($unsigned($signed((+reg743))))
                    begin
                      reg3507 <= wire724;
                    end
                  else
                    begin
                      reg3507 <= (reg3479[(2'h3):(2'h3)] ?
                          (reg742[(3'h5):(3'h4)] >= $signed(reg730)) : $signed({(!reg865)}));
                      reg3508 <= $unsigned({(~^(reg3481 ? reg3466 : (8'hb1)))});
                      reg3509 <= $unsigned($unsigned(($signed(reg3504) & reg3492[(3'h7):(3'h6)])));
                    end
                  if ((!(($unsigned((8'hab)) ?
                          reg828[(4'hb):(1'h1)] : (!reg833)) ?
                      reg832 : (8'hb0))))
                    begin
                      reg3510 <= ($signed($signed(reg807)) << reg3434);
                      reg3511 <= wire2031;
                    end
                  else
                    begin
                      reg3510 <= {(forvar3441 == forvar3449[(1'h0):(1'h0)])};
                      reg3511 <= (~&(reg3486[(4'hc):(4'ha)] ?
                          (|$signed(forvar3440)) : reg3497));
                    end
                end
            end
          if (((8'hb9) ?
              $unsigned(reg3449[(4'hc):(3'h6)]) : (+reg776[(1'h1):(1'h0)])))
            begin
              reg3512 <= (&(reg829 ?
                  (reg758[(1'h0):(1'h0)] << reg3444) : ($unsigned(reg3456) ^ $unsigned(reg837))));
              if ((!(((reg3452 ? reg738 : reg783) ?
                      (reg3436 < reg3438) : (reg813 < reg3498)) ?
                  (8'ha6) : $unsigned({(8'h9e)}))))
                begin
                  if (reg3474[(2'h3):(2'h3)])
                    begin
                      reg3513 <= {(($signed(reg3438) ?
                              $signed(forvar3452) : $unsigned((8'h9d))) + $signed((^reg844)))};
                      reg3514 <= (({reg3457} ?
                          $unsigned((!forvar3465)) : reg3438[(3'h6):(3'h4)]) > {reg3513});
                      reg3515 <= $unsigned((~|((^reg786) ^ reg737[(1'h1):(1'h0)])));
                      reg3516 <= ($unsigned(({reg784} && reg759)) ?
                          reg808 : reg3451);
                    end
                  else
                    begin
                      reg3513 <= {$unsigned(($unsigned((8'haf)) ^~ (~reg3429)))};
                      reg3514 <= ((((+reg776) ?
                                  ((8'hb6) ? reg3500 : reg3498) : reg763) ?
                              (((8'hb0) | (8'h9c)) << (reg3487 <<< reg819)) : ((reg819 * reg776) ?
                                  $unsigned(forvar3452) : reg3501[(1'h1):(1'h0)])) ?
                          {($unsigned(reg850) ^~ $signed(reg763))} : (|reg863[(2'h2):(2'h2)]));
                    end
                end
              else
                begin
                  for (forvar3513 = (1'h0); (forvar3513 < (1'h1)); forvar3513 = (forvar3513 + (1'h1)))
                    begin
                      reg3514 <= reg3457[(4'he):(3'h7)];
                      reg3515 <= (reg3458[(4'h8):(3'h4)] ? reg860 : reg818);
                      reg3516 <= $unsigned($signed((reg819[(1'h1):(1'h0)] ?
                          $unsigned(reg764) : wire726[(2'h2):(2'h2)])));
                    end
                end
              for (forvar3517 = (1'h0); (forvar3517 < (2'h2)); forvar3517 = (forvar3517 + (1'h1)))
                begin
                  if ((~$signed(reg3483)))
                    begin
                      reg3518 <= (((|{forvar3447}) != reg3436) * (($signed(reg743) ?
                              reg3473 : $signed(reg763)) ?
                          reg794 : $unsigned(reg759)));
                      reg3519 <= ($unsigned($unsigned($unsigned(reg802))) && {(-(reg777 ?
                              wire2033 : forvar3452))});
                      reg3520 <= ((wire725[(1'h0):(1'h0)] <= $unsigned((&wire3425))) <<< reg855[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg3518 <= ({reg791[(2'h2):(1'h0)]} ?
                          $unsigned($unsigned($unsigned(reg734))) : (^~(reg757[(3'h6):(2'h2)] - $signed(reg790))));
                      reg3519 <= reg3445[(2'h3):(1'h0)];
                      reg3520 <= reg795[(2'h2):(2'h2)];
                      reg3521 <= $unsigned(({((8'ha0) ^~ forvar3461)} & $unsigned($unsigned(forvar3486))));
                    end
                  for (forvar3522 = (1'h0); (forvar3522 < (2'h3)); forvar3522 = (forvar3522 + (1'h1)))
                    begin
                      reg3523 <= (~|{reg761[(3'h6):(3'h5)]});
                      reg3524 <= ($signed(($signed(reg806) ?
                          (^reg829) : ((8'had) >>> reg788))) ^~ (^($signed(reg771) << (~reg3520))));
                    end
                end
              reg3525 <= ((reg800 ?
                  $unsigned((^~reg3443)) : $unsigned((reg854 ?
                      forvar3465 : reg831))) <= $signed((~|$unsigned(reg750))));
            end
          else
            begin
              for (forvar3512 = (1'h0); (forvar3512 < (1'h1)); forvar3512 = (forvar3512 + (1'h1)))
                begin
                  for (forvar3513 = (1'h0); (forvar3513 < (2'h2)); forvar3513 = (forvar3513 + (1'h1)))
                    begin
                      reg3514 <= reg806;
                      reg3515 <= $signed(reg750[(2'h3):(2'h3)]);
                      reg3516 <= $signed(((~|{reg736}) >>> reg859[(2'h3):(1'h0)]));
                      reg3517 <= reg791;
                    end
                end
              if (reg3500)
                begin
                  if ({forvar3471[(3'h6):(2'h3)]})
                    begin
                      reg3518 <= ($unsigned(reg824[(4'h8):(4'h8)]) < $signed({reg750}));
                      reg3519 <= ($unsigned($signed(reg759)) | reg762);
                    end
                  else
                    begin
                      reg3518 <= $signed((~|reg753));
                      reg3519 <= ($unsigned((~$signed(reg756))) - $signed(((reg3519 & reg854) ?
                          (~reg757) : reg832[(4'h9):(2'h2)])));
                      reg3520 <= (reg3493[(3'h4):(1'h1)] == (|(&(~reg3459))));
                      reg3521 <= reg853;
                    end
                  for (forvar3522 = (1'h0); (forvar3522 < (1'h1)); forvar3522 = (forvar3522 + (1'h1)))
                    begin
                      reg3523 <= forvar3468[(2'h3):(2'h2)];
                      reg3524 <= ($signed(forvar3468) ?
                          (($unsigned(reg3499) ? $unsigned(reg3452) : reg729) ?
                              $signed(reg824) : reg3447) : (reg3467[(1'h0):(1'h0)] | $unsigned({reg3437})));
                    end
                end
              else
                begin
                  for (forvar3518 = (1'h0); (forvar3518 < (2'h2)); forvar3518 = (forvar3518 + (1'h1)))
                    begin
                      reg3519 <= $signed(($unsigned({reg818}) << $unsigned($unsigned(reg864))));
                      reg3520 <= $unsigned((|$signed($signed(reg3499))));
                      reg3521 <= reg785[(3'h6):(2'h2)];
                      reg3522 <= (forvar3458 != $unsigned(((^reg848) ?
                          reg3469 : $signed(reg3433))));
                    end
                  if (reg849[(4'hb):(4'h8)])
                    begin
                      reg3523 <= ($unsigned($unsigned(reg781[(2'h3):(2'h2)])) * $signed((reg734[(4'ha):(1'h0)] ?
                          forvar3467 : reg819)));
                      reg3524 <= (({((8'hb1) + reg732)} && (|(wire727 == reg3499))) ?
                          reg817 : reg3514[(4'h8):(1'h0)]);
                      reg3525 <= {reg3466[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg3523 <= ({reg3437[(3'h5):(1'h0)]} & reg3479[(3'h7):(3'h5)]);
                    end
                end
            end
        end
      if ($signed($unsigned((~|$unsigned(reg3482)))))
        begin
          if ($signed((reg3470[(1'h0):(1'h0)] - $signed($signed(reg759)))))
            begin
              if ($signed($unsigned((8'had))))
                begin
                  reg3526 <= (~&($signed(wire724) ?
                      ($unsigned(forvar3482) ?
                          (reg772 ^ forvar3468) : reg823) : $unsigned(forvar3461)));
                  if ($signed((reg844[(1'h1):(1'h0)] <= $unsigned(reg861[(1'h1):(1'h1)]))))
                    begin
                      reg3527 <= $signed($unsigned(reg3491[(4'h9):(2'h3)]));
                      reg3528 <= ((!reg3508[(1'h0):(1'h0)]) >= reg747);
                      reg3529 <= (-(reg3483 - forvar3496[(2'h2):(1'h0)]));
                      reg3530 <= reg3469[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3527 <= $signed((reg855[(2'h3):(2'h2)] ?
                          $signed($unsigned(reg3470)) : reg3454));
                    end
                  if (reg736[(3'h6):(3'h6)])
                    begin
                      reg3531 <= $unsigned((-$unsigned((reg3429 ?
                          wire724 : forvar3427))));
                      reg3532 <= $signed(($unsigned($signed(wire727)) ?
                          (8'ha2) : $signed(reg3483)));
                    end
                  else
                    begin
                      reg3531 <= (~^reg3513);
                      reg3532 <= reg3460[(2'h3):(1'h1)];
                    end
                end
              else
                begin
                  if ({{(((8'ha8) <= (8'h9c)) ? (~&reg3532) : {reg3527})}})
                    begin
                      reg3526 <= reg797;
                      reg3527 <= reg748;
                      reg3528 <= (^~((-reg786[(3'h5):(2'h3)]) & $unsigned($signed(reg838))));
                    end
                  else
                    begin
                      reg3526 <= (reg803[(1'h0):(1'h0)] >>> ($unsigned(((8'hb1) <= reg3526)) == (reg861 != {reg3479})));
                      reg3527 <= $signed($unsigned({$signed(forvar3468)}));
                      reg3528 <= reg783[(3'h6):(3'h5)];
                    end
                  if (($signed(reg3487[(4'h9):(4'h8)]) >>> reg731[(1'h1):(1'h1)]))
                    begin
                      reg3529 <= $unsigned(forvar3513[(2'h3):(2'h3)]);
                      reg3530 <= ($unsigned(((reg3430 - (8'haf)) ?
                          reg3527[(4'h9):(2'h3)] : (reg3429 ?
                              reg3472 : reg781))) << reg849[(1'h1):(1'h1)]);
                      reg3531 <= $signed(reg3522[(2'h3):(2'h2)]);
                      reg3532 <= $unsigned($unsigned({(~&forvar3450)}));
                    end
                  else
                    begin
                      reg3529 <= (($unsigned((|reg3443)) ?
                          (8'hae) : (~|reg3444[(1'h1):(1'h1)])) >= reg791[(1'h1):(1'h1)]);
                      reg3530 <= $unsigned((8'ha0));
                    end
                  for (forvar3533 = (1'h0); (forvar3533 < (2'h3)); forvar3533 = (forvar3533 + (1'h1)))
                    begin
                      reg3534 <= $unsigned(reg737[(1'h0):(1'h0)]);
                      reg3535 <= $signed($signed($signed($unsigned(reg3467))));
                      reg3536 <= (-reg828[(3'h7):(3'h4)]);
                    end
                end
              reg3537 <= $unsigned((8'hb3));
              for (forvar3538 = (1'h0); (forvar3538 < (1'h1)); forvar3538 = (forvar3538 + (1'h1)))
                begin
                  if (reg774)
                    begin
                      reg3539 <= ((8'hba) ? reg802[(4'hb):(3'h4)] : reg3455);
                      reg3540 <= reg744;
                    end
                  else
                    begin
                      reg3539 <= ($unsigned({forvar3458}) ?
                          (({(8'hae)} ?
                              $unsigned(reg800) : $unsigned(reg786)) ^~ ((reg3481 + reg3473) ?
                              reg791 : $unsigned((8'hb2)))) : (~|forvar3468[(1'h0):(1'h0)]));
                      reg3540 <= reg3434[(3'h4):(2'h3)];
                      reg3541 <= $unsigned((~&$signed((reg3483 | reg736))));
                      reg3542 <= (|$unsigned($unsigned((reg3466 ?
                          reg815 : reg3516))));
                    end
                  if ($unsigned(((~$signed(reg770)) ?
                      reg790 : $unsigned($signed(reg3532)))))
                    begin
                      reg3543 <= reg743;
                      reg3544 <= (^$unsigned($unsigned((reg836 == forvar3471))));
                      reg3545 <= $unsigned({(reg3517[(3'h7):(3'h5)] ?
                              $signed(reg3536) : (!reg3455))});
                      reg3546 <= $signed(forvar3461);
                    end
                  else
                    begin
                      reg3543 <= {$unsigned(($unsigned(reg843) && $signed(reg3438)))};
                    end
                  reg3547 <= (&((reg3435 ?
                      reg3515 : $signed(reg801)) <= (8'hab)));
                end
            end
          else
            begin
              if (reg3546[(1'h0):(1'h0)])
                begin
                  if (($signed($unsigned($unsigned((8'ha0)))) ?
                      (!(~&{reg3514})) : forvar3471[(4'hb):(1'h0)]))
                    begin
                      reg3526 <= forvar3450;
                      reg3527 <= {(reg865 ? reg3499 : reg733[(2'h2):(1'h1)])};
                    end
                  else
                    begin
                      reg3526 <= $unsigned(reg3463[(3'h7):(3'h6)]);
                      reg3527 <= reg861;
                    end
                end
              else
                begin
                  reg3526 <= {$unsigned(forvar3513)};
                  if ($signed(((~reg3515) ?
                      ($unsigned(reg840) > reg3546[(2'h3):(2'h2)]) : ((reg3437 && reg3437) ?
                          $signed(reg838) : forvar3461))))
                    begin
                      reg3527 <= (+reg837[(3'h5):(3'h4)]);
                      reg3528 <= reg3451;
                      reg3529 <= ($unsigned((((8'hba) ? reg823 : (8'hb4)) ?
                          reg763 : $signed(reg3514))) && $unsigned(reg745));
                    end
                  else
                    begin
                      reg3527 <= (^((+(8'hb1)) == (reg865 > ((8'ha3) ^ wire724))));
                      reg3528 <= {reg747[(2'h3):(2'h2)]};
                      reg3529 <= reg749[(4'hc):(3'h6)];
                      reg3530 <= (~reg3436[(2'h2):(1'h0)]);
                    end
                end
              for (forvar3531 = (1'h0); (forvar3531 < (1'h1)); forvar3531 = (forvar3531 + (1'h1)))
                begin
                  reg3532 <= {$unsigned($unsigned($unsigned(reg3542)))};
                end
            end
          if ($signed($unsigned(reg794)))
            begin
              reg3548 <= $signed({{reg3499}});
            end
          else
            begin
              if (($unsigned(((reg757 ?
                      reg3535 : (8'ha8)) ~^ ((8'h9c) + forvar3475))) ?
                  (($signed((8'hba)) + reg762[(3'h4):(1'h1)]) >> $unsigned((~&reg3432))) : $signed($unsigned(reg3445[(1'h0):(1'h0)]))))
                begin
                  if ($signed(forvar3476))
                    begin
                      reg3548 <= (|reg3504[(3'h5):(1'h1)]);
                      reg3549 <= $signed(((reg3474 >> (~&reg856)) ?
                          reg729 : reg781));
                      reg3550 <= forvar3428[(3'h5):(1'h1)];
                      reg3551 <= reg781;
                    end
                  else
                    begin
                      reg3548 <= $signed(forvar3471[(4'h8):(3'h5)]);
                    end
                  for (forvar3552 = (1'h0); (forvar3552 < (2'h2)); forvar3552 = (forvar3552 + (1'h1)))
                    begin
                      reg3553 <= reg3448;
                      reg3554 <= {($unsigned(((8'ha5) ?
                              reg3506 : reg3472)) || reg820)};
                    end
                  if (((^forvar3496) <= (+(forvar3467[(2'h2):(1'h0)] <= $unsigned(reg802)))))
                    begin
                      reg3555 <= (($unsigned((~&reg3463)) ?
                              (-(~&reg784)) : ((reg3509 && reg3490) * reg771)) ?
                          (^reg805[(3'h6):(2'h2)]) : (reg802 <= wire723[(1'h0):(1'h0)]));
                      reg3556 <= reg3438[(1'h1):(1'h0)];
                      reg3557 <= (($unsigned(forvar3495) * $signed((reg798 ^ reg814))) ?
                          reg3505[(2'h3):(1'h1)] : reg741[(2'h2):(2'h2)]);
                      reg3558 <= $unsigned({reg3467[(3'h6):(2'h3)]});
                    end
                  else
                    begin
                      reg3555 <= ((+reg863[(2'h3):(2'h3)]) <<< {(-(reg3504 + wire727))});
                      reg3556 <= (reg3444 >= $unsigned((|(reg825 > (8'hb7)))));
                      reg3557 <= reg3461;
                    end
                end
              else
                begin
                  for (forvar3548 = (1'h0); (forvar3548 < (2'h2)); forvar3548 = (forvar3548 + (1'h1)))
                    begin
                      reg3549 <= ($unsigned(reg3489) - reg744);
                      reg3550 <= $unsigned(reg3522);
                      reg3551 <= ((8'hb4) <= $unsigned(reg824[(3'h6):(3'h4)]));
                    end
                end
              reg3559 <= reg825[(4'ha):(3'h4)];
              for (forvar3560 = (1'h0); (forvar3560 < (1'h0)); forvar3560 = (forvar3560 + (1'h1)))
                begin
                  for (forvar3561 = (1'h0); (forvar3561 < (1'h1)); forvar3561 = (forvar3561 + (1'h1)))
                    begin
                      reg3562 <= (^~forvar3496[(1'h0):(1'h0)]);
                      reg3563 <= ((&reg3516) ?
                          (($unsigned(reg802) ?
                                  reg3473[(2'h3):(2'h2)] : forvar3450) ?
                              $signed({(8'hae)}) : (^forvar3449)) : (8'hb2));
                      reg3564 <= ($signed(($signed(reg829) & reg3448)) == $unsigned(reg3555));
                      reg3565 <= reg3513[(2'h2):(2'h2)];
                    end
                  reg3566 <= $unsigned(($unsigned($signed(reg831)) ?
                      $unsigned($unsigned(reg3437)) : ($unsigned(reg3515) >>> reg3490[(3'h5):(1'h0)])));
                  if (forvar3548[(2'h3):(1'h0)])
                    begin
                      reg3567 <= reg856[(1'h0):(1'h0)];
                      reg3568 <= (^~reg818);
                    end
                  else
                    begin
                      reg3567 <= {(~|$unsigned((^(8'ha7))))};
                      reg3568 <= {forvar3561[(3'h5):(2'h3)]};
                      reg3569 <= reg3535[(3'h5):(1'h1)];
                    end
                end
            end
        end
      else
        begin
          for (forvar3526 = (1'h0); (forvar3526 < (1'h1)); forvar3526 = (forvar3526 + (1'h1)))
            begin
              for (forvar3527 = (1'h0); (forvar3527 < (1'h1)); forvar3527 = (forvar3527 + (1'h1)))
                begin
                  if ($signed((8'hb7)))
                    begin
                      reg3528 <= forvar3458;
                      reg3529 <= ((($signed(reg863) ?
                              (+reg760) : forvar3453[(2'h2):(2'h2)]) ?
                          $signed(reg775) : reg3567[(3'h4):(2'h3)]) - (($unsigned(reg823) != reg3472[(4'he):(1'h1)]) ?
                          $unsigned((reg751 >>> reg762)) : $signed((reg851 ?
                              reg3438 : reg3448))));
                    end
                  else
                    begin
                      reg3528 <= ($signed(((~|forvar3441) ?
                          (forvar3476 >= forvar3560) : reg3442)) > reg3540[(2'h3):(2'h2)]);
                    end
                  for (forvar3530 = (1'h0); (forvar3530 < (2'h3)); forvar3530 = (forvar3530 + (1'h1)))
                    begin
                      reg3531 <= reg3461;
                      reg3532 <= $unsigned(($signed($unsigned(reg802)) ?
                          $unsigned((~^reg805)) : reg861));
                    end
                  for (forvar3533 = (1'h0); (forvar3533 < (1'h1)); forvar3533 = (forvar3533 + (1'h1)))
                    begin
                      reg3534 <= $unsigned(reg3451);
                      reg3535 <= (&$unsigned((~|{reg3463})));
                      reg3536 <= (8'hb4);
                      reg3537 <= (&((~&{reg3542}) ?
                          $signed((reg833 + (8'hb7))) : (~&wire725)));
                    end
                end
              if ($unsigned(reg833))
                begin
                  if ((reg865[(1'h1):(1'h0)] << (reg3500[(1'h0):(1'h0)] ?
                      (reg794 ?
                          (&reg3531) : $unsigned((8'haf))) : $signed(forvar3527[(3'h4):(3'h4)]))))
                    begin
                      reg3538 <= $signed(reg797);
                    end
                  else
                    begin
                      reg3538 <= {$unsigned(reg848)};
                      reg3539 <= (-(reg818 ?
                          $unsigned($signed((8'hb9))) : (~reg740)));
                    end
                  if ($signed(({(reg3454 - reg794)} & $signed((forvar3450 ?
                      reg3543 : forvar3447)))))
                    begin
                      reg3540 <= wire3425[(3'h7):(2'h3)];
                    end
                  else
                    begin
                      reg3540 <= forvar3533[(1'h0):(1'h0)];
                      reg3541 <= $signed(reg793[(4'hb):(1'h0)]);
                      reg3542 <= $unsigned(reg736);
                      reg3543 <= $signed($unsigned(((!(8'haa)) ?
                          $signed(reg3554) : (^~(8'hb6)))));
                    end
                  reg3544 <= $unsigned((^~$unsigned($unsigned((8'ha5)))));
                  for (forvar3545 = (1'h0); (forvar3545 < (1'h0)); forvar3545 = (forvar3545 + (1'h1)))
                    begin
                      reg3546 <= (8'hb8);
                      reg3547 <= (+$signed(($unsigned(reg3501) ?
                          reg3531[(2'h3):(1'h0)] : (reg3544 ^ (8'hb8)))));
                    end
                end
              else
                begin
                  for (forvar3538 = (1'h0); (forvar3538 < (2'h3)); forvar3538 = (forvar3538 + (1'h1)))
                    begin
                      reg3539 <= ($signed(((reg3448 < forvar3471) || (reg3567 ?
                          reg3502 : forvar3456))) != (+$unsigned((8'hb1))));
                      reg3540 <= (^~{reg3452});
                    end
                end
              for (forvar3548 = (1'h0); (forvar3548 < (1'h1)); forvar3548 = (forvar3548 + (1'h1)))
                begin
                  for (forvar3549 = (1'h0); (forvar3549 < (2'h2)); forvar3549 = (forvar3549 + (1'h1)))
                    begin
                      reg3550 <= {(forvar3512 ?
                              ((~reg3438) ?
                                  reg856[(3'h6):(3'h5)] : (^reg3438)) : $signed((~&(8'hab))))};
                      reg3551 <= $unsigned($unsigned(((reg738 < (8'haa)) ~^ reg3460[(1'h0):(1'h0)])));
                      reg3552 <= $unsigned(({((8'hb1) ?
                              reg3507 : reg852)} >>> (&$unsigned((8'haf)))));
                    end
                  for (forvar3553 = (1'h0); (forvar3553 < (2'h3)); forvar3553 = (forvar3553 + (1'h1)))
                    begin
                      reg3554 <= ((8'ha5) ?
                          (((reg3457 ?
                              forvar3517 : (8'hb6)) ^ $signed((8'ha8))) + $unsigned((reg769 >= reg824))) : $unsigned(reg3443));
                      reg3555 <= reg3488;
                      reg3556 <= reg815[(4'h8):(3'h7)];
                      reg3557 <= {((~|reg851) && $unsigned(reg3545))};
                    end
                end
              for (forvar3558 = (1'h0); (forvar3558 < (1'h1)); forvar3558 = (forvar3558 + (1'h1)))
                begin
                  for (forvar3559 = (1'h0); (forvar3559 < (2'h3)); forvar3559 = (forvar3559 + (1'h1)))
                    begin
                      reg3560 <= (~$signed({{(8'hb3)}}));
                      reg3561 <= reg803[(1'h0):(1'h0)];
                      reg3562 <= {(|((~^reg3448) >= ((8'hb9) ?
                              reg743 : reg788)))};
                    end
                  if (((+reg854) << $unsigned((-(~^reg798)))))
                    begin
                      reg3563 <= (|$signed(forvar3495[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg3563 <= reg3541[(4'h8):(3'h7)];
                      reg3564 <= (reg845 ?
                          (|$unsigned({reg735})) : {$signed($unsigned(forvar3517))});
                      reg3565 <= $unsigned(($unsigned((^~reg794)) <<< (8'ha9)));
                      reg3566 <= $signed($unsigned($unsigned((reg3481 == reg3485))));
                    end
                end
            end
        end
      if (reg3442)
        begin
          for (forvar3570 = (1'h0); (forvar3570 < (2'h3)); forvar3570 = (forvar3570 + (1'h1)))
            begin
              reg3571 <= (|(8'hac));
            end
          reg3572 <= ($signed($unsigned($signed((8'ha4)))) ^~ reg3511[(3'h4):(2'h3)]);
        end
      else
        begin
          if ($signed((^$signed({reg3482}))))
            begin
              if (((((~|reg831) && (reg761 ?
                      forvar3475 : (8'h9d))) * (~^$unsigned(reg3487))) ?
                  reg824[(3'h5):(3'h5)] : (!(reg3510[(3'h6):(3'h4)] ^ (reg3532 >= reg808)))))
                begin
                  if (((!reg792[(3'h4):(2'h2)]) ?
                      (reg3527[(4'h8):(3'h6)] < reg3512[(2'h3):(2'h3)]) : (8'ha7)))
                    begin
                      reg3570 <= (($unsigned($unsigned(reg3571)) & reg838[(3'h5):(1'h0)]) != reg836[(2'h3):(2'h3)]);
                      reg3571 <= $unsigned($unsigned((~|reg782[(2'h2):(2'h2)])));
                    end
                  else
                    begin
                      reg3570 <= (reg3512[(2'h3):(2'h3)] ?
                          (^((reg748 ? (8'hb8) : reg751) & reg3456)) : (8'ha4));
                      reg3571 <= $unsigned(reg3493[(2'h2):(1'h1)]);
                      reg3572 <= $signed($unsigned($unsigned((^~reg772))));
                    end
                  for (forvar3573 = (1'h0); (forvar3573 < (2'h2)); forvar3573 = (forvar3573 + (1'h1)))
                    begin
                      reg3574 <= {reg3489[(2'h2):(1'h0)]};
                    end
                  reg3575 <= (~^((wire724 ?
                          reg798[(3'h5):(2'h3)] : $signed(reg3462)) ?
                      $signed($signed(reg3483)) : ($signed(reg853) ?
                          $unsigned((8'hb3)) : (reg761 ^~ forvar3471))));
                end
              else
                begin
                  for (forvar3570 = (1'h0); (forvar3570 < (1'h1)); forvar3570 = (forvar3570 + (1'h1)))
                    begin
                      reg3571 <= ($signed($signed(wire725)) && {(&reg822)});
                    end
                end
              reg3576 <= $signed(forvar3512);
            end
          else
            begin
              if ((^$signed({(~^reg3499)})))
                begin
                  reg3570 <= reg3545[(2'h3):(1'h1)];
                  reg3571 <= (reg3512 ^ ((((8'hb7) >> forvar3538) - $unsigned((8'hb9))) ?
                      reg749 : {$signed(reg3477)}));
                  if ((forvar3552 ?
                      {(((8'ha6) + (8'hb7)) ?
                              $unsigned((8'ha9)) : (reg3464 ?
                                  reg744 : reg3554))} : $unsigned($signed(reg3566[(1'h1):(1'h1)]))))
                    begin
                      reg3572 <= $signed({reg776});
                      reg3573 <= $unsigned(reg3523);
                      reg3574 <= (~^(^~$signed(reg3480)));
                      reg3575 <= $unsigned(reg808);
                    end
                  else
                    begin
                      reg3572 <= (^(reg755[(3'h5):(3'h4)] & $unsigned($signed(reg3497))));
                      reg3573 <= ((((!(8'h9c)) ^ reg3513) <<< (^forvar3559)) ?
                          reg3520[(1'h1):(1'h1)] : reg764[(2'h2):(1'h0)]);
                      reg3574 <= reg3442[(1'h1):(1'h1)];
                      reg3575 <= {$signed(((reg829 < reg737) | $unsigned(reg3571)))};
                    end
                end
              else
                begin
                  for (forvar3570 = (1'h0); (forvar3570 < (2'h3)); forvar3570 = (forvar3570 + (1'h1)))
                    begin
                      reg3571 <= {($unsigned((reg3505 ^ reg3519)) ?
                              ({wire3425} ^~ (+reg3537)) : {$unsigned(reg3548)})};
                      reg3572 <= ($unsigned(($unsigned(reg738) ?
                              forvar3553[(4'he):(3'h6)] : forvar3548[(2'h3):(1'h0)])) ?
                          (reg3501[(1'h0):(1'h0)] >= $signed((reg3485 ?
                              reg825 : reg3432))) : reg3484[(3'h5):(2'h2)]);
                    end
                  for (forvar3573 = (1'h0); (forvar3573 < (2'h2)); forvar3573 = (forvar3573 + (1'h1)))
                    begin
                      reg3574 <= $unsigned((&reg3490[(3'h5):(1'h0)]));
                    end
                  reg3575 <= (reg3555[(3'h6):(3'h5)] ?
                      $unsigned($unsigned({wire2033})) : (reg825 < reg3485));
                end
              for (forvar3576 = (1'h0); (forvar3576 < (1'h1)); forvar3576 = (forvar3576 + (1'h1)))
                begin
                  for (forvar3577 = (1'h0); (forvar3577 < (1'h0)); forvar3577 = (forvar3577 + (1'h1)))
                    begin
                      reg3578 <= $signed(((|reg3500[(1'h1):(1'h1)]) - $unsigned((^~reg3478))));
                      reg3579 <= reg823[(2'h3):(1'h1)];
                      reg3580 <= reg815;
                    end
                  for (forvar3581 = (1'h0); (forvar3581 < (2'h2)); forvar3581 = (forvar3581 + (1'h1)))
                    begin
                      reg3582 <= (reg3494[(3'h5):(2'h3)] * reg855[(3'h5):(2'h2)]);
                      reg3583 <= (^~reg3482);
                    end
                  if ({((|(~reg794)) ? $unsigned($signed(reg737)) : reg3465)})
                    begin
                      reg3584 <= (~^(^~reg3522[(2'h3):(2'h2)]));
                      reg3585 <= ((8'h9d) ?
                          reg3452 : forvar3552[(1'h0):(1'h0)]);
                      reg3586 <= ((|$signed($signed(reg3578))) ?
                          (8'hb6) : $signed($signed(reg3555[(4'h8):(4'h8)])));
                      reg3587 <= (^~$unsigned(reg3439));
                    end
                  else
                    begin
                      reg3584 <= (~$unsigned((~^{reg776})));
                      reg3585 <= (^~(^~$unsigned($signed(reg838))));
                      reg3586 <= ({{(reg841 ?
                                  forvar3530 : reg3448)}} != $unsigned(reg3548[(3'h4):(2'h2)]));
                    end
                  if ((8'hba))
                    begin
                      reg3588 <= forvar3446[(4'hd):(4'h9)];
                    end
                  else
                    begin
                      reg3588 <= reg855[(1'h1):(1'h1)];
                      reg3589 <= forvar3545;
                    end
                end
            end
          if ((+((~|wire725[(1'h0):(1'h0)]) >>> (reg859 ?
              (~&(8'ha4)) : (reg3432 ? reg3578 : reg792)))))
            begin
              reg3590 <= (^(|(+(forvar3559 ? reg3569 : reg3443))));
              if ($signed(((~(reg3562 ? reg3445 : reg783)) && reg3431)))
                begin
                  reg3591 <= $unsigned((~((+reg3531) ?
                      forvar3449[(2'h2):(2'h2)] : $unsigned(forvar3513))));
                  reg3592 <= ($signed(reg783) ?
                      ((&(reg808 ^ reg3572)) >= ((reg3572 ?
                              forvar3581 : reg825) ?
                          {(8'hab)} : {forvar3441})) : (($unsigned(reg3485) + reg3529) ?
                          {reg739[(3'h5):(2'h2)]} : reg3444[(1'h0):(1'h0)]));
                  if (reg728[(3'h6):(1'h1)])
                    begin
                      reg3593 <= (reg3448 ?
                          reg3445 : (reg3525[(2'h3):(2'h3)] == (reg3542 + (reg3490 ?
                              reg3437 : reg750))));
                      reg3594 <= (-($unsigned($signed(reg741)) ?
                          (~^$signed(reg3463)) : $unsigned({reg3562})));
                      reg3595 <= {reg3459};
                    end
                  else
                    begin
                      reg3593 <= reg3471;
                      reg3594 <= forvar3464;
                    end
                  for (forvar3596 = (1'h0); (forvar3596 < (1'h0)); forvar3596 = (forvar3596 + (1'h1)))
                    begin
                      reg3597 <= ((((8'ha7) >= (reg813 << reg3582)) > {(-reg3539)}) ^ (8'hb0));
                      reg3598 <= $signed(forvar3538);
                      reg3599 <= {$unsigned((reg3501 > reg3549[(2'h2):(1'h0)]))};
                      reg3600 <= ((^((reg3436 ?
                          reg813 : (8'hb0)) & (forvar3517 ?
                          (8'ha9) : reg3554))) << ($signed((forvar3513 >= (8'hab))) & {$signed(forvar3471)}));
                    end
                end
              else
                begin
                  for (forvar3591 = (1'h0); (forvar3591 < (2'h2)); forvar3591 = (forvar3591 + (1'h1)))
                    begin
                      reg3592 <= $unsigned(forvar3467[(3'h5):(2'h3)]);
                    end
                end
              reg3601 <= (^~((-$signed(reg836)) ?
                  $signed((~^reg3536)) : ($unsigned(reg860) ?
                      $signed(reg864) : reg3526)));
              reg3602 <= ((((^~reg831) ?
                          $unsigned(forvar3596) : (forvar3461 ?
                              reg3573 : forvar3570)) ?
                      $unsigned($signed((8'hb1))) : {{reg3563}}) ?
                  ((~|reg3598) - reg728) : reg3555);
            end
          else
            begin
              for (forvar3590 = (1'h0); (forvar3590 < (1'h1)); forvar3590 = (forvar3590 + (1'h1)))
                begin
                  for (forvar3591 = (1'h0); (forvar3591 < (2'h2)); forvar3591 = (forvar3591 + (1'h1)))
                    begin
                      reg3592 <= ((+reg3569[(4'h9):(1'h1)]) ?
                          $unsigned(((reg3561 > (8'hb8)) >= (reg808 | reg856))) : (forvar3461[(1'h0):(1'h0)] << reg864[(1'h0):(1'h0)]));
                    end
                end
            end
          for (forvar3603 = (1'h0); (forvar3603 < (2'h3)); forvar3603 = (forvar3603 + (1'h1)))
            begin
              for (forvar3604 = (1'h0); (forvar3604 < (1'h1)); forvar3604 = (forvar3604 + (1'h1)))
                begin
                  if ($signed(((reg3447[(4'hb):(4'ha)] - (reg3494 ?
                          reg758 : reg752)) ?
                      (reg3583[(1'h1):(1'h0)] + $signed(reg855)) : (+forvar3596))))
                    begin
                      reg3605 <= reg781[(3'h4):(2'h2)];
                      reg3606 <= reg3519;
                    end
                  else
                    begin
                      reg3605 <= reg3510;
                      reg3606 <= reg3454[(1'h1):(1'h1)];
                      reg3607 <= {reg775[(4'ha):(3'h5)]};
                      reg3608 <= ({reg3515} ?
                          $unsigned(reg784) : {($unsigned(reg3431) ^~ $unsigned(reg3452))});
                    end
                  for (forvar3609 = (1'h0); (forvar3609 < (2'h3)); forvar3609 = (forvar3609 + (1'h1)))
                    begin
                      reg3610 <= $unsigned($signed(((~&forvar3596) ?
                          reg747[(1'h0):(1'h0)] : reg814[(1'h0):(1'h0)])));
                      reg3611 <= ((forvar3461[(2'h3):(1'h0)] * ((reg3520 | reg864) ?
                              (reg3491 ^~ reg846) : reg3460)) ?
                          ((~|$unsigned(reg3469)) + ($signed(reg806) ^ (reg3476 ?
                              reg828 : reg3576))) : ($unsigned(reg744) ?
                              $signed(reg809) : (^~$signed(reg786))));
                      reg3612 <= $signed((^(|forvar3526)));
                    end
                  for (forvar3613 = (1'h0); (forvar3613 < (1'h1)); forvar3613 = (forvar3613 + (1'h1)))
                    begin
                      reg3614 <= (8'ha7);
                      reg3615 <= (((forvar3538 && $unsigned(reg3567)) ?
                              (~(reg3525 - reg734)) : reg3551[(1'h0):(1'h0)]) ?
                          $unsigned($unsigned((forvar3513 == reg3447))) : $unsigned(reg3524));
                      reg3616 <= {($unsigned(reg3483[(2'h2):(2'h2)]) * $signed(((8'h9e) ?
                              reg738 : (8'haa))))};
                      reg3617 <= (^(&$unsigned((reg3578 >>> (8'ha6)))));
                    end
                  if (({((wire726 >>> reg794) ?
                              $signed(reg810) : reg790[(4'he):(4'hc)])} ?
                      forvar3440[(4'he):(4'hc)] : (reg3592 ~^ (~|(forvar3495 - reg825)))))
                    begin
                      reg3618 <= reg3532[(3'h6):(2'h2)];
                      reg3619 <= reg749[(1'h0):(1'h0)];
                      reg3620 <= reg3438;
                      reg3621 <= (~|({forvar3552} * ((!(8'ha6)) | ((8'hb4) ?
                          reg3514 : reg784))));
                    end
                  else
                    begin
                      reg3618 <= $unsigned($signed($unsigned((reg3471 ?
                          (8'haa) : reg3506))));
                      reg3619 <= {({$signed(reg3552)} && ((reg795 ?
                                  reg3547 : reg3497) ?
                              $unsigned((8'haa)) : $signed(reg3559)))};
                      reg3620 <= ((~^($unsigned(reg765) ?
                          (reg3473 ?
                              reg3471 : reg799) : $unsigned(reg793))) != reg777[(3'h7):(1'h1)]);
                      reg3621 <= ((((!(8'ha3)) ?
                              (8'haa) : (wire3425 >>> reg3448)) != {(reg3528 ?
                                  reg782 : reg769)}) ?
                          $signed(($signed(reg768) ?
                              (reg747 ?
                                  reg819 : reg3579) : $unsigned(forvar3545))) : $unsigned(({reg3530} == (reg761 ~^ reg793))));
                    end
                end
              for (forvar3622 = (1'h0); (forvar3622 < (1'h1)); forvar3622 = (forvar3622 + (1'h1)))
                begin
                  if ((($unsigned((^~reg3433)) ?
                          (^~(~wire727)) : ((reg3454 ^~ reg3508) ?
                              (~&reg738) : forvar3522[(2'h2):(1'h1)])) ?
                      (~|($signed(forvar3553) ?
                          (forvar3591 ?
                              reg3510 : reg3456) : reg3464[(1'h1):(1'h0)])) : ((8'ha1) ?
                          ((forvar3482 ? reg860 : reg799) ?
                              reg802[(4'ha):(3'h6)] : reg3521[(3'h6):(1'h0)]) : reg3550[(2'h2):(1'h1)])))
                    begin
                      reg3623 <= $unsigned((!(~^(reg3566 ? reg765 : (8'had)))));
                      reg3624 <= $signed($signed(reg730[(2'h2):(1'h0)]));
                      reg3625 <= $unsigned((reg3437[(4'h8):(4'h8)] | (8'haf)));
                      reg3626 <= {reg846};
                    end
                  else
                    begin
                      reg3623 <= (($signed(reg3485) > ((reg791 ^ reg792) ?
                              {forvar3526} : (forvar3427 ? reg806 : (8'ha2)))) ?
                          reg758 : $signed(reg3623));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      reg3627 <= (&$signed(reg3548[(2'h3):(2'h2)]));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module513  (y, clk, wire518, wire517, wire516, wire515, wire514);
  output wire [(32'h916):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire518;
  input wire [(4'hc):(1'h0)] wire517;
  input wire signed [(3'h6):(1'h0)] wire516;
  input wire [(3'h4):(1'h0)] wire515;
  input wire signed [(4'hd):(1'h0)] wire514;
  wire signed [(3'h6):(1'h0)] wire717;
  wire [(3'h7):(1'h0)] wire716;
  wire [(4'hd):(1'h0)] wire715;
  reg [(4'h9):(1'h0)] reg714 = (1'h0);
  reg [(2'h3):(1'h0)] reg713 = (1'h0);
  reg [(4'he):(1'h0)] reg701 = (1'h0);
  reg [(4'hc):(1'h0)] reg712 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg711 = (1'h0);
  reg [(5'h10):(1'h0)] reg710 = (1'h0);
  reg [(3'h5):(1'h0)] reg709 = (1'h0);
  reg signed [(4'he):(1'h0)] reg708 = (1'h0);
  reg [(4'hc):(1'h0)] reg707 = (1'h0);
  reg [(2'h3):(1'h0)] reg706 = (1'h0);
  reg [(3'h4):(1'h0)] reg704 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg703 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg702 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg700 = (1'h0);
  reg [(2'h3):(1'h0)] reg699 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg698 = (1'h0);
  reg [(4'h9):(1'h0)] reg697 = (1'h0);
  reg [(3'h5):(1'h0)] reg696 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg695 = (1'h0);
  reg [(4'hd):(1'h0)] reg693 = (1'h0);
  reg [(2'h2):(1'h0)] reg692 = (1'h0);
  reg [(2'h3):(1'h0)] reg691 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg690 = (1'h0);
  reg [(2'h2):(1'h0)] reg689 = (1'h0);
  reg [(4'hd):(1'h0)] reg688 = (1'h0);
  reg [(4'hf):(1'h0)] reg687 = (1'h0);
  reg signed [(4'he):(1'h0)] reg685 = (1'h0);
  reg [(4'h8):(1'h0)] reg683 = (1'h0);
  reg [(4'hb):(1'h0)] reg671 = (1'h0);
  reg [(3'h4):(1'h0)] reg658 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg657 = (1'h0);
  reg [(4'he):(1'h0)] reg653 = (1'h0);
  reg [(4'h8):(1'h0)] reg648 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg647 = (1'h0);
  reg [(2'h3):(1'h0)] reg645 = (1'h0);
  reg signed [(4'he):(1'h0)] reg684 = (1'h0);
  reg [(4'hf):(1'h0)] reg682 = (1'h0);
  reg [(4'h9):(1'h0)] reg674 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg668 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg681 = (1'h0);
  reg [(4'hc):(1'h0)] reg680 = (1'h0);
  reg [(4'hc):(1'h0)] reg679 = (1'h0);
  reg [(3'h7):(1'h0)] reg678 = (1'h0);
  reg [(2'h3):(1'h0)] reg677 = (1'h0);
  reg [(3'h4):(1'h0)] reg676 = (1'h0);
  reg [(4'hc):(1'h0)] reg675 = (1'h0);
  reg [(4'hf):(1'h0)] reg673 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg672 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg670 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg669 = (1'h0);
  reg [(4'h9):(1'h0)] reg667 = (1'h0);
  reg [(4'hc):(1'h0)] reg666 = (1'h0);
  reg [(3'h7):(1'h0)] reg665 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg664 = (1'h0);
  reg [(3'h6):(1'h0)] reg663 = (1'h0);
  reg [(4'h8):(1'h0)] reg662 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg661 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg660 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg659 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg656 = (1'h0);
  reg [(3'h7):(1'h0)] reg655 = (1'h0);
  reg [(2'h2):(1'h0)] reg654 = (1'h0);
  reg [(3'h6):(1'h0)] reg652 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg651 = (1'h0);
  reg [(2'h3):(1'h0)] reg650 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg649 = (1'h0);
  reg [(3'h6):(1'h0)] reg646 = (1'h0);
  reg [(2'h2):(1'h0)] reg629 = (1'h0);
  reg [(2'h3):(1'h0)] reg636 = (1'h0);
  reg [(4'he):(1'h0)] reg635 = (1'h0);
  reg [(4'hc):(1'h0)] reg633 = (1'h0);
  reg [(4'hf):(1'h0)] reg644 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg643 = (1'h0);
  reg [(5'h10):(1'h0)] reg641 = (1'h0);
  reg [(2'h3):(1'h0)] reg640 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg638 = (1'h0);
  reg [(3'h7):(1'h0)] reg637 = (1'h0);
  reg [(4'h8):(1'h0)] reg634 = (1'h0);
  reg [(3'h4):(1'h0)] reg632 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg631 = (1'h0);
  reg [(3'h6):(1'h0)] reg630 = (1'h0);
  reg [(4'hd):(1'h0)] reg628 = (1'h0);
  reg [(5'h10):(1'h0)] reg625 = (1'h0);
  reg [(4'ha):(1'h0)] reg624 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg623 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg620 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg619 = (1'h0);
  reg signed [(4'he):(1'h0)] reg618 = (1'h0);
  reg [(5'h10):(1'h0)] reg616 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg602 = (1'h0);
  reg [(4'ha):(1'h0)] reg613 = (1'h0);
  reg [(4'ha):(1'h0)] reg612 = (1'h0);
  reg [(3'h5):(1'h0)] reg611 = (1'h0);
  reg [(3'h6):(1'h0)] reg610 = (1'h0);
  reg [(3'h6):(1'h0)] reg609 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg608 = (1'h0);
  reg [(3'h5):(1'h0)] reg607 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg606 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg605 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg604 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg603 = (1'h0);
  reg [(4'hd):(1'h0)] reg601 = (1'h0);
  reg [(4'hf):(1'h0)] reg600 = (1'h0);
  reg [(3'h5):(1'h0)] reg599 = (1'h0);
  reg [(4'h8):(1'h0)] reg598 = (1'h0);
  reg [(3'h6):(1'h0)] reg597 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg596 = (1'h0);
  reg [(4'hb):(1'h0)] reg594 = (1'h0);
  reg [(3'h6):(1'h0)] reg592 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg591 = (1'h0);
  reg [(3'h5):(1'h0)] reg590 = (1'h0);
  reg [(4'hb):(1'h0)] reg589 = (1'h0);
  reg [(4'hc):(1'h0)] reg588 = (1'h0);
  reg [(4'h9):(1'h0)] reg587 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg586 = (1'h0);
  reg [(3'h5):(1'h0)] reg585 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg584 = (1'h0);
  reg signed [(4'he):(1'h0)] reg583 = (1'h0);
  reg [(3'h6):(1'h0)] reg582 = (1'h0);
  reg [(5'h10):(1'h0)] reg580 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg579 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg576 = (1'h0);
  reg [(4'hf):(1'h0)] reg578 = (1'h0);
  reg [(5'h10):(1'h0)] reg577 = (1'h0);
  reg [(2'h3):(1'h0)] reg575 = (1'h0);
  reg [(4'hc):(1'h0)] reg574 = (1'h0);
  reg [(5'h10):(1'h0)] reg573 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg572 = (1'h0);
  reg [(4'hf):(1'h0)] reg571 = (1'h0);
  reg [(4'hd):(1'h0)] reg569 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg568 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg567 = (1'h0);
  reg [(4'h9):(1'h0)] reg563 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg556 = (1'h0);
  reg [(4'h9):(1'h0)] reg555 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg554 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg566 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg565 = (1'h0);
  reg [(5'h10):(1'h0)] reg564 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg562 = (1'h0);
  reg [(4'ha):(1'h0)] reg561 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg560 = (1'h0);
  reg [(4'hc):(1'h0)] reg559 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg558 = (1'h0);
  reg [(4'h9):(1'h0)] reg557 = (1'h0);
  reg [(4'hf):(1'h0)] reg553 = (1'h0);
  reg [(3'h4):(1'h0)] reg552 = (1'h0);
  reg [(4'hf):(1'h0)] reg543 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg538 = (1'h0);
  reg [(4'hc):(1'h0)] reg551 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg548 = (1'h0);
  reg [(5'h10):(1'h0)] reg547 = (1'h0);
  reg [(4'hf):(1'h0)] reg546 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg545 = (1'h0);
  reg signed [(4'he):(1'h0)] reg534 = (1'h0);
  reg [(3'h5):(1'h0)] reg542 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg541 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg540 = (1'h0);
  reg [(3'h5):(1'h0)] reg539 = (1'h0);
  reg [(4'hc):(1'h0)] reg537 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg536 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg535 = (1'h0);
  reg [(3'h4):(1'h0)] reg533 = (1'h0);
  reg [(4'h9):(1'h0)] reg532 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg531 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg530 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg527 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg526 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg524 = (1'h0);
  reg [(4'ha):(1'h0)] reg523 = (1'h0);
  reg [(3'h7):(1'h0)] reg522 = (1'h0);
  reg [(2'h3):(1'h0)] forvar710 = (1'h0);
  reg [(2'h3):(1'h0)] forvar709 = (1'h0);
  reg [(4'ha):(1'h0)] forvar700 = (1'h0);
  reg [(2'h2):(1'h0)] forvar695 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar705 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar701 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar694 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar686 = (1'h0);
  reg [(4'hb):(1'h0)] forvar681 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar677 = (1'h0);
  reg [(4'h9):(1'h0)] forvar672 = (1'h0);
  reg [(4'ha):(1'h0)] forvar670 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar664 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar663 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar660 = (1'h0);
  reg [(4'hf):(1'h0)] forvar651 = (1'h0);
  reg [(4'hb):(1'h0)] forvar646 = (1'h0);
  reg [(4'ha):(1'h0)] forvar683 = (1'h0);
  reg [(4'hf):(1'h0)] forvar678 = (1'h0);
  reg [(3'h7):(1'h0)] forvar676 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar674 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar671 = (1'h0);
  reg [(4'h9):(1'h0)] forvar668 = (1'h0);
  reg [(4'hf):(1'h0)] forvar658 = (1'h0);
  reg [(3'h6):(1'h0)] forvar657 = (1'h0);
  reg [(4'hf):(1'h0)] forvar653 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar648 = (1'h0);
  reg [(4'hc):(1'h0)] forvar647 = (1'h0);
  reg [(4'hd):(1'h0)] forvar645 = (1'h0);
  reg [(4'ha):(1'h0)] forvar630 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar632 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar642 = (1'h0);
  reg [(4'hc):(1'h0)] forvar639 = (1'h0);
  reg [(4'hb):(1'h0)] forvar636 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar635 = (1'h0);
  reg [(4'ha):(1'h0)] forvar633 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar629 = (1'h0);
  reg [(3'h6):(1'h0)] forvar627 = (1'h0);
  reg [(4'h9):(1'h0)] forvar626 = (1'h0);
  reg [(4'h8):(1'h0)] forvar622 = (1'h0);
  reg [(4'he):(1'h0)] forvar621 = (1'h0);
  reg [(4'h9):(1'h0)] forvar617 = (1'h0);
  reg [(3'h4):(1'h0)] forvar615 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar614 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar604 = (1'h0);
  reg [(2'h3):(1'h0)] forvar601 = (1'h0);
  reg [(3'h7):(1'h0)] forvar602 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar595 = (1'h0);
  reg [(4'hd):(1'h0)] forvar593 = (1'h0);
  reg [(3'h6):(1'h0)] forvar583 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar581 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar578 = (1'h0);
  reg [(2'h3):(1'h0)] forvar576 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar570 = (1'h0);
  reg [(4'h9):(1'h0)] forvar565 = (1'h0);
  reg [(4'hc):(1'h0)] forvar559 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar553 = (1'h0);
  reg [(4'hf):(1'h0)] forvar563 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar556 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar555 = (1'h0);
  reg [(4'hb):(1'h0)] forvar554 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar545 = (1'h0);
  reg [(4'h8):(1'h0)] forvar542 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar539 = (1'h0);
  reg [(4'hc):(1'h0)] forvar550 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar549 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar544 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar543 = (1'h0);
  reg [(4'hf):(1'h0)] forvar538 = (1'h0);
  reg [(4'hc):(1'h0)] forvar534 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar529 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar528 = (1'h0);
  reg [(4'hf):(1'h0)] forvar525 = (1'h0);
  reg [(4'ha):(1'h0)] forvar521 = (1'h0);
  reg [(4'he):(1'h0)] forvar520 = (1'h0);
  reg [(5'h10):(1'h0)] forvar519 = (1'h0);
  assign y = {wire717,
                 wire716,
                 wire715,
                 reg714,
                 reg713,
                 reg701,
                 reg712,
                 reg711,
                 reg710,
                 reg709,
                 reg708,
                 reg707,
                 reg706,
                 reg704,
                 reg703,
                 reg702,
                 reg700,
                 reg699,
                 reg698,
                 reg697,
                 reg696,
                 reg695,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg689,
                 reg688,
                 reg687,
                 reg685,
                 reg683,
                 reg671,
                 reg658,
                 reg657,
                 reg653,
                 reg648,
                 reg647,
                 reg645,
                 reg684,
                 reg682,
                 reg674,
                 reg668,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg676,
                 reg675,
                 reg673,
                 reg672,
                 reg670,
                 reg669,
                 reg667,
                 reg666,
                 reg665,
                 reg664,
                 reg663,
                 reg662,
                 reg661,
                 reg660,
                 reg659,
                 reg656,
                 reg655,
                 reg654,
                 reg652,
                 reg651,
                 reg650,
                 reg649,
                 reg646,
                 reg629,
                 reg636,
                 reg635,
                 reg633,
                 reg644,
                 reg643,
                 reg641,
                 reg640,
                 reg638,
                 reg637,
                 reg634,
                 reg632,
                 reg631,
                 reg630,
                 reg628,
                 reg625,
                 reg624,
                 reg623,
                 reg620,
                 reg619,
                 reg618,
                 reg616,
                 reg602,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg594,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg580,
                 reg579,
                 reg576,
                 reg578,
                 reg577,
                 reg575,
                 reg574,
                 reg573,
                 reg572,
                 reg571,
                 reg569,
                 reg568,
                 reg567,
                 reg563,
                 reg556,
                 reg555,
                 reg554,
                 reg566,
                 reg565,
                 reg564,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 reg553,
                 reg552,
                 reg543,
                 reg538,
                 reg551,
                 reg548,
                 reg547,
                 reg546,
                 reg545,
                 reg534,
                 reg542,
                 reg541,
                 reg540,
                 reg539,
                 reg537,
                 reg536,
                 reg535,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg527,
                 reg526,
                 reg524,
                 reg523,
                 reg522,
                 forvar710,
                 forvar709,
                 forvar700,
                 forvar695,
                 forvar705,
                 forvar701,
                 forvar694,
                 forvar686,
                 forvar681,
                 forvar677,
                 forvar672,
                 forvar670,
                 forvar664,
                 forvar663,
                 forvar660,
                 forvar651,
                 forvar646,
                 forvar683,
                 forvar678,
                 forvar676,
                 forvar674,
                 forvar671,
                 forvar668,
                 forvar658,
                 forvar657,
                 forvar653,
                 forvar648,
                 forvar647,
                 forvar645,
                 forvar630,
                 forvar632,
                 forvar642,
                 forvar639,
                 forvar636,
                 forvar635,
                 forvar633,
                 forvar629,
                 forvar627,
                 forvar626,
                 forvar622,
                 forvar621,
                 forvar617,
                 forvar615,
                 forvar614,
                 forvar604,
                 forvar601,
                 forvar602,
                 forvar595,
                 forvar593,
                 forvar583,
                 forvar581,
                 forvar578,
                 forvar576,
                 forvar570,
                 forvar565,
                 forvar559,
                 forvar553,
                 forvar563,
                 forvar556,
                 forvar555,
                 forvar554,
                 forvar545,
                 forvar542,
                 forvar539,
                 forvar550,
                 forvar549,
                 forvar544,
                 forvar543,
                 forvar538,
                 forvar534,
                 forvar529,
                 forvar528,
                 forvar525,
                 forvar521,
                 forvar520,
                 forvar519,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar519 = (1'h0); (forvar519 < (2'h2)); forvar519 = (forvar519 + (1'h1)))
        begin
          for (forvar520 = (1'h0); (forvar520 < (1'h1)); forvar520 = (forvar520 + (1'h1)))
            begin
              if (forvar519[(1'h1):(1'h0)])
                begin
                  for (forvar521 = (1'h0); (forvar521 < (1'h1)); forvar521 = (forvar521 + (1'h1)))
                    begin
                      reg522 <= (((&forvar520[(4'hd):(3'h5)]) ?
                              wire514[(4'h9):(1'h0)] : (+{(8'had)})) ?
                          forvar521[(3'h4):(2'h3)] : $signed((^$signed(forvar520))));
                      reg523 <= (wire516[(2'h2):(1'h1)] ?
                          (&$unsigned($signed(wire518))) : (wire518[(4'ha):(3'h5)] << reg522[(3'h6):(2'h3)]));
                      reg524 <= ($signed((~(wire516 ?
                          wire517 : wire516))) <= {((wire516 ?
                                  (8'hb7) : forvar521) ?
                              {(8'haf)} : reg522[(3'h5):(3'h4)])});
                    end
                  for (forvar525 = (1'h0); (forvar525 < (2'h3)); forvar525 = (forvar525 + (1'h1)))
                    begin
                      reg526 <= (reg523 ^ (^$signed(reg523[(2'h3):(2'h2)])));
                      reg527 <= $unsigned(forvar520);
                    end
                end
              else
                begin
                  for (forvar521 = (1'h0); (forvar521 < (2'h3)); forvar521 = (forvar521 + (1'h1)))
                    begin
                      reg522 <= wire517[(4'h8):(1'h1)];
                      reg523 <= $signed({reg527[(1'h0):(1'h0)]});
                      reg524 <= (forvar521[(1'h1):(1'h1)] && wire517);
                    end
                end
            end
          for (forvar528 = (1'h0); (forvar528 < (2'h3)); forvar528 = (forvar528 + (1'h1)))
            begin
              for (forvar529 = (1'h0); (forvar529 < (2'h2)); forvar529 = (forvar529 + (1'h1)))
                begin
                  if ((reg524[(3'h6):(3'h4)] ?
                      $signed(($signed((8'hb4)) >= {reg526})) : (reg527[(4'ha):(4'h9)] ?
                          forvar528 : reg524[(4'h8):(2'h3)])))
                    begin
                      reg530 <= ({((!wire517) >> forvar520)} ?
                          (reg524 | ((wire516 ? (8'ha8) : wire517) ?
                              $signed((8'hab)) : ((8'h9e) ?
                                  (8'ha1) : forvar525))) : (reg527 != wire516));
                      reg531 <= (wire517[(3'h5):(3'h5)] * $unsigned(($signed(reg526) ^ $unsigned(wire516))));
                    end
                  else
                    begin
                      reg530 <= (+$unsigned((~$unsigned(wire516))));
                      reg531 <= (!$unsigned(($unsigned(wire515) ^~ $signed(wire516))));
                      reg532 <= reg531;
                      reg533 <= $signed(({$unsigned((8'ha5))} ?
                          reg532 : $unsigned(reg527)));
                    end
                end
            end
          if (wire516[(1'h0):(1'h0)])
            begin
              if (forvar529[(3'h5):(1'h1)])
                begin
                  for (forvar534 = (1'h0); (forvar534 < (1'h0)); forvar534 = (forvar534 + (1'h1)))
                    begin
                      reg535 <= (^reg522[(3'h7):(1'h1)]);
                    end
                  reg536 <= $unsigned((-wire515));
                  reg537 <= ($unsigned(reg522[(3'h5):(3'h4)]) == (^wire515[(3'h4):(1'h1)]));
                  for (forvar538 = (1'h0); (forvar538 < (2'h2)); forvar538 = (forvar538 + (1'h1)))
                    begin
                      reg539 <= {$signed((~^forvar534[(1'h1):(1'h0)]))};
                      reg540 <= $unsigned($signed($signed((^~reg526))));
                      reg541 <= $signed(forvar521[(3'h4):(2'h2)]);
                      reg542 <= {wire517[(3'h5):(2'h3)]};
                    end
                end
              else
                begin
                  reg534 <= $signed(wire514[(4'hd):(1'h0)]);
                  reg535 <= reg526[(3'h7):(2'h2)];
                end
              for (forvar543 = (1'h0); (forvar543 < (2'h3)); forvar543 = (forvar543 + (1'h1)))
                begin
                  for (forvar544 = (1'h0); (forvar544 < (1'h1)); forvar544 = (forvar544 + (1'h1)))
                    begin
                      reg545 <= $signed(reg532[(3'h5):(1'h1)]);
                      reg546 <= reg533;
                      reg547 <= $unsigned((forvar528[(4'h8):(3'h7)] ?
                          reg541 : $signed($signed(wire517))));
                      reg548 <= $signed((~|$unsigned($unsigned(forvar528))));
                    end
                end
              for (forvar549 = (1'h0); (forvar549 < (1'h0)); forvar549 = (forvar549 + (1'h1)))
                begin
                  for (forvar550 = (1'h0); (forvar550 < (1'h1)); forvar550 = (forvar550 + (1'h1)))
                    begin
                      reg551 <= reg545[(4'hb):(4'hb)];
                    end
                end
            end
          else
            begin
              if ($signed((~^{(forvar550 ? wire518 : forvar525)})))
                begin
                  reg534 <= {$unsigned($unsigned((^~reg539)))};
                  if (reg540[(3'h5):(1'h0)])
                    begin
                      reg535 <= $signed($signed($signed(reg534)));
                      reg536 <= (^$signed({(forvar525 ^~ reg526)}));
                    end
                  else
                    begin
                      reg535 <= ((|(((8'ha0) + forvar549) < (8'hb1))) ?
                          ((~$signed(reg532)) ?
                              (+$unsigned(forvar550)) : (forvar549 ?
                                  reg548[(2'h3):(1'h0)] : reg537)) : reg542[(3'h5):(2'h2)]);
                    end
                  reg537 <= reg541;
                end
              else
                begin
                  if ((($unsigned(reg531[(2'h3):(2'h3)]) ?
                          (forvar529 ?
                              (8'ha9) : $unsigned(forvar549)) : (8'ha0)) ?
                      $signed(((reg531 ?
                          reg546 : reg539) ^ (8'ha5))) : (reg542 ?
                          {(&reg523)} : forvar550)))
                    begin
                      reg534 <= (($unsigned({forvar543}) ?
                          $signed(reg524) : ((reg537 != forvar550) ^ $signed(reg545))) != $signed(forvar529[(1'h0):(1'h0)]));
                      reg535 <= $unsigned(($unsigned((reg539 ?
                          (8'hb2) : reg530)) > $signed(forvar534)));
                      reg536 <= $signed((~^reg522));
                    end
                  else
                    begin
                      reg534 <= (+forvar534[(3'h7):(3'h4)]);
                    end
                  if ({($signed(reg536) != wire516)})
                    begin
                      reg537 <= ((reg524 ?
                          (&(forvar525 | reg534)) : reg527) * (wire516 ?
                          ((^~reg542) <= reg527[(3'h7):(1'h1)]) : forvar534));
                      reg538 <= ({reg545} - $unsigned($unsigned((wire518 ?
                          reg545 : reg542))));
                    end
                  else
                    begin
                      reg537 <= reg537;
                    end
                  for (forvar539 = (1'h0); (forvar539 < (1'h1)); forvar539 = (forvar539 + (1'h1)))
                    begin
                      reg540 <= ({(^~(reg548 ? reg546 : reg536))} | forvar539);
                      reg541 <= forvar544;
                    end
                  for (forvar542 = (1'h0); (forvar542 < (2'h3)); forvar542 = (forvar542 + (1'h1)))
                    begin
                      reg543 <= forvar539[(4'he):(4'h8)];
                    end
                end
              for (forvar544 = (1'h0); (forvar544 < (1'h0)); forvar544 = (forvar544 + (1'h1)))
                begin
                  for (forvar545 = (1'h0); (forvar545 < (1'h1)); forvar545 = (forvar545 + (1'h1)))
                    begin
                      reg546 <= (^~$signed(forvar529[(2'h3):(2'h3)]));
                      reg547 <= ((-($signed(forvar529) ?
                              $unsigned(reg548) : forvar528[(3'h6):(2'h2)])) ?
                          reg531[(3'h6):(2'h3)] : reg551);
                      reg548 <= ({wire518} ^ ($unsigned((reg534 ?
                          reg539 : reg545)) | $signed(((8'hab) & (8'h9e)))));
                    end
                end
            end
        end
      reg552 <= reg534;
      if (reg552[(2'h2):(1'h0)])
        begin
          reg553 <= $unsigned(forvar550);
          for (forvar554 = (1'h0); (forvar554 < (1'h0)); forvar554 = (forvar554 + (1'h1)))
            begin
              for (forvar555 = (1'h0); (forvar555 < (1'h1)); forvar555 = (forvar555 + (1'h1)))
                begin
                  for (forvar556 = (1'h0); (forvar556 < (2'h3)); forvar556 = (forvar556 + (1'h1)))
                    begin
                      reg557 <= ((($signed(reg551) ^~ reg534[(3'h4):(2'h3)]) == {{reg526}}) ?
                          (forvar545 << (^(forvar539 ?
                              (8'h9d) : forvar550))) : {((reg538 ?
                                  forvar525 : forvar542) || ((8'hac) ?
                                  reg551 : reg546))});
                    end
                end
              reg558 <= $unsigned($signed((+$unsigned(reg538))));
              if ($signed((^(&$signed(forvar525)))))
                begin
                  reg559 <= (|$unsigned(forvar539));
                  if ({((wire517 ^~ $unsigned((8'haa))) >> forvar528)})
                    begin
                      reg560 <= ({reg522[(2'h2):(1'h0)]} ?
                          ($signed(wire514[(3'h5):(3'h4)]) ?
                              (^$unsigned(reg537)) : (!(8'hb4))) : forvar555[(3'h6):(2'h2)]);
                      reg561 <= reg530;
                    end
                  else
                    begin
                      reg560 <= (reg548[(1'h0):(1'h0)] - reg542);
                      reg561 <= $signed({reg561[(3'h7):(1'h0)]});
                      reg562 <= reg531[(4'h9):(3'h6)];
                    end
                  for (forvar563 = (1'h0); (forvar563 < (1'h0)); forvar563 = (forvar563 + (1'h1)))
                    begin
                      reg564 <= (reg546 > $unsigned($signed($unsigned(forvar554))));
                      reg565 <= {(reg533[(3'h4):(1'h1)] ?
                              (~reg539[(3'h5):(2'h2)]) : (-(forvar554 ?
                                  reg522 : (8'hb0))))};
                      reg566 <= reg557;
                    end
                end
              else
                begin
                  if (reg557[(2'h2):(1'h0)])
                    begin
                      reg559 <= ($unsigned($unsigned(reg548[(1'h0):(1'h0)])) ?
                          wire514[(2'h3):(1'h0)] : $signed((reg545[(3'h6):(1'h1)] < (reg543 ?
                              reg559 : reg538))));
                      reg560 <= (8'h9d);
                      reg561 <= $signed((($signed(reg527) && (~|reg557)) ?
                          {$unsigned(reg557)} : $signed((reg545 <<< reg534))));
                    end
                  else
                    begin
                      reg559 <= (forvar554[(4'h8):(3'h7)] == $signed(reg527));
                      reg560 <= $signed(reg565);
                      reg561 <= (|(+reg530));
                    end
                end
            end
        end
      else
        begin
          for (forvar553 = (1'h0); (forvar553 < (1'h1)); forvar553 = (forvar553 + (1'h1)))
            begin
              reg554 <= reg535[(2'h2):(1'h0)];
              if ((forvar520 - $signed($unsigned((reg566 >>> forvar543)))))
                begin
                  if (($unsigned($signed((reg552 ?
                      forvar539 : forvar543))) >= $signed(($signed((8'ha8)) == ((8'hae) ?
                      reg530 : (8'h9f))))))
                    begin
                      reg555 <= $signed((&reg538));
                      reg556 <= {($signed($signed(reg552)) ?
                              forvar550 : (reg543 ?
                                  forvar545[(3'h4):(2'h2)] : $unsigned(reg533)))};
                      reg557 <= ((^~reg524) ?
                          $unsigned((reg535 ?
                              reg543[(4'hd):(2'h2)] : $unsigned(forvar525))) : ($unsigned({reg556}) != $signed($signed((8'hab)))));
                      reg558 <= $unsigned({$unsigned((reg537 > reg547))});
                    end
                  else
                    begin
                      reg555 <= $signed(reg527);
                    end
                  for (forvar559 = (1'h0); (forvar559 < (1'h1)); forvar559 = (forvar559 + (1'h1)))
                    begin
                      reg560 <= {($unsigned($signed((8'ha7))) == (~$signed(wire518)))};
                      reg561 <= (!forvar549);
                      reg562 <= reg557;
                    end
                  if (forvar543[(4'h8):(3'h5)])
                    begin
                      reg563 <= $unsigned(reg554);
                    end
                  else
                    begin
                      reg563 <= reg531[(1'h1):(1'h1)];
                      reg564 <= $signed($signed(forvar538[(4'he):(4'hb)]));
                    end
                end
              else
                begin
                  if (((forvar525 ?
                          (^(^~reg562)) : ({reg536} ?
                              (~^reg532) : (^forvar543))) ?
                      reg548[(3'h5):(1'h1)] : reg551[(3'h4):(1'h1)]))
                    begin
                      reg555 <= reg547[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg555 <= reg532[(1'h0):(1'h0)];
                      reg556 <= forvar542;
                      reg557 <= wire517;
                      reg558 <= {{{(reg555 ? reg546 : forvar525)}}};
                    end
                end
              for (forvar565 = (1'h0); (forvar565 < (2'h2)); forvar565 = (forvar565 + (1'h1)))
                begin
                  if ((~^$unsigned($unsigned($signed(forvar542)))))
                    begin
                      reg566 <= $unsigned((((reg553 * forvar555) - $unsigned(forvar555)) ?
                          $signed((forvar520 || reg552)) : (~|forvar550[(1'h1):(1'h1)])));
                      reg567 <= $unsigned((^~(^(+reg537))));
                    end
                  else
                    begin
                      reg566 <= $unsigned($signed(($unsigned(reg562) ?
                          reg562[(2'h3):(2'h3)] : $signed((8'ha3)))));
                      reg567 <= $signed(((reg556[(2'h2):(1'h1)] <= forvar520) ?
                          (^~reg542[(2'h2):(1'h1)]) : ($signed(reg552) ?
                              {reg554} : forvar519[(4'ha):(4'ha)])));
                      reg568 <= (^$unsigned(reg522));
                      reg569 <= $unsigned(forvar556[(4'hd):(4'hb)]);
                    end
                  for (forvar570 = (1'h0); (forvar570 < (1'h0)); forvar570 = (forvar570 + (1'h1)))
                    begin
                      reg571 <= {({$signed(forvar542)} >>> (~(forvar534 ?
                              forvar538 : reg558)))};
                      reg572 <= $signed((|{$signed(reg568)}));
                    end
                  if ($signed(((-$signed(reg567)) ?
                      ({forvar559} | (forvar528 ?
                          reg561 : reg540)) : (((8'hb9) << (8'ha9)) << forvar529))))
                    begin
                      reg573 <= (($signed((reg524 != (8'hb8))) ?
                              (~|(8'h9d)) : reg564[(3'h7):(3'h5)]) ?
                          ((reg555[(4'h8):(3'h7)] ^ $signed(reg551)) >= forvar538[(3'h7):(1'h0)]) : (~$signed($signed(reg564))));
                      reg574 <= reg556[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg573 <= (~|$unsigned(forvar555[(2'h2):(1'h1)]));
                      reg574 <= reg561[(4'ha):(1'h1)];
                      reg575 <= ($signed(({forvar559} ?
                              reg548[(3'h5):(1'h0)] : (reg572 <= reg535))) ?
                          reg524 : {forvar543});
                    end
                end
              if (reg531[(4'ha):(3'h6)])
                begin
                  for (forvar576 = (1'h0); (forvar576 < (2'h3)); forvar576 = (forvar576 + (1'h1)))
                    begin
                      reg577 <= (reg575 > (&(|$signed(forvar520))));
                      reg578 <= (~&{$signed($unsigned((8'h9d)))});
                    end
                end
              else
                begin
                  if ((({$signed((8'hba))} ^~ $unsigned(reg526)) > (-((8'ha0) ?
                      {forvar542} : $unsigned(forvar576)))))
                    begin
                      reg576 <= (reg546 ? reg562 : forvar554[(3'h7):(3'h6)]);
                      reg577 <= (((|(wire518 + reg541)) ?
                          reg561[(2'h2):(1'h0)] : {(forvar550 ?
                                  reg568 : (8'hb2))}) + (reg547 ?
                          (8'hb8) : (forvar559[(1'h0):(1'h0)] && (8'hb2))));
                    end
                  else
                    begin
                      reg576 <= reg533;
                    end
                  for (forvar578 = (1'h0); (forvar578 < (2'h2)); forvar578 = (forvar578 + (1'h1)))
                    begin
                      reg579 <= (^(~(&(forvar549 * forvar555))));
                      reg580 <= reg533[(3'h4):(3'h4)];
                    end
                end
            end
          for (forvar581 = (1'h0); (forvar581 < (2'h3)); forvar581 = (forvar581 + (1'h1)))
            begin
              reg582 <= reg554;
              if ((~&(8'hae)))
                begin
                  reg583 <= ($unsigned(reg541) >= $unsigned(forvar553[(2'h3):(1'h0)]));
                  if ($unsigned((((^forvar542) > $unsigned((8'hb9))) + ((reg535 ?
                          reg562 : reg524) ?
                      (reg540 ? reg556 : reg537) : (^forvar550)))))
                    begin
                      reg584 <= ($signed(reg545[(2'h2):(1'h1)]) ?
                          (reg582 >= $signed((~&forvar525))) : ({(forvar519 >> reg531)} ?
                              (~^((8'h9d) ?
                                  reg524 : forvar545)) : $unsigned((forvar534 >>> reg583))));
                      reg585 <= reg534;
                    end
                  else
                    begin
                      reg584 <= ($unsigned((reg576[(2'h3):(2'h3)] ?
                              forvar542[(3'h5):(1'h1)] : forvar542[(1'h0):(1'h0)])) ?
                          $unsigned($signed($unsigned(reg566))) : forvar570);
                      reg585 <= reg573[(4'hf):(3'h4)];
                      reg586 <= (-(8'hb4));
                    end
                end
              else
                begin
                  for (forvar583 = (1'h0); (forvar583 < (1'h1)); forvar583 = (forvar583 + (1'h1)))
                    begin
                      reg584 <= forvar581[(3'h4):(3'h4)];
                    end
                  if ((&(^~$signed((forvar555 <<< forvar534)))))
                    begin
                      reg585 <= (($unsigned((&forvar521)) >= $unsigned($unsigned(reg561))) ~^ $signed((^~$unsigned(reg524))));
                      reg586 <= ((reg522[(1'h1):(1'h1)] ?
                              ((^reg572) ?
                                  (forvar544 ?
                                      forvar553 : (8'h9e)) : (^~(8'hb6))) : (forvar549 ?
                                  (!(8'ha8)) : (reg572 ? reg565 : forvar554))) ?
                          {forvar529[(1'h1):(1'h1)]} : forvar545[(3'h6):(3'h4)]);
                    end
                  else
                    begin
                      reg585 <= {$signed((!(^~(8'hb4))))};
                      reg586 <= wire514[(2'h2):(1'h1)];
                      reg587 <= (reg527 | (!((reg548 ? forvar576 : forvar563) ?
                          (reg532 ?
                              forvar545 : reg538) : (forvar565 || forvar555))));
                      reg588 <= (~&(&{(forvar519 ? reg546 : (8'hb9))}));
                    end
                  if (reg555[(3'h6):(1'h0)])
                    begin
                      reg589 <= ((reg542[(3'h5):(2'h2)] ?
                          ({reg548} > $unsigned((8'hac))) : ($signed(reg586) ?
                              (reg542 ^ reg566) : {reg571})) <<< (reg527 < reg585));
                      reg590 <= $signed(forvar570[(3'h5):(3'h4)]);
                      reg591 <= ({(^~(reg567 ?
                              forvar538 : forvar570))} & reg527);
                      reg592 <= {wire517};
                    end
                  else
                    begin
                      reg589 <= (($signed($unsigned(forvar578)) ?
                          ($signed((8'hb4)) < $unsigned((8'hb0))) : (~(&reg565))) * (reg543[(3'h6):(1'h1)] ?
                          $signed((wire514 ? reg530 : reg538)) : (-{reg533})));
                      reg590 <= $signed($unsigned(((&reg556) ^~ {reg580})));
                      reg591 <= $unsigned($signed(((&(8'hb9)) ?
                          $signed(reg523) : forvar549[(2'h3):(1'h1)])));
                    end
                  for (forvar593 = (1'h0); (forvar593 < (1'h1)); forvar593 = (forvar593 + (1'h1)))
                    begin
                      reg594 <= (-(^(reg560 > (reg575 ^ (8'h9d)))));
                    end
                end
              for (forvar595 = (1'h0); (forvar595 < (1'h1)); forvar595 = (forvar595 + (1'h1)))
                begin
                  if (($signed(((&reg552) >> $unsigned(forvar576))) * $signed($signed($unsigned((8'ha5))))))
                    begin
                      reg596 <= (!($unsigned($signed(reg559)) < (!reg577[(3'h7):(3'h4)])));
                      reg597 <= forvar578[(2'h3):(1'h0)];
                      reg598 <= forvar570;
                      reg599 <= ((!($unsigned(wire517) - reg589)) ?
                          (reg562[(3'h4):(2'h2)] ?
                              ((reg571 < reg591) != $unsigned(forvar570)) : {(8'h9c)}) : ($signed(forvar525[(1'h0):(1'h0)]) - forvar570));
                    end
                  else
                    begin
                      reg596 <= forvar538;
                      reg597 <= {forvar559};
                      reg598 <= (^~$signed((|$unsigned(reg524))));
                    end
                  if ($unsigned((-(forvar570[(2'h2):(1'h1)] < (reg535 >= reg576)))))
                    begin
                      reg600 <= (^~$signed(forvar593));
                    end
                  else
                    begin
                      reg600 <= $signed((&wire517[(1'h0):(1'h0)]));
                    end
                end
              if (($signed(((reg569 - forvar543) << {forvar528})) >> $unsigned(reg535)))
                begin
                  reg601 <= (|reg575[(2'h2):(1'h0)]);
                  for (forvar602 = (1'h0); (forvar602 < (1'h0)); forvar602 = (forvar602 + (1'h1)))
                    begin
                      reg603 <= ((8'hb8) ? reg541 : reg590);
                      reg604 <= $unsigned(((forvar570[(3'h6):(2'h3)] || reg569[(3'h4):(2'h2)]) ?
                          (^$unsigned(forvar520)) : ({reg597} + $signed(reg566))));
                      reg605 <= (+$unsigned((|reg578[(3'h5):(2'h3)])));
                    end
                  if ((~^(~^(^~$signed(reg540)))))
                    begin
                      reg606 <= (~forvar556);
                      reg607 <= reg591;
                      reg608 <= $signed(((|$signed(reg531)) ?
                          $unsigned($unsigned(wire517)) : ($signed(reg565) == $signed(reg596))));
                      reg609 <= (reg582 || $signed(forvar544[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg606 <= ($unsigned($signed($unsigned(reg569))) ?
                          forvar539[(1'h0):(1'h0)] : reg546);
                      reg607 <= ($signed(forvar519[(1'h0):(1'h0)]) && (|$signed($signed(reg537))));
                      reg608 <= ($signed($signed($unsigned(reg601))) << {$signed({(8'had)})});
                    end
                  if (($signed($signed((~^(8'ha6)))) ?
                      $signed(reg539) : ($unsigned(reg531) ?
                          (&forvar553[(1'h0):(1'h0)]) : $unsigned(forvar534[(4'ha):(1'h0)]))))
                    begin
                      reg610 <= $unsigned(reg527[(4'ha):(3'h6)]);
                      reg611 <= ($signed(reg561[(2'h3):(1'h0)]) ?
                          $signed(reg587) : ({forvar593[(4'h8):(1'h0)]} <<< (~|(forvar550 ?
                              reg530 : (8'haa)))));
                      reg612 <= forvar554;
                      reg613 <= (forvar563 + $signed(reg538[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg610 <= (reg524[(1'h1):(1'h0)] ?
                          $unsigned((^(reg561 ? reg587 : reg572))) : reg536);
                      reg611 <= $signed($signed((forvar593[(3'h4):(2'h3)] & {reg542})));
                      reg612 <= $signed((reg554 ?
                          reg537[(4'h9):(1'h0)] : (reg559[(4'hc):(2'h3)] ?
                              forvar563[(2'h3):(2'h2)] : reg572[(3'h5):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar601 = (1'h0); (forvar601 < (2'h2)); forvar601 = (forvar601 + (1'h1)))
                    begin
                      reg602 <= (~|reg557);
                      reg603 <= reg553;
                    end
                  for (forvar604 = (1'h0); (forvar604 < (1'h1)); forvar604 = (forvar604 + (1'h1)))
                    begin
                      reg605 <= $signed($unsigned(reg539));
                    end
                end
            end
          for (forvar614 = (1'h0); (forvar614 < (1'h0)); forvar614 = (forvar614 + (1'h1)))
            begin
              for (forvar615 = (1'h0); (forvar615 < (1'h0)); forvar615 = (forvar615 + (1'h1)))
                begin
                  reg616 <= $signed($unsigned($unsigned((~&reg574))));
                  for (forvar617 = (1'h0); (forvar617 < (1'h0)); forvar617 = (forvar617 + (1'h1)))
                    begin
                      reg618 <= (forvar544[(1'h0):(1'h0)] >>> (reg527[(3'h5):(2'h2)] ?
                          $unsigned({reg616}) : (~&$signed(forvar576))));
                      reg619 <= reg563;
                      reg620 <= (({((8'hb8) > reg531)} ^~ ((forvar615 >= reg522) ?
                              (reg609 != reg548) : reg573[(3'h6):(1'h1)])) ?
                          reg572 : ({$signed((8'hb5))} ?
                              reg575 : $unsigned($unsigned(reg569))));
                    end
                end
              for (forvar621 = (1'h0); (forvar621 < (1'h0)); forvar621 = (forvar621 + (1'h1)))
                begin
                  for (forvar622 = (1'h0); (forvar622 < (2'h3)); forvar622 = (forvar622 + (1'h1)))
                    begin
                      reg623 <= $unsigned($signed(((+reg559) ?
                          {reg547} : (reg573 ? forvar576 : reg567))));
                      reg624 <= (&$unsigned((8'ha2)));
                      reg625 <= ((8'had) | (((^~reg598) && $signed(forvar529)) ^ (reg585[(3'h5):(1'h1)] ?
                          reg535[(3'h7):(1'h0)] : (reg538 ?
                              (8'haa) : forvar525))));
                    end
                end
              for (forvar626 = (1'h0); (forvar626 < (1'h0)); forvar626 = (forvar626 + (1'h1)))
                begin
                  for (forvar627 = (1'h0); (forvar627 < (1'h1)); forvar627 = (forvar627 + (1'h1)))
                    begin
                      reg628 <= reg605[(3'h4):(1'h1)];
                    end
                end
            end
          if ($signed((reg620 ?
              $signed((reg561 ~^ reg599)) : (((8'hb2) ? reg565 : forvar539) ?
                  (~&reg599) : $signed(reg534)))))
            begin
              if ((^((&forvar529) && (forvar538[(4'hd):(4'hb)] ?
                  forvar525[(3'h7):(2'h3)] : (reg572 ? reg600 : reg612)))))
                begin
                  for (forvar629 = (1'h0); (forvar629 < (2'h2)); forvar629 = (forvar629 + (1'h1)))
                    begin
                      reg630 <= $signed((~^reg539));
                    end
                  if ((reg623[(2'h2):(1'h0)] & (|{(reg552 ?
                          reg560 : forvar593)})))
                    begin
                      reg631 <= ((((forvar554 ?
                                  reg563 : reg601) >= (&forvar563)) ?
                              $signed(forvar525) : {$unsigned(reg562)}) ?
                          $signed((+$unsigned((8'ha8)))) : $signed(($unsigned(reg551) < (reg602 != reg607))));
                    end
                  else
                    begin
                      reg631 <= reg576;
                      reg632 <= reg567;
                    end
                  for (forvar633 = (1'h0); (forvar633 < (2'h2)); forvar633 = (forvar633 + (1'h1)))
                    begin
                      reg634 <= ((($unsigned(reg524) >= (~forvar617)) + (reg591[(2'h2):(2'h2)] ^~ $signed((8'hb3)))) ?
                          (!(+reg562)) : reg620);
                    end
                end
              else
                begin
                  for (forvar629 = (1'h0); (forvar629 < (2'h3)); forvar629 = (forvar629 + (1'h1)))
                    begin
                      reg630 <= reg530[(2'h3):(1'h1)];
                      reg631 <= $signed(reg567);
                    end
                end
              for (forvar635 = (1'h0); (forvar635 < (1'h0)); forvar635 = (forvar635 + (1'h1)))
                begin
                  for (forvar636 = (1'h0); (forvar636 < (2'h2)); forvar636 = (forvar636 + (1'h1)))
                    begin
                      reg637 <= reg591[(1'h1):(1'h0)];
                      reg638 <= $unsigned(reg559);
                    end
                  for (forvar639 = (1'h0); (forvar639 < (1'h0)); forvar639 = (forvar639 + (1'h1)))
                    begin
                      reg640 <= (+(((-reg591) >> reg558) ?
                          $signed(reg573[(3'h6):(2'h2)]) : (reg522 ?
                              ((8'hb0) ?
                                  (8'hb0) : reg553) : (reg565 + reg603))));
                    end
                  reg641 <= (8'hb3);
                  for (forvar642 = (1'h0); (forvar642 < (1'h0)); forvar642 = (forvar642 + (1'h1)))
                    begin
                      reg643 <= $signed((reg634 > wire516));
                      reg644 <= reg562;
                    end
                end
            end
          else
            begin
              if ($unsigned((8'ha8)))
                begin
                  for (forvar629 = (1'h0); (forvar629 < (2'h3)); forvar629 = (forvar629 + (1'h1)))
                    begin
                      reg630 <= $unsigned((!($unsigned((8'ha7)) ?
                          {reg565} : (8'ha7))));
                      reg631 <= {(8'h9c)};
                    end
                  for (forvar632 = (1'h0); (forvar632 < (1'h0)); forvar632 = (forvar632 + (1'h1)))
                    begin
                      reg633 <= {reg610[(1'h0):(1'h0)]};
                      reg634 <= (((reg605[(3'h4):(1'h0)] || (reg538 > reg588)) + $signed((wire515 ?
                          reg599 : (8'h9d)))) ^ reg625[(3'h7):(1'h1)]);
                      reg635 <= reg554[(3'h5):(3'h5)];
                      reg636 <= wire517[(3'h5):(3'h4)];
                    end
                end
              else
                begin
                  reg629 <= reg561;
                  for (forvar630 = (1'h0); (forvar630 < (1'h0)); forvar630 = (forvar630 + (1'h1)))
                    begin
                      reg631 <= ($unsigned($unsigned($unsigned((8'hb1)))) ?
                          reg602 : reg558);
                    end
                  if (forvar626[(1'h1):(1'h1)])
                    begin
                      reg632 <= (~|(($signed(reg579) <= forvar635) && reg613[(4'h9):(2'h3)]));
                      reg633 <= wire517;
                      reg634 <= ($signed($signed(forvar629[(3'h7):(3'h4)])) || (reg640[(1'h0):(1'h0)] || $unsigned({wire518})));
                    end
                  else
                    begin
                      reg632 <= reg526;
                    end
                  reg635 <= $unsigned((($signed(reg589) ?
                      (-reg598) : forvar626[(4'h9):(2'h2)]) <= $signed($signed(reg597))));
                end
            end
        end
      if (forvar554[(3'h5):(3'h5)])
        begin
          for (forvar645 = (1'h0); (forvar645 < (2'h2)); forvar645 = (forvar645 + (1'h1)))
            begin
              reg646 <= (((reg597[(1'h0):(1'h0)] + $signed(forvar529)) ?
                      forvar617 : ($unsigned((8'ha3)) ?
                          (|reg624) : (!reg638))) ?
                  (((reg538 || (8'hb9)) ?
                          reg601[(3'h7):(3'h5)] : $unsigned(forvar632)) ?
                      (~(wire514 ?
                          reg535 : forvar639)) : (!(~^reg588))) : reg588[(4'hb):(2'h3)]);
              for (forvar647 = (1'h0); (forvar647 < (1'h1)); forvar647 = (forvar647 + (1'h1)))
                begin
                  for (forvar648 = (1'h0); (forvar648 < (2'h3)); forvar648 = (forvar648 + (1'h1)))
                    begin
                      reg649 <= reg594;
                    end
                  if ($unsigned((|{reg597})))
                    begin
                      reg650 <= $unsigned((reg625 << {reg649[(1'h1):(1'h1)]}));
                      reg651 <= reg569;
                    end
                  else
                    begin
                      reg650 <= $unsigned($signed((8'hae)));
                      reg651 <= $unsigned({((forvar521 ? reg619 : forvar544) ?
                              $unsigned(reg583) : (reg620 ?
                                  reg537 : (8'hb4)))});
                      reg652 <= forvar538;
                    end
                  for (forvar653 = (1'h0); (forvar653 < (2'h3)); forvar653 = (forvar653 + (1'h1)))
                    begin
                      reg654 <= $signed((8'hb0));
                      reg655 <= $unsigned($unsigned(reg613[(2'h3):(2'h3)]));
                    end
                  reg656 <= reg567;
                end
              for (forvar657 = (1'h0); (forvar657 < (2'h2)); forvar657 = (forvar657 + (1'h1)))
                begin
                  for (forvar658 = (1'h0); (forvar658 < (1'h0)); forvar658 = (forvar658 + (1'h1)))
                    begin
                      reg659 <= ($unsigned($unsigned(reg557[(1'h1):(1'h1)])) + (8'ha4));
                      reg660 <= {$unsigned(forvar635[(4'hd):(3'h5)])};
                      reg661 <= $unsigned((8'hac));
                      reg662 <= $unsigned((reg561 <= $unsigned($signed(reg534))));
                    end
                  if (reg602)
                    begin
                      reg663 <= ({$signed(((8'ha2) ? reg545 : forvar604))} ?
                          $signed((reg566[(4'h9):(3'h5)] - reg577)) : ({forvar647[(3'h4):(2'h3)]} <<< $unsigned((~^reg560))));
                      reg664 <= (&(+{reg631[(2'h2):(1'h1)]}));
                      reg665 <= $unsigned(({(&forvar563)} ?
                          {{reg556}} : ({(8'had)} >= (8'ha4))));
                    end
                  else
                    begin
                      reg663 <= {((forvar539 >>> (forvar555 ?
                              reg537 : reg652)) & (8'hab))};
                      reg664 <= $unsigned($signed({{forvar629}}));
                      reg665 <= ($unsigned((8'ha1)) & reg569[(4'h9):(1'h0)]);
                      reg666 <= reg606;
                    end
                  if ($signed((forvar632 ?
                      (~reg624[(4'h8):(1'h1)]) : (reg540[(2'h3):(2'h2)] ?
                          (reg548 ? forvar556 : reg600) : (reg558 ?
                              (8'hae) : reg586)))))
                    begin
                      reg667 <= reg638;
                    end
                  else
                    begin
                      reg667 <= ((($signed(reg631) ?
                              (forvar647 ?
                                  reg603 : (8'hba)) : reg552[(2'h2):(1'h1)]) ?
                          forvar601[(2'h3):(2'h3)] : reg663[(1'h1):(1'h0)]) >>> (~|forvar617[(2'h2):(1'h0)]));
                    end
                end
              if (((reg636 ?
                  $unsigned((reg602 ~^ reg652)) : (reg613[(4'ha):(4'h9)] == $signed(reg611))) & ((reg583 | ((8'hac) ?
                      forvar633 : reg650)) ?
                  $signed({reg578}) : $signed((~|reg661)))))
                begin
                  for (forvar668 = (1'h0); (forvar668 < (2'h3)); forvar668 = (forvar668 + (1'h1)))
                    begin
                      reg669 <= (8'had);
                      reg670 <= (wire517[(4'hc):(4'h9)] ? reg663 : (8'hb4));
                    end
                  for (forvar671 = (1'h0); (forvar671 < (1'h0)); forvar671 = (forvar671 + (1'h1)))
                    begin
                      reg672 <= $unsigned($signed(reg524[(4'h9):(4'h9)]));
                      reg673 <= reg573;
                    end
                  for (forvar674 = (1'h0); (forvar674 < (2'h3)); forvar674 = (forvar674 + (1'h1)))
                    begin
                      reg675 <= (forvar521 ?
                          ({{reg660}} > reg574) : (reg554[(3'h6):(3'h5)] < forvar539));
                      reg676 <= $signed((&($unsigned(reg597) <<< (reg579 ?
                          reg612 : forvar639))));
                      reg677 <= reg656[(3'h6):(2'h3)];
                    end
                  if ((reg572[(1'h0):(1'h0)] ?
                      reg574[(4'h8):(3'h4)] : (!$unsigned((forvar555 ?
                          reg606 : forvar626)))))
                    begin
                      reg678 <= reg591;
                      reg679 <= (($unsigned(reg663[(3'h4):(2'h3)]) ?
                              forvar525[(2'h2):(1'h0)] : (8'hb8)) ?
                          (reg555[(4'h9):(1'h1)] ?
                              $unsigned($signed(reg640)) : {reg565[(1'h1):(1'h0)]}) : forvar534[(2'h3):(1'h0)]);
                      reg680 <= {reg602};
                      reg681 <= $signed($signed(forvar553[(4'hc):(4'hc)]));
                    end
                  else
                    begin
                      reg678 <= (8'hb3);
                    end
                end
              else
                begin
                  if (reg590)
                    begin
                      reg668 <= $unsigned(forvar668[(4'h8):(1'h0)]);
                    end
                  else
                    begin
                      reg668 <= reg616;
                      reg669 <= reg532;
                      reg670 <= $signed($unsigned((8'hba)));
                    end
                  for (forvar671 = (1'h0); (forvar671 < (1'h1)); forvar671 = (forvar671 + (1'h1)))
                    begin
                      reg672 <= $signed({$signed((reg589 ? reg677 : reg613))});
                      reg673 <= (reg608[(2'h2):(1'h1)] ^~ $signed(reg670[(2'h2):(1'h0)]));
                      reg674 <= reg598[(3'h6):(1'h0)];
                      reg675 <= {((-reg583[(4'he):(3'h7)]) ?
                              reg590[(3'h4):(1'h0)] : (-$unsigned(reg566)))};
                    end
                  for (forvar676 = (1'h0); (forvar676 < (2'h3)); forvar676 = (forvar676 + (1'h1)))
                    begin
                      reg677 <= {{(((8'hb0) ?
                                  forvar543 : (8'hb6)) >> {reg556})}};
                    end
                  for (forvar678 = (1'h0); (forvar678 < (1'h1)); forvar678 = (forvar678 + (1'h1)))
                    begin
                      reg679 <= reg573;
                      reg680 <= forvar602;
                      reg681 <= (({reg656} == $signed(forvar622)) >>> (forvar538 ?
                          (8'ha1) : (|(reg523 ? forvar555 : reg634))));
                    end
                end
            end
          reg682 <= forvar632;
          for (forvar683 = (1'h0); (forvar683 < (1'h0)); forvar683 = (forvar683 + (1'h1)))
            begin
              reg684 <= reg678;
            end
        end
      else
        begin
          reg645 <= forvar602;
          for (forvar646 = (1'h0); (forvar646 < (2'h3)); forvar646 = (forvar646 + (1'h1)))
            begin
              if ($signed((-((reg565 < reg651) ? forvar544 : reg668))))
                begin
                  reg647 <= ($unsigned((forvar627 - (forvar627 <<< reg660))) * ((forvar550[(4'hc):(3'h6)] <= (reg638 * forvar520)) ?
                      ($unsigned((8'ha3)) * {forvar648}) : $signed($signed(forvar578))));
                  for (forvar648 = (1'h0); (forvar648 < (1'h0)); forvar648 = (forvar648 + (1'h1)))
                    begin
                      reg649 <= ((^$signed($unsigned(forvar671))) ?
                          (|($unsigned(reg546) ?
                              ((8'ha2) & reg673) : reg523[(2'h2):(1'h0)])) : $signed((forvar555 < $signed(forvar545))));
                      reg650 <= reg582[(3'h5):(1'h1)];
                      reg651 <= reg524[(4'h9):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar647 = (1'h0); (forvar647 < (2'h2)); forvar647 = (forvar647 + (1'h1)))
                    begin
                      reg648 <= (^~$unsigned((8'hb7)));
                      reg649 <= (($unsigned((forvar555 + reg551)) << (reg553 < $unsigned((8'h9e)))) ?
                          ({(forvar636 ? (8'ha6) : forvar534)} ?
                              forvar629[(1'h1):(1'h1)] : $unsigned((reg523 ?
                                  reg599 : reg625))) : reg536[(2'h3):(2'h3)]);
                      reg650 <= (forvar519 * (~|forvar614[(3'h6):(3'h6)]));
                    end
                  for (forvar651 = (1'h0); (forvar651 < (1'h1)); forvar651 = (forvar651 + (1'h1)))
                    begin
                      reg652 <= $signed((($unsigned(reg597) <= $signed((8'ha9))) ?
                          $unsigned(reg585[(1'h1):(1'h1)]) : ($unsigned(forvar632) ~^ $unsigned(forvar534))));
                      reg653 <= (~|($unsigned((reg682 << reg651)) || {forvar617[(3'h4):(1'h1)]}));
                      reg654 <= $unsigned(reg603);
                      reg655 <= reg630;
                    end
                  if ((|(((reg679 + (8'ha7)) ?
                          $unsigned(reg606) : $signed(forvar534)) ?
                      {$signed(forvar550)} : (&(~reg580)))))
                    begin
                      reg656 <= (|reg668);
                      reg657 <= reg661;
                      reg658 <= ((+{(reg588 ? reg577 : (8'haf))}) ?
                          ($unsigned($unsigned(reg587)) ?
                              ({forvar539} * $signed(wire517)) : $signed({reg667})) : reg539);
                      reg659 <= forvar657[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg656 <= $unsigned(wire514[(2'h3):(1'h0)]);
                      reg657 <= (+reg576[(4'ha):(3'h6)]);
                      reg658 <= $signed($signed((-{forvar658})));
                      reg659 <= $signed((&(~|(reg586 >= reg650))));
                    end
                  for (forvar660 = (1'h0); (forvar660 < (2'h2)); forvar660 = (forvar660 + (1'h1)))
                    begin
                      reg661 <= reg522[(2'h2):(1'h0)];
                      reg662 <= $unsigned(reg658);
                    end
                end
            end
          if ((&$unsigned(($signed(wire515) ?
              (reg530 ? (8'ha6) : (8'ha0)) : (reg665 & (8'hac))))))
            begin
              for (forvar663 = (1'h0); (forvar663 < (1'h0)); forvar663 = (forvar663 + (1'h1)))
                begin
                  if ($unsigned(forvar519[(4'hf):(2'h3)]))
                    begin
                      reg664 <= reg604[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg664 <= {{forvar617}};
                      reg665 <= reg591;
                      reg666 <= $unsigned($signed($signed((reg562 << forvar565))));
                      reg667 <= (+(8'ha4));
                    end
                end
            end
          else
            begin
              for (forvar663 = (1'h0); (forvar663 < (2'h3)); forvar663 = (forvar663 + (1'h1)))
                begin
                  for (forvar664 = (1'h0); (forvar664 < (2'h2)); forvar664 = (forvar664 + (1'h1)))
                    begin
                      reg665 <= (((reg541 ?
                                  $signed(reg670) : (forvar627 ?
                                      reg636 : reg646)) ?
                              {reg579} : wire515) ?
                          reg583[(2'h3):(2'h2)] : $signed($signed((reg644 ?
                              reg576 : forvar629))));
                      reg666 <= $signed((^({reg650} ?
                          $unsigned(forvar653) : forvar664[(4'h9):(2'h3)])));
                    end
                  reg667 <= reg548[(1'h0):(1'h0)];
                end
              for (forvar668 = (1'h0); (forvar668 < (1'h1)); forvar668 = (forvar668 + (1'h1)))
                begin
                  reg669 <= $signed($unsigned(((forvar647 != (8'hb3)) ?
                      (forvar636 + forvar576) : forvar520)));
                end
              if ($signed($signed(({reg628} ?
                  (reg532 ? forvar627 : reg588) : $unsigned(reg562)))))
                begin
                  reg670 <= (-reg578[(4'h9):(4'h9)]);
                  if ($signed((forvar550 ?
                      $unsigned((reg675 ?
                          forvar639 : reg583)) : forvar668[(3'h4):(1'h1)])))
                    begin
                      reg671 <= {$signed(((forvar554 | forvar538) ?
                              $signed(forvar648) : $signed(forvar651)))};
                      reg672 <= ((reg640[(2'h3):(1'h0)] ?
                              reg647[(1'h0):(1'h0)] : $unsigned((reg584 - (8'ha3)))) ?
                          (|$unsigned(((8'h9f) > forvar678))) : reg663[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg671 <= (^$signed($unsigned($signed((8'hb0)))));
                      reg672 <= (forvar645[(4'hc):(2'h2)] || (~|reg666[(3'h4):(3'h4)]));
                      reg673 <= (+($signed($unsigned(forvar671)) ?
                          ((!reg573) ?
                              wire514[(3'h4):(2'h3)] : {reg610}) : reg670[(1'h1):(1'h1)]));
                      reg674 <= (~^(|(8'hb4)));
                    end
                  if ((reg530[(3'h6):(1'h1)] == (-$unsigned((8'hab)))))
                    begin
                      reg675 <= forvar647;
                      reg676 <= $unsigned((&{reg589[(1'h0):(1'h0)]}));
                      reg677 <= ((+forvar556) ?
                          $signed((~$signed(forvar565))) : ($unsigned(((8'ha2) ?
                                  forvar581 : (8'ha4))) ?
                              ($signed(reg612) + {reg575}) : reg643[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg675 <= (forvar651 >> ($signed((forvar676 & reg567)) ?
                          ((reg607 ~^ reg657) ?
                              (-reg551) : $unsigned(reg616)) : $unsigned($signed(forvar653))));
                      reg676 <= (reg684 ?
                          $signed(($unsigned(forvar648) && {reg657})) : $signed(((8'haf) ?
                              $signed((8'h9e)) : ((8'ha7) ?
                                  forvar678 : reg585))));
                      reg677 <= reg637;
                    end
                end
              else
                begin
                  for (forvar670 = (1'h0); (forvar670 < (1'h0)); forvar670 = (forvar670 + (1'h1)))
                    begin
                      reg671 <= reg638;
                    end
                  for (forvar672 = (1'h0); (forvar672 < (2'h3)); forvar672 = (forvar672 + (1'h1)))
                    begin
                      reg673 <= reg589[(3'h7):(2'h3)];
                    end
                  for (forvar674 = (1'h0); (forvar674 < (2'h3)); forvar674 = (forvar674 + (1'h1)))
                    begin
                      reg675 <= $signed(({reg640} ?
                          reg646 : ($unsigned(reg654) ?
                              (reg566 ?
                                  (8'hac) : reg548) : $unsigned(reg629))));
                      reg676 <= reg572;
                    end
                  for (forvar677 = (1'h0); (forvar677 < (2'h3)); forvar677 = (forvar677 + (1'h1)))
                    begin
                      reg678 <= forvar595;
                      reg679 <= $unsigned(forvar525[(3'h4):(1'h0)]);
                      reg680 <= reg659;
                    end
                end
              if (reg602)
                begin
                  for (forvar681 = (1'h0); (forvar681 < (1'h0)); forvar681 = (forvar681 + (1'h1)))
                    begin
                      reg682 <= reg619;
                      reg683 <= $signed(($signed(((8'ha0) >>> (8'had))) && forvar663));
                      reg684 <= $unsigned($unsigned($signed(forvar676)));
                      reg685 <= ({$unsigned((forvar651 <<< reg532))} <<< (8'ha2));
                    end
                  for (forvar686 = (1'h0); (forvar686 < (1'h0)); forvar686 = (forvar686 + (1'h1)))
                    begin
                      reg687 <= forvar595;
                      reg688 <= ((reg683[(1'h0):(1'h0)] ?
                          reg638[(2'h3):(1'h1)] : (reg579[(2'h2):(2'h2)] && {reg578})) ^~ $unsigned(((reg598 >= forvar630) >> $signed(reg632))));
                      reg689 <= $unsigned($signed((&{(8'h9f)})));
                    end
                  reg690 <= {(8'hb1)};
                  if ($unsigned(reg647[(4'h8):(3'h4)]))
                    begin
                      reg691 <= {(reg690 ?
                              reg539[(1'h1):(1'h1)] : $signed(reg590))};
                      reg692 <= $unsigned($unsigned($signed(forvar645)));
                      reg693 <= forvar647[(3'h5):(1'h0)];
                    end
                  else
                    begin
                      reg691 <= (^(((forvar658 ? reg673 : (8'ha0)) ?
                              (~&(8'haa)) : {reg533}) ?
                          {reg532} : $signed(reg693)));
                    end
                end
              else
                begin
                  for (forvar681 = (1'h0); (forvar681 < (2'h2)); forvar681 = (forvar681 + (1'h1)))
                    begin
                      reg682 <= $signed($signed(((^reg678) ?
                          $unsigned(forvar576) : forvar630[(4'h9):(3'h6)])));
                      reg683 <= $unsigned(reg672[(4'h9):(2'h3)]);
                    end
                  reg684 <= ({reg596[(3'h5):(1'h0)]} ?
                      {((reg675 ?
                              reg576 : reg648) || reg559[(4'h8):(3'h4)])} : (|(^~$signed(reg628))));
                  reg685 <= $unsigned((^~$signed($unsigned(reg573))));
                end
            end
          if ((~^$signed(reg524)))
            begin
              for (forvar694 = (1'h0); (forvar694 < (2'h3)); forvar694 = (forvar694 + (1'h1)))
                begin
                  if ($signed(($signed((reg655 ? reg646 : reg648)) ?
                      (forvar647[(4'hc):(3'h7)] ?
                          $unsigned(reg636) : ((8'ha9) ?
                              forvar520 : (8'hb9))) : (!$unsigned(reg645)))))
                    begin
                      reg695 <= $signed(($unsigned({reg548}) ?
                          (~&(forvar593 <<< reg541)) : ((forvar683 ?
                              reg543 : forvar542) + (!forvar565))));
                      reg696 <= reg536[(3'h4):(1'h1)];
                      reg697 <= $unsigned(($unsigned((^wire517)) ?
                          ($unsigned(reg602) ?
                              $unsigned(forvar556) : (forvar615 ?
                                  forvar651 : reg580)) : $unsigned((|reg535))));
                    end
                  else
                    begin
                      reg695 <= {reg678};
                      reg696 <= reg599;
                      reg697 <= $signed(((8'hac) ^ (reg556 ?
                          (reg599 ? (8'hb9) : forvar639) : reg568)));
                    end
                  if (($unsigned((!$unsigned(forvar544))) ?
                      $unsigned((^{reg654})) : (~reg658[(2'h2):(2'h2)])))
                    begin
                      reg698 <= ({$signed(reg633)} ?
                          ((forvar539 ?
                                  (forvar539 ^ reg648) : $signed(forvar615)) ?
                              forvar629[(4'hf):(4'h8)] : $unsigned($unsigned(reg656))) : reg650);
                      reg699 <= ($signed((~|reg571)) ?
                          $signed(reg612) : reg608);
                    end
                  else
                    begin
                      reg698 <= $signed(reg690[(4'hb):(3'h6)]);
                      reg699 <= reg524[(1'h0):(1'h0)];
                    end
                end
              reg700 <= reg693;
              for (forvar701 = (1'h0); (forvar701 < (1'h0)); forvar701 = (forvar701 + (1'h1)))
                begin
                  if (reg547)
                    begin
                      reg702 <= $unsigned({((8'ha3) >= $signed(reg628))});
                      reg703 <= $unsigned(reg567[(4'h8):(4'h8)]);
                    end
                  else
                    begin
                      reg702 <= (reg603 ?
                          $unsigned((+reg623)) : (!((reg576 | forvar528) ?
                              (forvar545 + reg548) : reg663)));
                      reg703 <= (reg558 ?
                          $signed((reg523[(1'h0):(1'h0)] ?
                              ((8'ha7) ?
                                  reg531 : forvar604) : (-(8'hae)))) : $unsigned(((~|(8'hab)) && $unsigned(reg535))));
                      reg704 <= wire514;
                    end
                  for (forvar705 = (1'h0); (forvar705 < (2'h2)); forvar705 = (forvar705 + (1'h1)))
                    begin
                      reg706 <= (-($unsigned($signed(forvar553)) ?
                          ($signed(reg527) ?
                              reg693 : reg607) : (!$unsigned(reg568))));
                      reg707 <= reg649;
                      reg708 <= (8'hb0);
                    end
                  if ((+reg645))
                    begin
                      reg709 <= (reg662[(2'h3):(1'h1)] | (($unsigned((8'hb1)) << $signed(reg661)) ?
                          $unsigned(((8'ha6) || (8'haa))) : (reg579 ?
                              $unsigned(reg649) : $signed(reg693))));
                      reg710 <= {$signed(($signed(forvar604) ?
                              (8'ha8) : {reg558}))};
                      reg711 <= $unsigned($signed((~{forvar621})));
                      reg712 <= {(&(~&(~|(8'hb2))))};
                    end
                  else
                    begin
                      reg709 <= ($signed((((8'ha5) ?
                              reg524 : reg531) <= (reg711 ^~ (8'ha7)))) ?
                          $unsigned($unsigned(forvar648[(1'h1):(1'h1)])) : $signed(($signed((8'hb9)) < (|reg556))));
                    end
                end
            end
          else
            begin
              for (forvar694 = (1'h0); (forvar694 < (1'h1)); forvar694 = (forvar694 + (1'h1)))
                begin
                  for (forvar695 = (1'h0); (forvar695 < (1'h1)); forvar695 = (forvar695 + (1'h1)))
                    begin
                      reg696 <= $unsigned((($unsigned(reg660) + {reg661}) ?
                          ($signed((8'hb9)) <= (|reg562)) : (&reg541[(4'ha):(2'h3)])));
                      reg697 <= $unsigned(((-(reg576 ?
                          reg522 : (8'ha5))) ^ reg630));
                      reg698 <= $signed({$unsigned((~(8'ha8)))});
                    end
                  reg699 <= ({$unsigned({(8'h9f)})} & $signed($unsigned(reg636[(1'h1):(1'h1)])));
                  for (forvar700 = (1'h0); (forvar700 < (2'h2)); forvar700 = (forvar700 + (1'h1)))
                    begin
                      reg701 <= $unsigned(forvar646);
                      reg702 <= $signed($signed(reg530));
                      reg703 <= (reg649 * reg685);
                      reg704 <= (+(|($unsigned(reg692) < (forvar642 | forvar694))));
                    end
                end
              for (forvar705 = (1'h0); (forvar705 < (1'h1)); forvar705 = (forvar705 + (1'h1)))
                begin
                  if ((8'hab))
                    begin
                      reg706 <= reg685[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg706 <= $unsigned({((reg677 ?
                              forvar559 : reg681) != $unsigned(reg629))});
                      reg707 <= $signed((forvar542[(3'h6):(3'h4)] ^~ $unsigned($unsigned(forvar700))));
                    end
                  reg708 <= reg671[(4'hb):(3'h7)];
                end
              for (forvar709 = (1'h0); (forvar709 < (2'h2)); forvar709 = (forvar709 + (1'h1)))
                begin
                  for (forvar710 = (1'h0); (forvar710 < (1'h0)); forvar710 = (forvar710 + (1'h1)))
                    begin
                      reg711 <= ($signed($signed((reg530 << reg611))) ?
                          (&reg578[(4'he):(3'h4)]) : (((^~reg590) ?
                                  forvar646[(1'h0):(1'h0)] : $signed(reg660)) ?
                              reg546 : $unsigned({reg700})));
                      reg712 <= (8'hb6);
                      reg713 <= forvar651[(4'hc):(3'h5)];
                      reg714 <= {($signed((reg556 ?
                              reg555 : (8'ha5))) ^~ ($unsigned((8'ha0)) ?
                              reg641[(1'h0):(1'h0)] : $signed(forvar544)))};
                    end
                end
            end
        end
    end
  assign wire715 = $signed(reg714);
  assign wire716 = $signed($unsigned($unsigned((^reg706))));
  assign wire717 = (-reg605);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2034  (y, clk, wire2038, wire2037, wire2036, wire2035);
  output wire [(32'h5e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire2038;
  input wire signed [(4'h8):(1'h0)] wire2037;
  input wire [(4'hc):(1'h0)] wire2036;
  input wire [(3'h5):(1'h0)] wire2035;
  wire signed [(4'he):(1'h0)] wire3424;
  wire signed [(4'hd):(1'h0)] wire3423;
  wire [(5'h10):(1'h0)] wire3422;
  wire signed [(4'ha):(1'h0)] wire3421;
  wire [(4'hd):(1'h0)] wire3420;
  wire [(2'h2):(1'h0)] wire3419;
  wire signed [(2'h3):(1'h0)] wire3417;
  wire signed [(4'h8):(1'h0)] wire3044;
  wire signed [(4'he):(1'h0)] wire3042;
  assign y = {wire3424,
                 wire3423,
                 wire3422,
                 wire3421,
                 wire3420,
                 wire3419,
                 wire3417,
                 wire3044,
                 wire3042,
                 (1'h0)};
  module2039 #() modinst3043 (wire3042, clk, wire2035, wire2038, wire2036, wire2037, (8'ha0));
  assign wire3044 = ({wire2037[(3'h4):(2'h3)]} ?
                        ((^~(&wire2035)) ?
                            wire2035 : (wire2036 ^ $unsigned((8'hb1)))) : $unsigned((~&$signed((8'hb5)))));
  module3045 #() modinst3418 (wire3417, clk, wire3044, wire3042, wire2037, wire2035);
  assign wire3419 = ((^(!(wire3044 >= wire3044))) >= wire2035);
  assign wire3420 = wire3419[(2'h2):(2'h2)];
  assign wire3421 = {wire3417};
  assign wire3422 = ($unsigned((wire3042 * wire3042)) ?
                        ($unsigned(wire2036[(2'h3):(2'h2)]) >= {wire3419[(2'h2):(2'h2)]}) : wire3042[(4'h9):(2'h2)]);
  assign wire3423 = ($unsigned(({wire3421} != $unsigned(wire3417))) ?
                        wire2035[(3'h4):(3'h4)] : $signed(wire3422[(3'h5):(2'h3)]));
  assign wire3424 = ((wire3421[(1'h0):(1'h0)] ?
                            $unsigned($unsigned(wire2038)) : wire3422) ?
                        (~&wire3417) : (~^wire2036[(4'h9):(3'h6)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module867
#(parameter param2030 = (&(~&({(8'hb8)} ? ((8'hb6) ? (8'hb6) : (8'ha7)) : {(8'hb3)}))))
(y, clk, wire871, wire870, wire869, wire868);
  output wire [(32'h6cd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire871;
  input wire signed [(2'h3):(1'h0)] wire870;
  input wire signed [(5'h10):(1'h0)] wire869;
  input wire signed [(4'hb):(1'h0)] wire868;
  wire signed [(4'hc):(1'h0)] wire1972;
  wire [(2'h2):(1'h0)] wire1971;
  wire [(4'hd):(1'h0)] wire1969;
  wire signed [(5'h10):(1'h0)] wire979;
  wire [(3'h6):(1'h0)] wire978;
  wire signed [(3'h7):(1'h0)] wire977;
  wire signed [(2'h3):(1'h0)] wire951;
  wire [(3'h5):(1'h0)] wire950;
  wire signed [(4'h9):(1'h0)] wire873;
  wire [(4'hd):(1'h0)] wire872;
  reg signed [(5'h10):(1'h0)] reg2016 = (1'h0);
  reg [(3'h4):(1'h0)] reg2029 = (1'h0);
  reg [(4'hb):(1'h0)] reg2028 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2027 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2025 = (1'h0);
  reg [(4'hb):(1'h0)] reg2023 = (1'h0);
  reg [(4'hf):(1'h0)] reg2022 = (1'h0);
  reg [(3'h7):(1'h0)] reg2021 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2019 = (1'h0);
  reg [(5'h10):(1'h0)] reg2018 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2017 = (1'h0);
  reg [(4'hd):(1'h0)] reg2010 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2013 = (1'h0);
  reg [(4'hc):(1'h0)] reg2012 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2011 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2009 = (1'h0);
  reg [(4'he):(1'h0)] reg2007 = (1'h0);
  reg [(4'hb):(1'h0)] reg2006 = (1'h0);
  reg [(4'he):(1'h0)] reg2004 = (1'h0);
  reg [(3'h6):(1'h0)] reg2003 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2002 = (1'h0);
  reg [(3'h6):(1'h0)] reg2001 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2000 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1999 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1998 = (1'h0);
  reg [(4'hd):(1'h0)] reg1997 = (1'h0);
  reg [(4'hd):(1'h0)] reg1996 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1994 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1993 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1991 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1990 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1989 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1987 = (1'h0);
  reg [(5'h10):(1'h0)] reg1984 = (1'h0);
  reg [(3'h6):(1'h0)] reg1983 = (1'h0);
  reg [(4'hd):(1'h0)] reg1982 = (1'h0);
  reg [(3'h5):(1'h0)] reg1981 = (1'h0);
  reg [(3'h4):(1'h0)] reg1980 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1978 = (1'h0);
  reg [(2'h2):(1'h0)] reg1977 = (1'h0);
  reg [(4'hc):(1'h0)] reg876 = (1'h0);
  reg [(4'h8):(1'h0)] reg877 = (1'h0);
  reg [(4'hb):(1'h0)] reg878 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg880 = (1'h0);
  reg [(4'h8):(1'h0)] reg881 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg882 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg879 = (1'h0);
  reg [(3'h5):(1'h0)] reg883 = (1'h0);
  reg [(4'hb):(1'h0)] reg884 = (1'h0);
  reg [(3'h4):(1'h0)] reg886 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg887 = (1'h0);
  reg [(4'hf):(1'h0)] reg888 = (1'h0);
  reg [(3'h4):(1'h0)] reg889 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg891 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg892 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg893 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg894 = (1'h0);
  reg [(3'h6):(1'h0)] reg896 = (1'h0);
  reg signed [(4'he):(1'h0)] reg897 = (1'h0);
  reg [(4'hd):(1'h0)] reg898 = (1'h0);
  reg [(3'h4):(1'h0)] reg899 = (1'h0);
  reg [(4'hd):(1'h0)] reg900 = (1'h0);
  reg [(4'hb):(1'h0)] reg885 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg902 = (1'h0);
  reg [(3'h5):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg904 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg906 = (1'h0);
  reg [(2'h3):(1'h0)] reg905 = (1'h0);
  reg [(4'hb):(1'h0)] reg907 = (1'h0);
  reg [(4'h8):(1'h0)] reg908 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg909 = (1'h0);
  reg [(4'h8):(1'h0)] reg910 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg911 = (1'h0);
  reg [(3'h4):(1'h0)] reg912 = (1'h0);
  reg [(4'he):(1'h0)] reg914 = (1'h0);
  reg [(2'h2):(1'h0)] reg915 = (1'h0);
  reg [(2'h2):(1'h0)] reg916 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg917 = (1'h0);
  reg [(4'h8):(1'h0)] reg919 = (1'h0);
  reg [(2'h3):(1'h0)] reg920 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg921 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg923 = (1'h0);
  reg [(5'h10):(1'h0)] reg924 = (1'h0);
  reg [(4'hc):(1'h0)] reg925 = (1'h0);
  reg [(4'hf):(1'h0)] reg926 = (1'h0);
  reg [(3'h7):(1'h0)] reg927 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg922 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg928 = (1'h0);
  reg [(4'hb):(1'h0)] reg930 = (1'h0);
  reg [(3'h4):(1'h0)] reg931 = (1'h0);
  reg [(4'hd):(1'h0)] reg932 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg929 = (1'h0);
  reg [(4'ha):(1'h0)] reg933 = (1'h0);
  reg [(4'ha):(1'h0)] reg934 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg935 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg936 = (1'h0);
  reg [(4'hb):(1'h0)] reg937 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg938 = (1'h0);
  reg [(2'h3):(1'h0)] reg939 = (1'h0);
  reg [(3'h6):(1'h0)] reg940 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg941 = (1'h0);
  reg [(2'h2):(1'h0)] reg942 = (1'h0);
  reg [(4'hf):(1'h0)] reg943 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg944 = (1'h0);
  reg [(4'hf):(1'h0)] reg945 = (1'h0);
  reg signed [(4'he):(1'h0)] reg946 = (1'h0);
  reg [(2'h3):(1'h0)] reg947 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg949 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg953 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg954 = (1'h0);
  reg [(4'he):(1'h0)] reg955 = (1'h0);
  reg [(4'hf):(1'h0)] reg956 = (1'h0);
  reg [(4'ha):(1'h0)] reg958 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg960 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg961 = (1'h0);
  reg [(5'h10):(1'h0)] reg962 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg963 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg957 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg959 = (1'h0);
  reg [(4'h9):(1'h0)] reg964 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg966 = (1'h0);
  reg [(4'ha):(1'h0)] reg967 = (1'h0);
  reg [(4'hb):(1'h0)] reg968 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg969 = (1'h0);
  reg [(4'h8):(1'h0)] reg970 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg965 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg972 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg973 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg974 = (1'h0);
  reg [(4'hb):(1'h0)] reg975 = (1'h0);
  reg [(3'h5):(1'h0)] reg976 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2026 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2024 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2020 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2016 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2015 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2014 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2010 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2008 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1998 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2005 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1995 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1992 = (1'h0);
  reg [(4'he):(1'h0)] forvar1988 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1986 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1985 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1979 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1976 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1975 = (1'h0);
  reg [(4'he):(1'h0)] forvar1974 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1973 = (1'h0);
  reg [(5'h10):(1'h0)] forvar971 = (1'h0);
  reg [(4'hb):(1'h0)] forvar965 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar959 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar957 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar952 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar948 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar942 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar929 = (1'h0);
  reg [(4'h9):(1'h0)] forvar924 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar920 = (1'h0);
  reg [(4'hd):(1'h0)] forvar922 = (1'h0);
  reg [(5'h10):(1'h0)] forvar918 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar913 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar906 = (1'h0);
  reg [(2'h2):(1'h0)] forvar905 = (1'h0);
  reg [(4'he):(1'h0)] forvar901 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar880 = (1'h0);
  reg [(2'h2):(1'h0)] forvar895 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar890 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar885 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar881 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar879 = (1'h0);
  reg [(4'he):(1'h0)] forvar875 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar874 = (1'h0);
  assign y = {wire1972,
                 wire1971,
                 wire1969,
                 wire979,
                 wire978,
                 wire977,
                 wire951,
                 wire950,
                 wire873,
                 wire872,
                 reg2016,
                 reg2029,
                 reg2028,
                 reg2027,
                 reg2025,
                 reg2023,
                 reg2022,
                 reg2021,
                 reg2019,
                 reg2018,
                 reg2017,
                 reg2010,
                 reg2013,
                 reg2012,
                 reg2011,
                 reg2009,
                 reg2007,
                 reg2006,
                 reg2004,
                 reg2003,
                 reg2002,
                 reg2001,
                 reg2000,
                 reg1999,
                 reg1998,
                 reg1997,
                 reg1996,
                 reg1994,
                 reg1993,
                 reg1991,
                 reg1990,
                 reg1989,
                 reg1987,
                 reg1984,
                 reg1983,
                 reg1982,
                 reg1981,
                 reg1980,
                 reg1978,
                 reg1977,
                 reg876,
                 reg877,
                 reg878,
                 reg880,
                 reg881,
                 reg882,
                 reg879,
                 reg883,
                 reg884,
                 reg886,
                 reg887,
                 reg888,
                 reg889,
                 reg891,
                 reg892,
                 reg893,
                 reg894,
                 reg896,
                 reg897,
                 reg898,
                 reg899,
                 reg900,
                 reg885,
                 reg902,
                 reg903,
                 reg904,
                 reg906,
                 reg905,
                 reg907,
                 reg908,
                 reg909,
                 reg910,
                 reg911,
                 reg912,
                 reg914,
                 reg915,
                 reg916,
                 reg917,
                 reg919,
                 reg920,
                 reg921,
                 reg923,
                 reg924,
                 reg925,
                 reg926,
                 reg927,
                 reg922,
                 reg928,
                 reg930,
                 reg931,
                 reg932,
                 reg929,
                 reg933,
                 reg934,
                 reg935,
                 reg936,
                 reg937,
                 reg938,
                 reg939,
                 reg940,
                 reg941,
                 reg942,
                 reg943,
                 reg944,
                 reg945,
                 reg946,
                 reg947,
                 reg949,
                 reg953,
                 reg954,
                 reg955,
                 reg956,
                 reg958,
                 reg960,
                 reg961,
                 reg962,
                 reg963,
                 reg957,
                 reg959,
                 reg964,
                 reg966,
                 reg967,
                 reg968,
                 reg969,
                 reg970,
                 reg965,
                 reg972,
                 reg973,
                 reg974,
                 reg975,
                 reg976,
                 forvar2026,
                 forvar2024,
                 forvar2020,
                 forvar2016,
                 forvar2015,
                 forvar2014,
                 forvar2010,
                 forvar2008,
                 forvar1998,
                 forvar2005,
                 forvar1995,
                 forvar1992,
                 forvar1988,
                 forvar1986,
                 forvar1985,
                 forvar1979,
                 forvar1976,
                 forvar1975,
                 forvar1974,
                 forvar1973,
                 forvar971,
                 forvar965,
                 forvar959,
                 forvar957,
                 forvar952,
                 forvar948,
                 forvar942,
                 forvar929,
                 forvar924,
                 forvar920,
                 forvar922,
                 forvar918,
                 forvar913,
                 forvar906,
                 forvar905,
                 forvar901,
                 forvar880,
                 forvar895,
                 forvar890,
                 forvar885,
                 forvar881,
                 forvar879,
                 forvar875,
                 forvar874,
                 (1'h0)};
  assign wire872 = wire871;
  assign wire873 = wire872;
  always
    @(posedge clk) begin
      for (forvar874 = (1'h0); (forvar874 < (2'h3)); forvar874 = (forvar874 + (1'h1)))
        begin
          for (forvar875 = (1'h0); (forvar875 < (1'h0)); forvar875 = (forvar875 + (1'h1)))
            begin
              reg876 <= wire871[(3'h5):(3'h5)];
            end
          if ($signed($signed({(^wire871)})))
            begin
              if ($unsigned(forvar875))
                begin
                  if ((8'hb5))
                    begin
                      reg877 <= wire870;
                      reg878 <= {(!$unsigned((wire868 ? forvar875 : wire870)))};
                    end
                  else
                    begin
                      reg877 <= ($unsigned(forvar875) ?
                          $signed($unsigned($signed(forvar875))) : $signed((8'ha3)));
                      reg878 <= ($signed((&(wire869 ^ wire873))) ?
                          wire868[(3'h5):(3'h4)] : (reg878 ?
                              ((&wire870) + (forvar874 + wire869)) : reg878[(4'h9):(3'h6)]));
                    end
                  for (forvar879 = (1'h0); (forvar879 < (2'h3)); forvar879 = (forvar879 + (1'h1)))
                    begin
                      reg880 <= wire869[(4'hb):(4'hb)];
                      reg881 <= reg880[(3'h7):(3'h6)];
                      reg882 <= wire871;
                    end
                end
              else
                begin
                  reg877 <= ($unsigned((&(8'hba))) ?
                      {((wire870 << reg880) ?
                              forvar875 : $unsigned(wire871))} : ((reg880 ?
                              reg877[(1'h0):(1'h0)] : (-reg881)) ?
                          $signed(wire872) : (&(reg876 < wire873))));
                  if (wire870)
                    begin
                      reg878 <= forvar875[(2'h3):(1'h1)];
                      reg879 <= (reg878 == ($signed((wire868 & reg877)) ?
                          reg882 : reg880[(4'ha):(1'h1)]));
                      reg880 <= wire869[(4'h9):(1'h0)];
                    end
                  else
                    begin
                      reg878 <= (^~(wire869 & reg882));
                      reg879 <= ($signed($unsigned($signed(wire869))) || (-{wire871[(2'h2):(2'h2)]}));
                    end
                  for (forvar881 = (1'h0); (forvar881 < (1'h0)); forvar881 = (forvar881 + (1'h1)))
                    begin
                      reg882 <= forvar874;
                      reg883 <= $unsigned(reg881[(3'h6):(3'h5)]);
                    end
                end
              if (($unsigned($unsigned((reg881 < (8'hb0)))) ?
                  reg880 : $signed(reg879[(2'h3):(1'h0)])))
                begin
                  reg884 <= (!(8'h9d));
                  for (forvar885 = (1'h0); (forvar885 < (2'h3)); forvar885 = (forvar885 + (1'h1)))
                    begin
                      reg886 <= (reg880[(3'h5):(3'h4)] ^~ (reg881 << $unsigned($signed(wire870))));
                      reg887 <= (8'ha7);
                      reg888 <= reg886;
                    end
                end
              else
                begin
                  reg884 <= ($signed($signed((|(8'hb9)))) & ($signed((reg878 >>> wire871)) <= wire873[(4'h9):(4'h8)]));
                  for (forvar885 = (1'h0); (forvar885 < (2'h3)); forvar885 = (forvar885 + (1'h1)))
                    begin
                      reg886 <= (-$signed(reg881[(3'h5):(2'h3)]));
                      reg887 <= (&{{$signed(reg886)}});
                      reg888 <= ({((^reg880) >= (wire872 ~^ forvar885))} ?
                          (($signed(reg879) | wire872[(3'h4):(2'h2)]) ?
                              forvar881 : {$unsigned(reg879)}) : {wire870[(2'h3):(2'h2)]});
                    end
                  reg889 <= ($unsigned(forvar885) || $unsigned({(wire871 ?
                          wire870 : reg883)}));
                end
              for (forvar890 = (1'h0); (forvar890 < (2'h3)); forvar890 = (forvar890 + (1'h1)))
                begin
                  if (reg876)
                    begin
                      reg891 <= $unsigned($unsigned($unsigned((reg889 ?
                          (8'h9d) : wire869))));
                      reg892 <= reg888[(3'h5):(1'h1)];
                      reg893 <= reg892[(4'h9):(3'h6)];
                    end
                  else
                    begin
                      reg891 <= (reg881[(2'h2):(1'h1)] + {$unsigned($signed(reg877))});
                      reg892 <= ((reg883[(2'h2):(1'h1)] ?
                              (~reg889) : $signed($unsigned(forvar874))) ?
                          ($unsigned($unsigned((8'ha9))) ~^ wire871[(3'h6):(1'h1)]) : (($signed((8'hb1)) ?
                                  forvar879[(4'h8):(1'h1)] : reg893) ?
                              wire868 : $signed(((8'ha5) - forvar885))));
                      reg893 <= ($unsigned($signed(((8'ha8) >>> reg883))) - $signed(forvar881[(3'h4):(2'h2)]));
                      reg894 <= (8'ha2);
                    end
                  for (forvar895 = (1'h0); (forvar895 < (2'h3)); forvar895 = (forvar895 + (1'h1)))
                    begin
                      reg896 <= ($signed((wire872 * (reg887 ?
                              forvar895 : reg880))) ?
                          forvar890[(3'h5):(3'h4)] : $signed(reg891[(2'h2):(1'h1)]));
                      reg897 <= (forvar890 << $unsigned(reg886[(2'h2):(2'h2)]));
                    end
                  reg898 <= $unsigned((8'hba));
                  if ({$unsigned(wire871)})
                    begin
                      reg899 <= reg887;
                      reg900 <= $unsigned($unsigned((reg898 ?
                          (reg877 ? reg879 : wire870) : $unsigned((8'hb3)))));
                    end
                  else
                    begin
                      reg899 <= ((wire870[(1'h1):(1'h1)] >>> $signed((forvar881 ^~ (8'h9c)))) | {$unsigned($signed(reg889))});
                    end
                end
            end
          else
            begin
              if ($signed(($unsigned($signed(reg899)) ^ $signed((^~reg889)))))
                begin
                  reg877 <= (((~&reg879) ?
                      (-reg881) : (reg894[(2'h2):(2'h2)] ?
                          (~|reg878) : reg896)) == ($unsigned($signed(reg891)) ?
                      (8'ha4) : ((reg900 > forvar874) ?
                          $unsigned((8'ha3)) : (~&reg884))));
                end
              else
                begin
                  if (reg876[(1'h0):(1'h0)])
                    begin
                      reg877 <= (~|$unsigned($unsigned(reg898)));
                      reg878 <= {reg881};
                      reg879 <= reg887;
                    end
                  else
                    begin
                      reg877 <= $signed(reg894[(2'h2):(2'h2)]);
                    end
                  for (forvar880 = (1'h0); (forvar880 < (1'h0)); forvar880 = (forvar880 + (1'h1)))
                    begin
                      reg881 <= wire868;
                      reg882 <= ($signed((reg876[(3'h7):(3'h5)] && wire868[(4'ha):(4'ha)])) <= reg894);
                    end
                  if (((forvar875[(4'hb):(2'h2)] ?
                      $unsigned({forvar881}) : ($signed(reg896) ?
                          wire868 : $signed(reg879))) & (~((reg881 ?
                          wire868 : wire871) ?
                      forvar895 : forvar875))))
                    begin
                      reg883 <= ({{(forvar895 | (8'ha9))}} ?
                          $unsigned((^reg896[(3'h6):(3'h4)])) : (~$signed((forvar880 ?
                              (8'ha1) : (8'hb6)))));
                      reg884 <= {forvar881[(2'h3):(1'h1)]};
                    end
                  else
                    begin
                      reg883 <= $unsigned(wire869);
                      reg884 <= {forvar885};
                      reg885 <= ($signed(((+reg883) > (8'hb1))) && (|((reg878 ?
                              reg899 : forvar881) ?
                          (reg886 ?
                              wire870 : reg882) : reg880[(4'hc):(4'hb)])));
                    end
                end
            end
          for (forvar901 = (1'h0); (forvar901 < (1'h1)); forvar901 = (forvar901 + (1'h1)))
            begin
              reg902 <= ($signed($unsigned(reg893)) - (8'ha5));
              if ({(~^({(8'hb6)} ? reg902 : forvar880))})
                begin
                  if ($signed((reg898[(3'h7):(2'h3)] ?
                      ((reg886 ~^ reg877) >> (!forvar901)) : (-(forvar875 ?
                          reg893 : reg888)))))
                    begin
                      reg903 <= forvar885[(1'h1):(1'h1)];
                      reg904 <= (!{reg885});
                    end
                  else
                    begin
                      reg903 <= (reg904 ?
                          forvar895[(2'h2):(1'h0)] : $unsigned($signed($unsigned((8'hac)))));
                      reg904 <= ((|$unsigned(reg903)) ?
                          ((reg900[(3'h6):(3'h6)] >> $signed(reg877)) ?
                              (|(reg876 + forvar874)) : reg876) : (({reg904} >> ((8'ha3) ?
                                  wire870 : forvar881)) ?
                              forvar874[(2'h2):(1'h0)] : {{wire869}}));
                    end
                  for (forvar905 = (1'h0); (forvar905 < (1'h1)); forvar905 = (forvar905 + (1'h1)))
                    begin
                      reg906 <= ((forvar875[(2'h3):(2'h3)] & reg904[(4'ha):(3'h5)]) ?
                          {$signed(reg879[(3'h4):(3'h4)])} : (forvar885 ?
                              (^~((8'hb1) ~^ forvar880)) : $unsigned($signed(reg886))));
                    end
                end
              else
                begin
                  if ((&(~^$unsigned(reg888))))
                    begin
                      reg903 <= reg902[(2'h2):(2'h2)];
                      reg904 <= ((reg888 ?
                          {(reg878 >>> reg894)} : {$unsigned(reg885)}) == ({((8'ha2) ?
                              reg882 : (8'h9d))} || wire870));
                      reg905 <= $unsigned($signed((reg884 ~^ (reg876 ?
                          reg878 : wire869))));
                    end
                  else
                    begin
                      reg903 <= {$signed($signed($signed(forvar880)))};
                      reg904 <= reg898;
                    end
                  for (forvar906 = (1'h0); (forvar906 < (1'h1)); forvar906 = (forvar906 + (1'h1)))
                    begin
                      reg907 <= ($unsigned(($signed(reg903) <= $unsigned(forvar879))) & (((~|forvar885) ?
                              reg892[(2'h3):(2'h2)] : {(8'ha2)}) ?
                          $signed($signed(reg876)) : (~|(^forvar890))));
                      reg908 <= ($unsigned(reg887[(1'h0):(1'h0)]) ?
                          $signed(reg889[(3'h4):(2'h2)]) : (reg879 ?
                              reg898[(3'h4):(1'h0)] : ((reg898 ?
                                      reg894 : reg884) ?
                                  $signed(reg881) : $signed(reg898))));
                      reg909 <= ((~^$signed($signed((8'hac)))) ?
                          reg883[(2'h3):(2'h2)] : ((~(^reg906)) > $unsigned((^reg900))));
                      reg910 <= $unsigned((~&(reg909[(2'h3):(2'h2)] * $signed(wire872))));
                    end
                  if ((((^~(^forvar895)) ^~ $signed(reg876)) ?
                      reg877 : reg886[(1'h1):(1'h0)]))
                    begin
                      reg911 <= $signed(forvar901);
                    end
                  else
                    begin
                      reg911 <= (~$signed($unsigned($signed(reg887))));
                      reg912 <= $unsigned((~($signed(reg886) * forvar879[(3'h7):(3'h7)])));
                    end
                  for (forvar913 = (1'h0); (forvar913 < (1'h0)); forvar913 = (forvar913 + (1'h1)))
                    begin
                      reg914 <= $unsigned((~^$signed({reg882})));
                      reg915 <= $signed(($unsigned((~|reg877)) ?
                          $signed((forvar890 < reg878)) : (~|(reg886 ?
                              reg914 : reg876))));
                      reg916 <= wire870[(2'h3):(1'h1)];
                      reg917 <= reg910[(2'h3):(1'h1)];
                    end
                end
            end
          if ((forvar880 ?
              (8'ha3) : $signed($signed((reg894 ? forvar906 : reg916)))))
            begin
              for (forvar918 = (1'h0); (forvar918 < (1'h1)); forvar918 = (forvar918 + (1'h1)))
                begin
                  if ($unsigned({(&(reg896 - (8'h9f)))}))
                    begin
                      reg919 <= forvar901[(4'hc):(4'ha)];
                    end
                  else
                    begin
                      reg919 <= reg897[(3'h4):(3'h4)];
                      reg920 <= reg896[(2'h3):(2'h2)];
                      reg921 <= (reg885[(4'h8):(3'h6)] >>> (((^forvar875) ?
                              $signed(reg917) : (forvar875 ?
                                  forvar918 : forvar881)) ?
                          {(~|wire871)} : ((forvar879 ^ reg887) ?
                              (reg882 != forvar875) : {reg879})));
                    end
                  for (forvar922 = (1'h0); (forvar922 < (2'h3)); forvar922 = (forvar922 + (1'h1)))
                    begin
                      reg923 <= ((8'ha6) ?
                          $signed(reg886[(3'h4):(1'h0)]) : $unsigned({(reg893 > reg907)}));
                    end
                  if (({reg911} ? reg911 : forvar879[(3'h5):(3'h4)]))
                    begin
                      reg924 <= ((reg905[(2'h3):(1'h1)] - ($signed(reg909) ?
                          (8'haa) : $signed(reg892))) >>> $signed((forvar906[(4'h8):(2'h3)] ?
                          $signed(forvar895) : ((8'hb6) ? reg914 : reg921))));
                      reg925 <= {$unsigned($unsigned($unsigned(reg908)))};
                      reg926 <= (+((!(forvar922 & reg898)) ?
                          {(reg911 ? wire872 : reg917)} : ($signed(reg924) ?
                              (~reg879) : (forvar918 ~^ reg900))));
                    end
                  else
                    begin
                      reg924 <= ($unsigned($signed($unsigned(reg881))) >>> reg920[(2'h2):(2'h2)]);
                      reg925 <= reg920[(1'h1):(1'h1)];
                      reg926 <= reg907;
                    end
                  reg927 <= reg891;
                end
            end
          else
            begin
              for (forvar918 = (1'h0); (forvar918 < (2'h3)); forvar918 = (forvar918 + (1'h1)))
                begin
                  reg919 <= wire872[(4'ha):(3'h7)];
                  for (forvar920 = (1'h0); (forvar920 < (1'h1)); forvar920 = (forvar920 + (1'h1)))
                    begin
                      reg921 <= (((|(~^wire870)) ?
                              ((wire870 ? forvar913 : reg879) ?
                                  $unsigned(forvar879) : reg886[(1'h1):(1'h1)]) : (^~$signed((8'haf)))) ?
                          $signed((~|(!reg889))) : ({(reg907 >= reg903)} ?
                              {(reg886 ? reg876 : reg884)} : (reg909 ?
                                  (forvar906 << reg888) : (reg887 ?
                                      reg881 : reg882))));
                      reg922 <= reg920[(2'h2):(1'h1)];
                      reg923 <= reg914;
                    end
                end
              for (forvar924 = (1'h0); (forvar924 < (1'h0)); forvar924 = (forvar924 + (1'h1)))
                begin
                  reg925 <= $signed(((~^$signed(reg903)) ?
                      (8'hb4) : $signed(reg879)));
                end
              if (((($signed(reg889) | (&reg917)) ?
                  ((wire871 ?
                      reg888 : reg893) == $unsigned((8'ha8))) : $unsigned(reg892)) < $unsigned(({forvar885} ?
                  (~reg914) : $signed(forvar922)))))
                begin
                  reg926 <= (reg906 <<< {reg926[(4'hd):(3'h6)]});
                  reg927 <= (reg915[(2'h2):(1'h1)] < $unsigned(($signed(reg920) ?
                      $signed(reg923) : reg883[(1'h1):(1'h1)])));
                  if ($signed(reg897[(1'h1):(1'h0)]))
                    begin
                      reg928 <= (((reg903 ?
                              (reg909 ? reg881 : reg923) : (~&forvar875)) ?
                          $signed(((8'ha7) <= reg879)) : (&forvar890[(3'h7):(2'h3)])) <<< wire873);
                    end
                  else
                    begin
                      reg928 <= $signed((reg907 && forvar920[(3'h7):(2'h3)]));
                    end
                  for (forvar929 = (1'h0); (forvar929 < (2'h3)); forvar929 = (forvar929 + (1'h1)))
                    begin
                      reg930 <= {(reg926 ~^ {reg896})};
                      reg931 <= reg879;
                      reg932 <= $signed({((~^(8'hb2)) ~^ (reg902 ?
                              reg880 : reg886))});
                    end
                end
              else
                begin
                  if ($unsigned($unsigned(((!(8'ha7)) ?
                      (|reg896) : $signed(reg915)))))
                    begin
                      reg926 <= {($signed((^reg906)) ?
                              $signed($unsigned(reg879)) : {reg897[(4'hd):(4'hd)]})};
                      reg927 <= $unsigned(forvar920);
                    end
                  else
                    begin
                      reg926 <= (reg930 ^~ (8'hb8));
                      reg927 <= wire871;
                      reg928 <= (((&(reg917 ^ reg932)) ?
                          {{reg879}} : (reg910[(3'h7):(2'h2)] ?
                              reg903 : reg907[(3'h4):(1'h1)])) * reg885);
                    end
                  if ($signed(forvar881))
                    begin
                      reg929 <= (~^$unsigned(wire872[(2'h3):(1'h1)]));
                    end
                  else
                    begin
                      reg929 <= (&($signed($unsigned(reg897)) ?
                          $signed($signed((8'hb0))) : $signed(reg902[(2'h2):(1'h0)])));
                      reg930 <= $unsigned((reg932[(3'h4):(1'h1)] ?
                          $unsigned(((8'hb3) || reg882)) : ((wire870 ?
                              reg917 : (8'hb9)) >= (~(8'ha2)))));
                      reg931 <= $signed($signed({(-reg878)}));
                      reg932 <= (-$unsigned($unsigned($unsigned(reg927))));
                    end
                  if ($signed(reg896[(2'h2):(1'h1)]))
                    begin
                      reg933 <= $unsigned((({reg923} < (~&reg888)) <<< {$unsigned(reg896)}));
                      reg934 <= reg883;
                      reg935 <= (8'ha8);
                    end
                  else
                    begin
                      reg933 <= $unsigned($signed(reg888));
                      reg934 <= $signed((-({reg916} ? (~|reg921) : reg922)));
                      reg935 <= reg931;
                    end
                  if ({($unsigned(reg903[(2'h2):(1'h0)]) ?
                          {reg920[(2'h3):(1'h1)]} : ({(8'h9f)} ^~ {reg907}))})
                    begin
                      reg936 <= $unsigned(((+$signed(wire869)) ?
                          ((reg924 ? reg910 : reg881) ?
                              {reg893} : (reg914 ?
                                  forvar880 : reg907)) : $signed(((8'ha4) ?
                              reg925 : reg912))));
                      reg937 <= {forvar875[(1'h1):(1'h1)]};
                      reg938 <= {{reg907}};
                      reg939 <= (+(($signed(wire870) > forvar906) ?
                          {{reg912}} : $unsigned((~&reg891))));
                    end
                  else
                    begin
                      reg936 <= (~reg908);
                      reg937 <= forvar922[(4'ha):(3'h4)];
                    end
                end
              if (reg898)
                begin
                  if (((($unsigned(reg884) ? (reg933 != reg896) : reg892) ?
                          ((forvar895 == forvar913) & ((8'haa) ?
                              reg896 : reg879)) : reg931) ?
                      reg904 : $unsigned(({reg892} ?
                          reg915[(2'h2):(1'h1)] : ((8'h9c) ^ reg892)))))
                    begin
                      reg940 <= $unsigned((~|$signed((reg915 ?
                          reg914 : reg930))));
                      reg941 <= (((reg907 ?
                              reg905[(1'h1):(1'h1)] : ((8'hab) << reg931)) ?
                          reg908[(2'h3):(2'h3)] : forvar895[(1'h1):(1'h1)]) ~^ ($signed((8'hac)) >= {$signed(wire871)}));
                    end
                  else
                    begin
                      reg940 <= ((~^(~|(8'hae))) - forvar895);
                      reg941 <= reg923;
                      reg942 <= forvar874[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  if ($unsigned({reg878}))
                    begin
                      reg940 <= (~|$signed(((forvar885 && reg939) ?
                          (reg878 ^~ wire868) : wire873)));
                      reg941 <= {forvar905};
                    end
                  else
                    begin
                      reg940 <= ($unsigned(($signed(reg937) ?
                              $unsigned(forvar920) : (forvar901 <<< reg938))) ?
                          {(~|((8'ha8) <= reg919))} : (-($signed((8'hb4)) ?
                              reg936[(3'h5):(2'h3)] : $unsigned((8'ha5)))));
                      reg941 <= $unsigned($unsigned(((-reg914) <= (^reg893))));
                    end
                  for (forvar942 = (1'h0); (forvar942 < (2'h3)); forvar942 = (forvar942 + (1'h1)))
                    begin
                      reg943 <= ((!forvar885[(2'h3):(2'h2)]) ?
                          $unsigned(reg927[(3'h7):(3'h4)]) : forvar924);
                      reg944 <= reg878;
                      reg945 <= {$signed(reg894)};
                      reg946 <= (~^reg936[(1'h1):(1'h0)]);
                    end
                  reg947 <= (reg916 ?
                      (reg936 >>> ((8'hb7) ?
                          (^reg886) : reg897)) : forvar942[(4'ha):(3'h4)]);
                  for (forvar948 = (1'h0); (forvar948 < (1'h0)); forvar948 = (forvar948 + (1'h1)))
                    begin
                      reg949 <= (forvar924[(1'h1):(1'h0)] != reg877[(3'h6):(3'h5)]);
                    end
                end
            end
        end
    end
  assign wire950 = (reg911[(2'h2):(1'h1)] ?
                       $unsigned((|$unsigned(reg904))) : reg910);
  assign wire951 = wire871[(4'he):(3'h5)];
  always
    @(posedge clk) begin
      for (forvar952 = (1'h0); (forvar952 < (1'h0)); forvar952 = (forvar952 + (1'h1)))
        begin
          reg953 <= reg931[(2'h2):(2'h2)];
          if (($signed($signed((reg938 <<< reg930))) ?
              (reg876 ?
                  ($signed(forvar952) ^~ $signed(reg923)) : $unsigned(reg893)) : $signed(reg914[(3'h6):(2'h2)])))
            begin
              reg954 <= $signed({{$signed(reg885)}});
              if ($unsigned(reg954))
                begin
                  reg955 <= wire873;
                  reg956 <= (~&wire872[(3'h7):(3'h7)]);
                  for (forvar957 = (1'h0); (forvar957 < (1'h0)); forvar957 = (forvar957 + (1'h1)))
                    begin
                      reg958 <= wire870;
                    end
                  for (forvar959 = (1'h0); (forvar959 < (1'h1)); forvar959 = (forvar959 + (1'h1)))
                    begin
                      reg960 <= $unsigned($unsigned($unsigned((wire870 ?
                          reg922 : reg922))));
                      reg961 <= $unsigned(reg907[(1'h0):(1'h0)]);
                      reg962 <= reg956;
                      reg963 <= reg888;
                    end
                end
              else
                begin
                  if ($signed(reg879[(4'h9):(2'h2)]))
                    begin
                      reg955 <= (^~(($signed(wire872) ?
                          reg917 : reg906[(3'h5):(1'h1)]) >>> $signed((reg921 - reg878))));
                      reg956 <= {reg909[(3'h7):(2'h3)]};
                      reg957 <= reg919[(3'h4):(2'h2)];
                      reg958 <= reg879;
                    end
                  else
                    begin
                      reg955 <= $unsigned(reg915[(1'h1):(1'h0)]);
                    end
                  if (((((^reg925) ?
                          $unsigned(wire951) : reg928[(4'hb):(4'h8)]) && $signed($unsigned(reg923))) ?
                      (reg904 && reg902) : $signed(reg896)))
                    begin
                      reg959 <= (reg917[(2'h2):(2'h2)] ? reg925 : reg919);
                      reg960 <= $signed(reg925);
                      reg961 <= $signed((|reg938[(3'h4):(1'h0)]));
                      reg962 <= (~^reg955[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg959 <= (8'h9c);
                      reg960 <= reg946;
                    end
                end
              if (reg911[(1'h1):(1'h0)])
                begin
                  reg964 <= reg884[(1'h0):(1'h0)];
                  for (forvar965 = (1'h0); (forvar965 < (2'h2)); forvar965 = (forvar965 + (1'h1)))
                    begin
                      reg966 <= reg924[(4'hc):(3'h5)];
                      reg967 <= $signed(($unsigned($signed(reg941)) <<< $signed(reg963[(2'h2):(1'h1)])));
                    end
                  if ((8'ha0))
                    begin
                      reg968 <= reg928[(4'hc):(4'ha)];
                      reg969 <= wire868[(1'h0):(1'h0)];
                      reg970 <= (^reg893[(3'h7):(3'h4)]);
                    end
                  else
                    begin
                      reg968 <= ((8'h9e) ?
                          $unsigned(((&reg889) ?
                              ((8'haa) >>> reg894) : {forvar959})) : $signed($unsigned(reg893[(4'h8):(1'h1)])));
                      reg969 <= $signed($unsigned({reg898}));
                      reg970 <= wire871;
                    end
                end
              else
                begin
                  reg964 <= $signed((~|((8'hb7) ?
                      reg924[(4'h9):(3'h6)] : $unsigned(wire870))));
                  if ($signed((~((reg942 <= reg889) ?
                      {reg909} : $unsigned(reg933)))))
                    begin
                      reg965 <= ($unsigned($unsigned({reg888})) ?
                          $unsigned((!$signed(reg960))) : ((reg892 ?
                              $signed(reg924) : (reg967 >> reg887)) && (~^(^(8'h9c)))));
                      reg966 <= ($unsigned((~|(reg925 ? reg882 : reg957))) ?
                          $signed($unsigned((reg931 ?
                              (8'hae) : reg893))) : $signed(($unsigned(reg877) * $signed(reg940))));
                      reg967 <= (^~$signed(reg961[(4'h8):(1'h1)]));
                      reg968 <= wire868[(4'hb):(3'h7)];
                    end
                  else
                    begin
                      reg965 <= reg916[(2'h2):(1'h0)];
                    end
                  reg969 <= (~(8'hb4));
                  reg970 <= {(^~((&reg943) ?
                          $signed(reg970) : $signed((8'haf))))};
                end
              for (forvar971 = (1'h0); (forvar971 < (1'h1)); forvar971 = (forvar971 + (1'h1)))
                begin
                  reg972 <= $signed((8'hae));
                  if ((~|((reg897[(4'h8):(2'h2)] >> ((8'hb9) ?
                      reg899 : reg942)) ~^ reg942[(1'h1):(1'h1)])))
                    begin
                      reg973 <= $signed($signed((~^reg909)));
                      reg974 <= reg946;
                    end
                  else
                    begin
                      reg973 <= reg904[(3'h4):(1'h0)];
                      reg974 <= $unsigned((reg912 ?
                          wire950[(3'h5):(1'h0)] : (~|{forvar965})));
                      reg975 <= $unsigned((((reg945 != reg880) - (~|reg919)) ?
                          $signed(forvar971) : wire950));
                    end
                  reg976 <= ($unsigned($signed((reg967 + forvar959))) ?
                      $unsigned($signed(reg959)) : reg965[(3'h4):(3'h4)]);
                end
            end
          else
            begin
              reg954 <= (+{reg905[(2'h2):(1'h1)]});
            end
        end
    end
  assign wire977 = reg877[(2'h3):(2'h2)];
  assign wire978 = (8'hac);
  assign wire979 = reg934[(3'h6):(2'h3)];
  module980 #() modinst1970 (.wire985(reg963), .wire984(reg888), .wire981(reg943), .wire983(reg964), .wire982(reg907), .clk(clk), .y(wire1969));
  assign wire1971 = (-(&(^~(reg883 ? wire870 : reg946))));
  assign wire1972 = {$signed((^(-(8'hae))))};
  always
    @(posedge clk) begin
      for (forvar1973 = (1'h0); (forvar1973 < (2'h3)); forvar1973 = (forvar1973 + (1'h1)))
        begin
          for (forvar1974 = (1'h0); (forvar1974 < (1'h1)); forvar1974 = (forvar1974 + (1'h1)))
            begin
              for (forvar1975 = (1'h0); (forvar1975 < (1'h0)); forvar1975 = (forvar1975 + (1'h1)))
                begin
                  for (forvar1976 = (1'h0); (forvar1976 < (1'h0)); forvar1976 = (forvar1976 + (1'h1)))
                    begin
                      reg1977 <= ({$signed((8'h9e))} <= forvar1974);
                      reg1978 <= ((((reg958 << reg882) ?
                              (reg962 ?
                                  reg927 : wire1971) : (reg956 + reg949)) >= ({reg893} >> wire872)) ?
                          $signed(($signed(reg965) ?
                              $unsigned(reg958) : (reg967 <= reg943))) : reg893[(4'h8):(3'h6)]);
                    end
                  for (forvar1979 = (1'h0); (forvar1979 < (1'h1)); forvar1979 = (forvar1979 + (1'h1)))
                    begin
                      reg1980 <= ({$signed((wire871 ?
                              reg937 : reg943))} ^~ reg974);
                      reg1981 <= (reg942[(2'h2):(1'h0)] ?
                          (((reg920 == (8'ha5)) ?
                              ((8'h9d) - wire868) : $unsigned((8'hb1))) - $signed((reg900 >> reg940))) : {(&$unsigned((8'haa)))});
                      reg1982 <= reg898;
                      reg1983 <= $signed(($signed(reg884) ?
                          $unsigned((reg962 == reg949)) : reg907));
                    end
                end
              reg1984 <= ($unsigned(({reg1980} ?
                      {reg878} : reg945[(4'h9):(1'h0)])) ?
                  $unsigned(((^~reg974) && ((8'haa) ^~ reg881))) : (!$unsigned((^reg881))));
            end
          for (forvar1985 = (1'h0); (forvar1985 < (1'h1)); forvar1985 = (forvar1985 + (1'h1)))
            begin
              for (forvar1986 = (1'h0); (forvar1986 < (1'h1)); forvar1986 = (forvar1986 + (1'h1)))
                begin
                  reg1987 <= $signed($unsigned(reg903[(2'h2):(1'h0)]));
                  for (forvar1988 = (1'h0); (forvar1988 < (1'h1)); forvar1988 = (forvar1988 + (1'h1)))
                    begin
                      reg1989 <= $unsigned({(+(reg959 ? reg959 : reg899))});
                      reg1990 <= $signed((reg936 & {(reg945 <= reg970)}));
                    end
                  reg1991 <= (~&$unsigned($signed((^reg876))));
                  for (forvar1992 = (1'h0); (forvar1992 < (1'h1)); forvar1992 = (forvar1992 + (1'h1)))
                    begin
                      reg1993 <= (reg902[(4'hb):(2'h2)] <= wire872);
                      reg1994 <= reg966;
                    end
                end
              if ($unsigned(reg898[(2'h3):(1'h0)]))
                begin
                  for (forvar1995 = (1'h0); (forvar1995 < (2'h2)); forvar1995 = (forvar1995 + (1'h1)))
                    begin
                      reg1996 <= {{(reg939 ?
                                  reg929[(1'h1):(1'h0)] : reg906[(3'h5):(2'h2)])}};
                      reg1997 <= {(8'h9f)};
                      reg1998 <= reg955;
                    end
                  if (reg925[(3'h7):(3'h6)])
                    begin
                      reg1999 <= reg953;
                      reg2000 <= $signed((&({reg881} ~^ $signed(reg954))));
                      reg2001 <= (reg882 <<< (({reg912} ?
                          $signed(reg884) : (-reg945)) >= (reg954[(1'h0):(1'h0)] < (reg1994 >> (8'ha3)))));
                    end
                  else
                    begin
                      reg1999 <= $unsigned(reg938);
                    end
                  if (($unsigned($unsigned(reg940)) && reg920[(2'h2):(2'h2)]))
                    begin
                      reg2002 <= reg934;
                      reg2003 <= ((&$unsigned({reg921})) ? reg956 : forvar1975);
                      reg2004 <= (reg946 ?
                          $unsigned({$unsigned((8'hb3))}) : reg936[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg2002 <= reg942;
                    end
                  for (forvar2005 = (1'h0); (forvar2005 < (2'h3)); forvar2005 = (forvar2005 + (1'h1)))
                    begin
                      reg2006 <= reg885;
                    end
                end
              else
                begin
                  for (forvar1995 = (1'h0); (forvar1995 < (2'h2)); forvar1995 = (forvar1995 + (1'h1)))
                    begin
                      reg1996 <= ((&(^~(reg939 >>> reg883))) ?
                          forvar2005[(3'h4):(2'h2)] : reg909);
                      reg1997 <= reg1990[(1'h0):(1'h0)];
                    end
                  for (forvar1998 = (1'h0); (forvar1998 < (2'h2)); forvar1998 = (forvar1998 + (1'h1)))
                    begin
                      reg1999 <= forvar1986;
                      reg2000 <= reg923;
                      reg2001 <= reg973;
                    end
                  reg2002 <= reg965;
                end
              if (((8'hb6) + ((~^(reg921 ^~ wire1972)) ?
                  (~&(reg969 ^~ reg897)) : ($unsigned(reg931) | ((8'ha8) ?
                      reg947 : reg899)))))
                begin
                  reg2007 <= reg955[(2'h2):(1'h1)];
                  for (forvar2008 = (1'h0); (forvar2008 < (1'h0)); forvar2008 = (forvar2008 + (1'h1)))
                    begin
                      reg2009 <= ($unsigned(reg953) ?
                          (&(^~(|reg970))) : $unsigned($signed((reg903 ?
                              reg917 : reg936))));
                    end
                  for (forvar2010 = (1'h0); (forvar2010 < (2'h3)); forvar2010 = (forvar2010 + (1'h1)))
                    begin
                      reg2011 <= (($signed((reg907 ? (8'h9d) : wire1972)) ?
                          $signed($unsigned(reg877)) : reg942) - reg904[(3'h7):(3'h5)]);
                      reg2012 <= reg946;
                      reg2013 <= forvar2008[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  reg2007 <= $unsigned($unsigned($signed((reg1991 << reg958))));
                  for (forvar2008 = (1'h0); (forvar2008 < (1'h0)); forvar2008 = (forvar2008 + (1'h1)))
                    begin
                      reg2009 <= $signed((((reg1980 ?
                              reg953 : forvar1998) < (wire869 ^~ reg908)) ?
                          $unsigned((~wire978)) : reg2002[(4'ha):(4'ha)]));
                      reg2010 <= (forvar1986 ?
                          (((forvar1974 << reg887) ?
                              (^~reg946) : (reg949 ?
                                  reg926 : reg1977)) <<< ((reg972 ?
                              (8'h9f) : reg938) <<< reg933)) : (^(^~(8'hab))));
                      reg2011 <= reg935;
                      reg2012 <= forvar1974;
                    end
                end
            end
        end
      for (forvar2014 = (1'h0); (forvar2014 < (2'h2)); forvar2014 = (forvar2014 + (1'h1)))
        begin
          for (forvar2015 = (1'h0); (forvar2015 < (2'h3)); forvar2015 = (forvar2015 + (1'h1)))
            begin
              if ((~&($signed($signed(reg902)) ?
                  reg1989 : $unsigned($signed(reg946)))))
                begin
                  for (forvar2016 = (1'h0); (forvar2016 < (2'h3)); forvar2016 = (forvar2016 + (1'h1)))
                    begin
                      reg2017 <= $signed(((wire1971[(2'h2):(2'h2)] >> forvar2008) ?
                          (reg927[(1'h0):(1'h0)] >> $signed(forvar1992)) : reg927[(1'h1):(1'h0)]));
                      reg2018 <= $unsigned($unsigned($unsigned({forvar2008})));
                      reg2019 <= ((8'haa) || {((|(8'ha3)) + (reg892 ?
                              reg910 : reg891))});
                    end
                  for (forvar2020 = (1'h0); (forvar2020 < (2'h3)); forvar2020 = (forvar2020 + (1'h1)))
                    begin
                      reg2021 <= (+$signed({(reg1993 ? reg915 : reg1991)}));
                      reg2022 <= ($signed(reg924) - (($signed(reg885) ?
                          (reg966 ?
                              reg889 : reg917) : $unsigned(wire871)) != $signed((reg974 ?
                          (8'hb6) : reg887))));
                      reg2023 <= ((~|$unsigned((reg2002 < reg926))) ?
                          ((reg1993[(4'h9):(3'h7)] || $signed(reg884)) >>> $unsigned((reg891 ?
                              forvar1975 : reg879))) : ($signed($unsigned((8'hb7))) == $unsigned(reg936)));
                    end
                  for (forvar2024 = (1'h0); (forvar2024 < (1'h0)); forvar2024 = (forvar2024 + (1'h1)))
                    begin
                      reg2025 <= $unsigned((|reg959[(4'he):(4'he)]));
                    end
                  for (forvar2026 = (1'h0); (forvar2026 < (1'h1)); forvar2026 = (forvar2026 + (1'h1)))
                    begin
                      reg2027 <= reg1999[(4'hc):(4'ha)];
                      reg2028 <= (reg954 <<< $signed($signed((!(8'hb5)))));
                      reg2029 <= (8'hb9);
                    end
                end
              else
                begin
                  if (($unsigned({(~&forvar2008)}) * $signed(({(8'hac)} | $signed(reg976)))))
                    begin
                      reg2016 <= reg2021;
                      reg2017 <= $signed(reg962[(4'he):(3'h4)]);
                      reg2018 <= ((reg946 - {$unsigned(wire1971)}) ?
                          $unsigned(forvar2008) : ((8'ha1) ?
                              ($unsigned(reg894) ?
                                  {reg969} : (+wire1971)) : $signed(forvar2008)));
                      reg2019 <= $signed((&($unsigned(reg946) != (reg955 ?
                          reg905 : reg879))));
                    end
                  else
                    begin
                      reg2016 <= reg1989[(3'h5):(2'h2)];
                    end
                  for (forvar2020 = (1'h0); (forvar2020 < (1'h1)); forvar2020 = (forvar2020 + (1'h1)))
                    begin
                      reg2021 <= reg897[(2'h3):(2'h3)];
                    end
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module980  (y, clk, wire981, wire982, wire983, wire984, wire985);
  output wire [(32'h14ac):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire981;
  input wire [(4'hb):(1'h0)] wire982;
  input wire signed [(4'h9):(1'h0)] wire983;
  input wire [(2'h3):(1'h0)] wire984;
  input wire signed [(3'h4):(1'h0)] wire985;
  wire [(4'ha):(1'h0)] wire1968;
  wire [(3'h6):(1'h0)] wire1967;
  wire signed [(5'h10):(1'h0)] wire1908;
  wire signed [(4'hb):(1'h0)] wire1907;
  wire signed [(3'h6):(1'h0)] wire1861;
  wire signed [(4'hc):(1'h0)] wire1705;
  wire [(3'h4):(1'h0)] wire986;
  wire signed [(4'h8):(1'h0)] wire987;
  wire signed [(4'hd):(1'h0)] wire1146;
  wire [(4'hf):(1'h0)] wire1147;
  wire signed [(4'hc):(1'h0)] wire1658;
  reg [(4'hd):(1'h0)] reg1950 = (1'h0);
  reg [(4'hc):(1'h0)] reg1966 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1965 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1964 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1963 = (1'h0);
  reg [(4'hd):(1'h0)] reg1962 = (1'h0);
  reg [(5'h10):(1'h0)] reg1960 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1959 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1958 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1957 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1955 = (1'h0);
  reg [(4'he):(1'h0)] reg1954 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1946 = (1'h0);
  reg [(4'h9):(1'h0)] reg1953 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1952 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1951 = (1'h0);
  reg [(3'h4):(1'h0)] reg1949 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1948 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1947 = (1'h0);
  reg [(4'hf):(1'h0)] reg1945 = (1'h0);
  reg [(4'hd):(1'h0)] reg1944 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1943 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1941 = (1'h0);
  reg [(3'h5):(1'h0)] reg1940 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1939 = (1'h0);
  reg [(4'h9):(1'h0)] reg1937 = (1'h0);
  reg [(4'he):(1'h0)] reg1936 = (1'h0);
  reg [(4'hd):(1'h0)] reg1935 = (1'h0);
  reg [(4'h9):(1'h0)] reg1933 = (1'h0);
  reg [(4'h9):(1'h0)] reg1932 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1931 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1930 = (1'h0);
  reg [(4'hc):(1'h0)] reg1927 = (1'h0);
  reg [(5'h10):(1'h0)] reg1915 = (1'h0);
  reg [(5'h10):(1'h0)] reg1926 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1925 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1923 = (1'h0);
  reg [(2'h3):(1'h0)] reg1922 = (1'h0);
  reg [(4'hd):(1'h0)] reg1918 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1921 = (1'h0);
  reg [(2'h2):(1'h0)] reg1920 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1919 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1917 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1916 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1914 = (1'h0);
  reg [(4'hc):(1'h0)] reg1911 = (1'h0);
  reg [(4'he):(1'h0)] reg1910 = (1'h0);
  reg [(4'hc):(1'h0)] reg1906 = (1'h0);
  reg [(4'hb):(1'h0)] reg1905 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1904 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1903 = (1'h0);
  reg [(4'hb):(1'h0)] reg1902 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1901 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1900 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1899 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1898 = (1'h0);
  reg [(5'h10):(1'h0)] reg1897 = (1'h0);
  reg [(4'hf):(1'h0)] reg1896 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1895 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1894 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1888 = (1'h0);
  reg [(4'h9):(1'h0)] reg1887 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1883 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1871 = (1'h0);
  reg [(2'h3):(1'h0)] reg1893 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1892 = (1'h0);
  reg [(2'h2):(1'h0)] reg1891 = (1'h0);
  reg [(4'h9):(1'h0)] reg1890 = (1'h0);
  reg [(4'ha):(1'h0)] reg1889 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1886 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1885 = (1'h0);
  reg [(3'h5):(1'h0)] reg1878 = (1'h0);
  reg [(2'h3):(1'h0)] reg1882 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1881 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1880 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1879 = (1'h0);
  reg [(4'ha):(1'h0)] reg1877 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1876 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1875 = (1'h0);
  reg [(5'h10):(1'h0)] reg1874 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1873 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1872 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1870 = (1'h0);
  reg [(4'he):(1'h0)] reg1869 = (1'h0);
  reg [(2'h2):(1'h0)] reg1868 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1867 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1863 = (1'h0);
  reg [(3'h5):(1'h0)] reg1860 = (1'h0);
  reg [(2'h2):(1'h0)] reg1859 = (1'h0);
  reg [(3'h5):(1'h0)] reg1858 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1857 = (1'h0);
  reg [(4'ha):(1'h0)] reg1855 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1854 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1849 = (1'h0);
  reg [(4'he):(1'h0)] reg1851 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1850 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1848 = (1'h0);
  reg [(4'h8):(1'h0)] reg1847 = (1'h0);
  reg [(4'h9):(1'h0)] reg1846 = (1'h0);
  reg [(5'h10):(1'h0)] reg1845 = (1'h0);
  reg [(4'h8):(1'h0)] reg1844 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1843 = (1'h0);
  reg [(4'h9):(1'h0)] reg1842 = (1'h0);
  reg [(4'hb):(1'h0)] reg1839 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1838 = (1'h0);
  reg [(4'ha):(1'h0)] reg1836 = (1'h0);
  reg [(4'hc):(1'h0)] reg1835 = (1'h0);
  reg [(4'hc):(1'h0)] reg1834 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1833 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1832 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1831 = (1'h0);
  reg [(4'hd):(1'h0)] reg1830 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1829 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1828 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1824 = (1'h0);
  reg [(4'hd):(1'h0)] reg1823 = (1'h0);
  reg [(3'h4):(1'h0)] reg1822 = (1'h0);
  reg [(4'hb):(1'h0)] reg1821 = (1'h0);
  reg [(4'hd):(1'h0)] reg1819 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1818 = (1'h0);
  reg [(4'hf):(1'h0)] reg1817 = (1'h0);
  reg [(4'hf):(1'h0)] reg1816 = (1'h0);
  reg [(3'h7):(1'h0)] reg1814 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1813 = (1'h0);
  reg [(4'hd):(1'h0)] reg1812 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1809 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1808 = (1'h0);
  reg [(3'h6):(1'h0)] reg1807 = (1'h0);
  reg [(4'ha):(1'h0)] reg1806 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1803 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1801 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1800 = (1'h0);
  reg [(4'he):(1'h0)] reg1799 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1798 = (1'h0);
  reg [(4'hf):(1'h0)] reg1794 = (1'h0);
  reg [(3'h7):(1'h0)] reg1797 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1789 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1796 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1795 = (1'h0);
  reg [(4'h8):(1'h0)] reg1793 = (1'h0);
  reg [(4'hd):(1'h0)] reg1792 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1791 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1790 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1788 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1775 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1772 = (1'h0);
  reg [(3'h6):(1'h0)] reg1758 = (1'h0);
  reg [(3'h6):(1'h0)] reg1757 = (1'h0);
  reg [(4'hf):(1'h0)] reg1756 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1786 = (1'h0);
  reg [(5'h10):(1'h0)] reg1785 = (1'h0);
  reg [(5'h10):(1'h0)] reg1784 = (1'h0);
  reg [(2'h3):(1'h0)] reg1783 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1782 = (1'h0);
  reg [(2'h3):(1'h0)] reg1781 = (1'h0);
  reg [(5'h10):(1'h0)] reg1780 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1779 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1778 = (1'h0);
  reg [(4'hb):(1'h0)] reg1777 = (1'h0);
  reg [(3'h6):(1'h0)] reg1774 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1773 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1771 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1770 = (1'h0);
  reg [(2'h2):(1'h0)] reg1769 = (1'h0);
  reg [(2'h2):(1'h0)] reg1768 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1767 = (1'h0);
  reg [(4'hc):(1'h0)] reg1766 = (1'h0);
  reg [(2'h2):(1'h0)] reg1765 = (1'h0);
  reg [(3'h7):(1'h0)] reg1764 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1763 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1762 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1761 = (1'h0);
  reg [(3'h5):(1'h0)] reg1760 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1759 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1755 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1754 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1708 = (1'h0);
  reg [(4'hd):(1'h0)] reg1753 = (1'h0);
  reg [(4'h9):(1'h0)] reg1750 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1749 = (1'h0);
  reg [(2'h3):(1'h0)] reg1747 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1739 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1737 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1723 = (1'h0);
  reg [(4'hc):(1'h0)] reg1748 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1745 = (1'h0);
  reg [(2'h2):(1'h0)] reg1744 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1743 = (1'h0);
  reg [(3'h5):(1'h0)] reg1742 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1741 = (1'h0);
  reg [(4'he):(1'h0)] reg1740 = (1'h0);
  reg [(5'h10):(1'h0)] reg1731 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1726 = (1'h0);
  reg [(4'hf):(1'h0)] reg1738 = (1'h0);
  reg [(4'ha):(1'h0)] reg1736 = (1'h0);
  reg [(4'he):(1'h0)] reg1735 = (1'h0);
  reg [(3'h5):(1'h0)] reg1734 = (1'h0);
  reg [(4'hb):(1'h0)] reg1733 = (1'h0);
  reg [(4'ha):(1'h0)] reg1732 = (1'h0);
  reg [(4'ha):(1'h0)] reg1730 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1729 = (1'h0);
  reg [(4'h9):(1'h0)] reg1728 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1727 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1725 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1724 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1722 = (1'h0);
  reg [(2'h3):(1'h0)] reg1721 = (1'h0);
  reg [(3'h4):(1'h0)] reg1720 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1715 = (1'h0);
  reg [(4'hb):(1'h0)] reg1719 = (1'h0);
  reg [(4'hc):(1'h0)] reg1718 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1717 = (1'h0);
  reg [(4'hf):(1'h0)] reg1716 = (1'h0);
  reg [(3'h7):(1'h0)] reg1714 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1713 = (1'h0);
  reg [(4'h9):(1'h0)] reg1712 = (1'h0);
  reg [(3'h7):(1'h0)] reg1711 = (1'h0);
  reg [(2'h2):(1'h0)] reg1710 = (1'h0);
  reg [(4'hf):(1'h0)] reg1709 = (1'h0);
  reg [(5'h10):(1'h0)] reg1706 = (1'h0);
  reg [(5'h10):(1'h0)] reg1704 = (1'h0);
  reg [(4'hc):(1'h0)] reg1703 = (1'h0);
  reg [(4'hf):(1'h0)] reg1702 = (1'h0);
  reg [(4'ha):(1'h0)] reg1701 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1700 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1699 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1697 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1695 = (1'h0);
  reg [(4'hc):(1'h0)] reg1693 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1692 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1691 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1690 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1666 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1685 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1684 = (1'h0);
  reg [(3'h4):(1'h0)] reg1683 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1682 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1680 = (1'h0);
  reg [(3'h6):(1'h0)] reg1679 = (1'h0);
  reg [(3'h6):(1'h0)] reg1678 = (1'h0);
  reg [(4'h9):(1'h0)] reg1677 = (1'h0);
  reg [(4'he):(1'h0)] reg1676 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1675 = (1'h0);
  reg [(4'hb):(1'h0)] reg1673 = (1'h0);
  reg [(4'hb):(1'h0)] reg1671 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1670 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1669 = (1'h0);
  reg [(4'hb):(1'h0)] reg1668 = (1'h0);
  reg [(4'hb):(1'h0)] reg1665 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1664 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1663 = (1'h0);
  reg [(5'h10):(1'h0)] reg1662 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1660 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1097 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1090 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1145 = (1'h0);
  reg [(3'h7):(1'h0)] reg1144 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1143 = (1'h0);
  reg [(3'h4):(1'h0)] reg1142 = (1'h0);
  reg [(2'h2):(1'h0)] reg1141 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1139 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1138 = (1'h0);
  reg [(4'hf):(1'h0)] reg1137 = (1'h0);
  reg [(5'h10):(1'h0)] reg1135 = (1'h0);
  reg [(4'hd):(1'h0)] reg1134 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1133 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1131 = (1'h0);
  reg [(4'h9):(1'h0)] reg1127 = (1'h0);
  reg [(4'h8):(1'h0)] reg1132 = (1'h0);
  reg [(4'hd):(1'h0)] reg1130 = (1'h0);
  reg [(4'hb):(1'h0)] reg1129 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1128 = (1'h0);
  reg [(3'h4):(1'h0)] reg1126 = (1'h0);
  reg [(4'hd):(1'h0)] reg1125 = (1'h0);
  reg [(2'h2):(1'h0)] reg1124 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1123 = (1'h0);
  reg [(4'he):(1'h0)] reg1122 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1121 = (1'h0);
  reg [(4'h8):(1'h0)] reg1119 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1118 = (1'h0);
  reg [(3'h4):(1'h0)] reg1115 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1111 = (1'h0);
  reg [(3'h5):(1'h0)] reg1110 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1117 = (1'h0);
  reg [(3'h4):(1'h0)] reg1116 = (1'h0);
  reg [(3'h5):(1'h0)] reg1114 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1113 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1112 = (1'h0);
  reg [(2'h3):(1'h0)] reg1109 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1108 = (1'h0);
  reg [(2'h3):(1'h0)] reg1102 = (1'h0);
  reg [(4'h9):(1'h0)] reg1107 = (1'h0);
  reg [(2'h3):(1'h0)] reg1106 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1105 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1104 = (1'h0);
  reg [(3'h5):(1'h0)] reg1103 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1101 = (1'h0);
  reg [(3'h4):(1'h0)] reg1100 = (1'h0);
  reg [(4'hb):(1'h0)] reg1099 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1098 = (1'h0);
  reg [(3'h5):(1'h0)] reg1096 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1095 = (1'h0);
  reg [(4'hb):(1'h0)] reg1094 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1093 = (1'h0);
  reg [(5'h10):(1'h0)] reg1091 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1089 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1081 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1088 = (1'h0);
  reg [(4'ha):(1'h0)] reg1087 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1086 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1085 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1083 = (1'h0);
  reg [(3'h5):(1'h0)] reg1082 = (1'h0);
  reg [(4'ha):(1'h0)] reg1080 = (1'h0);
  reg [(3'h7):(1'h0)] reg1064 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1078 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1077 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1076 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1075 = (1'h0);
  reg [(2'h3):(1'h0)] reg1074 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1072 = (1'h0);
  reg [(4'hc):(1'h0)] reg1058 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1070 = (1'h0);
  reg [(4'h9):(1'h0)] reg1068 = (1'h0);
  reg [(4'hc):(1'h0)] reg1067 = (1'h0);
  reg [(2'h3):(1'h0)] reg1066 = (1'h0);
  reg [(4'h9):(1'h0)] reg1065 = (1'h0);
  reg [(4'ha):(1'h0)] reg1063 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1062 = (1'h0);
  reg [(4'hd):(1'h0)] reg1061 = (1'h0);
  reg [(4'ha):(1'h0)] reg1060 = (1'h0);
  reg [(2'h2):(1'h0)] reg1059 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1057 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1056 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1027 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1054 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1053 = (1'h0);
  reg [(3'h6):(1'h0)] reg1052 = (1'h0);
  reg [(3'h4):(1'h0)] reg1051 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1050 = (1'h0);
  reg [(4'h9):(1'h0)] reg1049 = (1'h0);
  reg [(3'h6):(1'h0)] reg1048 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1045 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1044 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1042 = (1'h0);
  reg [(2'h2):(1'h0)] reg1041 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1040 = (1'h0);
  reg [(4'ha):(1'h0)] reg1039 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1038 = (1'h0);
  reg [(2'h3):(1'h0)] reg1037 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1036 = (1'h0);
  reg [(2'h3):(1'h0)] reg1035 = (1'h0);
  reg [(4'hf):(1'h0)] reg1034 = (1'h0);
  reg [(2'h3):(1'h0)] reg1033 = (1'h0);
  reg [(3'h5):(1'h0)] reg1030 = (1'h0);
  reg [(2'h2):(1'h0)] reg1028 = (1'h0);
  reg [(3'h4):(1'h0)] reg1026 = (1'h0);
  reg [(4'hd):(1'h0)] reg1025 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1023 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1022 = (1'h0);
  reg [(4'he):(1'h0)] reg1021 = (1'h0);
  reg [(4'he):(1'h0)] reg1019 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1018 = (1'h0);
  reg [(3'h4):(1'h0)] reg1017 = (1'h0);
  reg [(4'hd):(1'h0)] reg1016 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1015 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1014 = (1'h0);
  reg [(4'hd):(1'h0)] reg1008 = (1'h0);
  reg [(4'ha):(1'h0)] reg1003 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1001 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg995 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg994 = (1'h0);
  reg [(3'h7):(1'h0)] reg1013 = (1'h0);
  reg [(2'h2):(1'h0)] reg1012 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1011 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1010 = (1'h0);
  reg [(4'he):(1'h0)] reg1009 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1007 = (1'h0);
  reg [(4'ha):(1'h0)] reg1006 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1005 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1004 = (1'h0);
  reg [(3'h5):(1'h0)] reg1002 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1000 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg999 = (1'h0);
  reg [(2'h3):(1'h0)] reg998 = (1'h0);
  reg [(3'h4):(1'h0)] reg997 = (1'h0);
  reg [(4'h8):(1'h0)] reg996 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg993 = (1'h0);
  reg [(2'h3):(1'h0)] reg992 = (1'h0);
  reg [(4'ha):(1'h0)] reg991 = (1'h0);
  reg [(4'h9):(1'h0)] reg990 = (1'h0);
  reg [(2'h3):(1'h0)] reg989 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1961 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1956 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1950 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1946 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1942 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1938 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1934 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1929 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1928 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1921 = (1'h0);
  reg [(4'he):(1'h0)] forvar1916 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1924 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1918 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1915 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1913 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1912 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1909 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1893 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1892 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1889 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1879 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1872 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1888 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1887 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1884 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1883 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1877 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1874 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1878 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1871 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1866 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1865 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1864 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1862 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1856 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1853 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1852 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1844 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1849 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1841 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1840 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1837 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1827 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1826 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1825 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1820 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1815 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1811 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1810 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1805 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1804 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1802 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1788 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1794 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1789 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1787 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1773 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1769 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1768 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1763 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1760 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1755 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1754 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1776 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1775 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1772 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1758 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1757 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1756 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1734 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1729 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1728 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1712 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1706 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1752 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1751 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1742 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1738 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1736 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1733 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1721 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1716 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1747 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1746 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1739 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1737 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1731 = (1'h0);
  reg [(4'he):(1'h0)] forvar1726 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1723 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1718 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1715 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1708 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1707 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1698 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1696 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1694 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1689 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1688 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1687 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1686 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1681 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1677 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1675 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1674 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1672 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1667 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1666 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1662 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1661 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1107 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1104 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1101 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1100 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1099 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1091 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1140 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1136 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1129 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1131 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1127 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1120 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1109 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1108 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1115 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1111 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1110 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1102 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1097 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1092 = (1'h0);
  reg [(4'he):(1'h0)] forvar1090 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1084 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1081 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1079 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1063 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1061 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1059 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1073 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1071 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1069 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1064 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1058 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1055 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1047 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1046 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1043 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1032 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1031 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1029 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1027 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1024 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1020 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1015 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1011 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1007 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1005 = (1'h0);
  reg [(4'ha):(1'h0)] forvar989 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1008 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1003 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1001 = (1'h0);
  reg [(2'h2):(1'h0)] forvar995 = (1'h0);
  reg [(4'he):(1'h0)] forvar994 = (1'h0);
  reg [(4'hb):(1'h0)] forvar990 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar988 = (1'h0);
  assign y = {wire1968,
                 wire1967,
                 wire1908,
                 wire1907,
                 wire1861,
                 wire1705,
                 wire986,
                 wire987,
                 wire1146,
                 wire1147,
                 wire1658,
                 reg1950,
                 reg1966,
                 reg1965,
                 reg1964,
                 reg1963,
                 reg1962,
                 reg1960,
                 reg1959,
                 reg1958,
                 reg1957,
                 reg1955,
                 reg1954,
                 reg1946,
                 reg1953,
                 reg1952,
                 reg1951,
                 reg1949,
                 reg1948,
                 reg1947,
                 reg1945,
                 reg1944,
                 reg1943,
                 reg1941,
                 reg1940,
                 reg1939,
                 reg1937,
                 reg1936,
                 reg1935,
                 reg1933,
                 reg1932,
                 reg1931,
                 reg1930,
                 reg1927,
                 reg1915,
                 reg1926,
                 reg1925,
                 reg1923,
                 reg1922,
                 reg1918,
                 reg1921,
                 reg1920,
                 reg1919,
                 reg1917,
                 reg1916,
                 reg1914,
                 reg1911,
                 reg1910,
                 reg1906,
                 reg1905,
                 reg1904,
                 reg1903,
                 reg1902,
                 reg1901,
                 reg1900,
                 reg1899,
                 reg1898,
                 reg1897,
                 reg1896,
                 reg1895,
                 reg1894,
                 reg1888,
                 reg1887,
                 reg1883,
                 reg1871,
                 reg1893,
                 reg1892,
                 reg1891,
                 reg1890,
                 reg1889,
                 reg1886,
                 reg1885,
                 reg1878,
                 reg1882,
                 reg1881,
                 reg1880,
                 reg1879,
                 reg1877,
                 reg1876,
                 reg1875,
                 reg1874,
                 reg1873,
                 reg1872,
                 reg1870,
                 reg1869,
                 reg1868,
                 reg1867,
                 reg1863,
                 reg1860,
                 reg1859,
                 reg1858,
                 reg1857,
                 reg1855,
                 reg1854,
                 reg1849,
                 reg1851,
                 reg1850,
                 reg1848,
                 reg1847,
                 reg1846,
                 reg1845,
                 reg1844,
                 reg1843,
                 reg1842,
                 reg1839,
                 reg1838,
                 reg1836,
                 reg1835,
                 reg1834,
                 reg1833,
                 reg1832,
                 reg1831,
                 reg1830,
                 reg1829,
                 reg1828,
                 reg1824,
                 reg1823,
                 reg1822,
                 reg1821,
                 reg1819,
                 reg1818,
                 reg1817,
                 reg1816,
                 reg1814,
                 reg1813,
                 reg1812,
                 reg1809,
                 reg1808,
                 reg1807,
                 reg1806,
                 reg1803,
                 reg1801,
                 reg1800,
                 reg1799,
                 reg1798,
                 reg1794,
                 reg1797,
                 reg1789,
                 reg1796,
                 reg1795,
                 reg1793,
                 reg1792,
                 reg1791,
                 reg1790,
                 reg1788,
                 reg1775,
                 reg1772,
                 reg1758,
                 reg1757,
                 reg1756,
                 reg1786,
                 reg1785,
                 reg1784,
                 reg1783,
                 reg1782,
                 reg1781,
                 reg1780,
                 reg1779,
                 reg1778,
                 reg1777,
                 reg1774,
                 reg1773,
                 reg1771,
                 reg1770,
                 reg1769,
                 reg1768,
                 reg1767,
                 reg1766,
                 reg1765,
                 reg1764,
                 reg1763,
                 reg1762,
                 reg1761,
                 reg1760,
                 reg1759,
                 reg1755,
                 reg1754,
                 reg1708,
                 reg1753,
                 reg1750,
                 reg1749,
                 reg1747,
                 reg1739,
                 reg1737,
                 reg1723,
                 reg1748,
                 reg1745,
                 reg1744,
                 reg1743,
                 reg1742,
                 reg1741,
                 reg1740,
                 reg1731,
                 reg1726,
                 reg1738,
                 reg1736,
                 reg1735,
                 reg1734,
                 reg1733,
                 reg1732,
                 reg1730,
                 reg1729,
                 reg1728,
                 reg1727,
                 reg1725,
                 reg1724,
                 reg1722,
                 reg1721,
                 reg1720,
                 reg1715,
                 reg1719,
                 reg1718,
                 reg1717,
                 reg1716,
                 reg1714,
                 reg1713,
                 reg1712,
                 reg1711,
                 reg1710,
                 reg1709,
                 reg1706,
                 reg1704,
                 reg1703,
                 reg1702,
                 reg1701,
                 reg1700,
                 reg1699,
                 reg1697,
                 reg1695,
                 reg1693,
                 reg1692,
                 reg1691,
                 reg1690,
                 reg1666,
                 reg1685,
                 reg1684,
                 reg1683,
                 reg1682,
                 reg1680,
                 reg1679,
                 reg1678,
                 reg1677,
                 reg1676,
                 reg1675,
                 reg1673,
                 reg1671,
                 reg1670,
                 reg1669,
                 reg1668,
                 reg1665,
                 reg1664,
                 reg1663,
                 reg1662,
                 reg1660,
                 reg1097,
                 reg1090,
                 reg1145,
                 reg1144,
                 reg1143,
                 reg1142,
                 reg1141,
                 reg1139,
                 reg1138,
                 reg1137,
                 reg1135,
                 reg1134,
                 reg1133,
                 reg1131,
                 reg1127,
                 reg1132,
                 reg1130,
                 reg1129,
                 reg1128,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1123,
                 reg1122,
                 reg1121,
                 reg1119,
                 reg1118,
                 reg1115,
                 reg1111,
                 reg1110,
                 reg1117,
                 reg1116,
                 reg1114,
                 reg1113,
                 reg1112,
                 reg1109,
                 reg1108,
                 reg1102,
                 reg1107,
                 reg1106,
                 reg1105,
                 reg1104,
                 reg1103,
                 reg1101,
                 reg1100,
                 reg1099,
                 reg1098,
                 reg1096,
                 reg1095,
                 reg1094,
                 reg1093,
                 reg1091,
                 reg1089,
                 reg1081,
                 reg1088,
                 reg1087,
                 reg1086,
                 reg1085,
                 reg1083,
                 reg1082,
                 reg1080,
                 reg1064,
                 reg1078,
                 reg1077,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg1072,
                 reg1058,
                 reg1070,
                 reg1068,
                 reg1067,
                 reg1066,
                 reg1065,
                 reg1063,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1057,
                 reg1056,
                 reg1027,
                 reg1054,
                 reg1053,
                 reg1052,
                 reg1051,
                 reg1050,
                 reg1049,
                 reg1048,
                 reg1045,
                 reg1044,
                 reg1042,
                 reg1041,
                 reg1040,
                 reg1039,
                 reg1038,
                 reg1037,
                 reg1036,
                 reg1035,
                 reg1034,
                 reg1033,
                 reg1030,
                 reg1028,
                 reg1026,
                 reg1025,
                 reg1023,
                 reg1022,
                 reg1021,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1016,
                 reg1015,
                 reg1014,
                 reg1008,
                 reg1003,
                 reg1001,
                 reg995,
                 reg994,
                 reg1013,
                 reg1012,
                 reg1011,
                 reg1010,
                 reg1009,
                 reg1007,
                 reg1006,
                 reg1005,
                 reg1004,
                 reg1002,
                 reg1000,
                 reg999,
                 reg998,
                 reg997,
                 reg996,
                 reg993,
                 reg992,
                 reg991,
                 reg990,
                 reg989,
                 forvar1961,
                 forvar1956,
                 forvar1950,
                 forvar1946,
                 forvar1942,
                 forvar1938,
                 forvar1934,
                 forvar1929,
                 forvar1928,
                 forvar1921,
                 forvar1916,
                 forvar1924,
                 forvar1918,
                 forvar1915,
                 forvar1913,
                 forvar1912,
                 forvar1909,
                 forvar1893,
                 forvar1892,
                 forvar1889,
                 forvar1879,
                 forvar1872,
                 forvar1888,
                 forvar1887,
                 forvar1884,
                 forvar1883,
                 forvar1877,
                 forvar1874,
                 forvar1878,
                 forvar1871,
                 forvar1866,
                 forvar1865,
                 forvar1864,
                 forvar1862,
                 forvar1856,
                 forvar1853,
                 forvar1852,
                 forvar1844,
                 forvar1849,
                 forvar1841,
                 forvar1840,
                 forvar1837,
                 forvar1827,
                 forvar1826,
                 forvar1825,
                 forvar1820,
                 forvar1815,
                 forvar1811,
                 forvar1810,
                 forvar1805,
                 forvar1804,
                 forvar1802,
                 forvar1788,
                 forvar1794,
                 forvar1789,
                 forvar1787,
                 forvar1773,
                 forvar1769,
                 forvar1768,
                 forvar1763,
                 forvar1760,
                 forvar1755,
                 forvar1754,
                 forvar1776,
                 forvar1775,
                 forvar1772,
                 forvar1758,
                 forvar1757,
                 forvar1756,
                 forvar1734,
                 forvar1729,
                 forvar1728,
                 forvar1712,
                 forvar1706,
                 forvar1752,
                 forvar1751,
                 forvar1742,
                 forvar1738,
                 forvar1736,
                 forvar1733,
                 forvar1721,
                 forvar1716,
                 forvar1747,
                 forvar1746,
                 forvar1739,
                 forvar1737,
                 forvar1731,
                 forvar1726,
                 forvar1723,
                 forvar1718,
                 forvar1715,
                 forvar1708,
                 forvar1707,
                 forvar1698,
                 forvar1696,
                 forvar1694,
                 forvar1689,
                 forvar1688,
                 forvar1687,
                 forvar1686,
                 forvar1681,
                 forvar1677,
                 forvar1675,
                 forvar1674,
                 forvar1672,
                 forvar1667,
                 forvar1666,
                 forvar1662,
                 forvar1661,
                 forvar1107,
                 forvar1104,
                 forvar1101,
                 forvar1100,
                 forvar1099,
                 forvar1091,
                 forvar1140,
                 forvar1136,
                 forvar1129,
                 forvar1131,
                 forvar1127,
                 forvar1120,
                 forvar1109,
                 forvar1108,
                 forvar1115,
                 forvar1111,
                 forvar1110,
                 forvar1102,
                 forvar1097,
                 forvar1092,
                 forvar1090,
                 forvar1084,
                 forvar1081,
                 forvar1079,
                 forvar1063,
                 forvar1061,
                 forvar1059,
                 forvar1073,
                 forvar1071,
                 forvar1069,
                 forvar1064,
                 forvar1058,
                 forvar1055,
                 forvar1047,
                 forvar1046,
                 forvar1043,
                 forvar1032,
                 forvar1031,
                 forvar1029,
                 forvar1027,
                 forvar1024,
                 forvar1020,
                 forvar1015,
                 forvar1011,
                 forvar1007,
                 forvar1005,
                 forvar989,
                 forvar1008,
                 forvar1003,
                 forvar1001,
                 forvar995,
                 forvar994,
                 forvar990,
                 forvar988,
                 (1'h0)};
  assign wire986 = wire985[(2'h2):(1'h1)];
  assign wire987 = (wire982 ?
                       $signed(((wire985 != wire984) - wire981[(4'h8):(1'h1)])) : (~&$signed((wire986 * wire981))));
  always
    @(posedge clk) begin
      for (forvar988 = (1'h0); (forvar988 < (1'h0)); forvar988 = (forvar988 + (1'h1)))
        begin
          if ($signed(({wire981} && $signed((wire983 ? forvar988 : wire986)))))
            begin
              if (wire986[(2'h3):(1'h1)])
                begin
                  reg989 <= (wire981[(4'ha):(2'h3)] ?
                      $signed($signed($unsigned(wire983))) : wire987);
                  if (((wire986[(2'h3):(2'h3)] ?
                          wire986[(1'h1):(1'h0)] : (~(~&reg989))) ?
                      $unsigned((-(-wire983))) : (wire981[(2'h2):(1'h0)] ?
                          $unsigned(wire986) : (~|wire982))))
                    begin
                      reg990 <= (($signed($signed(wire981)) >> (~|$unsigned((8'hb6)))) ?
                          wire982[(3'h5):(3'h4)] : $signed(wire984[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg990 <= $signed((~&$unsigned((wire987 + (8'hba)))));
                      reg991 <= ($unsigned(wire981) ?
                          {$signed($signed(wire982))} : (~&wire985[(1'h0):(1'h0)]));
                      reg992 <= ($signed(wire984) && (wire982[(4'ha):(1'h1)] ?
                          $signed(((8'ha3) && wire985)) : wire987[(3'h7):(3'h4)]));
                      reg993 <= ({(!(!wire985))} ?
                          {$unsigned(((8'hb9) ? reg989 : reg989))} : reg990);
                    end
                end
              else
                begin
                  reg989 <= (wire982 ?
                      (8'h9d) : $signed($unsigned((^~wire987))));
                  for (forvar990 = (1'h0); (forvar990 < (1'h0)); forvar990 = (forvar990 + (1'h1)))
                    begin
                      reg991 <= $unsigned(reg989);
                      reg992 <= (wire982 << reg989[(2'h3):(2'h3)]);
                      reg993 <= $unsigned(($signed({wire982}) == $unsigned(reg989[(2'h3):(2'h2)])));
                    end
                end
              for (forvar994 = (1'h0); (forvar994 < (1'h0)); forvar994 = (forvar994 + (1'h1)))
                begin
                  for (forvar995 = (1'h0); (forvar995 < (2'h2)); forvar995 = (forvar995 + (1'h1)))
                    begin
                      reg996 <= (^~$unsigned(((~^wire985) ?
                          (forvar994 ?
                              wire987 : forvar994) : $unsigned(forvar988))));
                      reg997 <= ({reg993} ?
                          $signed(($signed(wire982) < (wire987 ?
                              wire981 : wire981))) : $unsigned(reg991));
                    end
                  if (((~|$signed($unsigned(forvar994))) ?
                      forvar995 : $signed((8'had))))
                    begin
                      reg998 <= ($unsigned($signed((+forvar990))) ?
                          {$unsigned(reg990[(3'h5):(3'h4)])} : wire986[(1'h0):(1'h0)]);
                      reg999 <= (~reg989[(2'h3):(1'h1)]);
                      reg1000 <= {$signed((!reg999))};
                    end
                  else
                    begin
                      reg998 <= reg991;
                      reg999 <= (!(~&wire987));
                    end
                end
              for (forvar1001 = (1'h0); (forvar1001 < (1'h1)); forvar1001 = (forvar1001 + (1'h1)))
                begin
                  reg1002 <= {$signed((wire983[(3'h6):(2'h3)] | (^(8'ha4))))};
                  for (forvar1003 = (1'h0); (forvar1003 < (1'h0)); forvar1003 = (forvar1003 + (1'h1)))
                    begin
                      reg1004 <= reg1002[(3'h4):(2'h2)];
                      reg1005 <= (^(~&(+$signed((8'hb3)))));
                      reg1006 <= forvar990;
                      reg1007 <= (|($signed(wire987) ?
                          forvar995 : (wire986 - (&reg993))));
                    end
                  for (forvar1008 = (1'h0); (forvar1008 < (1'h1)); forvar1008 = (forvar1008 + (1'h1)))
                    begin
                      reg1009 <= reg991[(4'h9):(1'h0)];
                      reg1010 <= (forvar1008[(3'h7):(3'h4)] ~^ reg991[(3'h7):(2'h2)]);
                      reg1011 <= (($unsigned($unsigned(forvar1001)) ?
                          reg1000[(1'h1):(1'h0)] : $unsigned(reg991)) >> forvar1001[(4'h9):(3'h7)]);
                    end
                  if ($unsigned((-(^forvar995[(1'h1):(1'h0)]))))
                    begin
                      reg1012 <= (forvar995 ?
                          (+$unsigned(reg997)) : ({reg1005} ?
                              reg1000[(3'h5):(1'h1)] : (8'had)));
                    end
                  else
                    begin
                      reg1012 <= reg1004;
                      reg1013 <= $signed(reg1009);
                    end
                end
            end
          else
            begin
              for (forvar989 = (1'h0); (forvar989 < (1'h0)); forvar989 = (forvar989 + (1'h1)))
                begin
                  for (forvar990 = (1'h0); (forvar990 < (2'h3)); forvar990 = (forvar990 + (1'h1)))
                    begin
                      reg991 <= wire984[(1'h1):(1'h0)];
                    end
                  if ({reg1011})
                    begin
                      reg992 <= wire986;
                      reg993 <= (reg1002 && forvar994[(4'ha):(4'h9)]);
                      reg994 <= $unsigned(forvar1008[(1'h0):(1'h0)]);
                      reg995 <= $signed((!{reg1005}));
                    end
                  else
                    begin
                      reg992 <= reg1012[(1'h1):(1'h0)];
                    end
                  if ((~&reg997))
                    begin
                      reg996 <= (reg1005 ?
                          wire983 : $signed($unsigned((~^reg1007))));
                      reg997 <= $unsigned(forvar988);
                      reg998 <= (~(((!reg997) ?
                              (reg997 ^~ reg998) : (wire983 && forvar1008)) ?
                          $signed({(8'ha5)}) : {$unsigned(forvar994)}));
                      reg999 <= (~&($signed(forvar1001) + wire985[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg996 <= (!reg1010[(4'hb):(2'h3)]);
                      reg997 <= {($signed((reg1006 + (8'hb1))) > wire987)};
                      reg998 <= (~|$unsigned($signed($unsigned((8'hae)))));
                    end
                  if ((reg1004 >>> ((reg1004[(3'h6):(2'h3)] << $signed((8'hb7))) == reg1009[(2'h2):(1'h1)])))
                    begin
                      reg1000 <= ($unsigned(((~(8'h9d)) ?
                          (-wire982) : wire985)) || ((~&(reg998 == forvar1008)) ?
                          ({forvar1008} >>> wire985[(3'h4):(2'h2)]) : (|(forvar988 & reg992))));
                      reg1001 <= $unsigned(reg1013[(3'h4):(3'h4)]);
                      reg1002 <= $unsigned(reg994);
                      reg1003 <= ($unsigned(((8'ha3) ?
                              $signed(forvar1008) : (^~forvar1003))) ?
                          (wire981[(4'he):(4'hd)] && $signed($unsigned(reg1009))) : ($signed((forvar1001 ?
                              reg992 : (8'ha1))) ~^ $unsigned((8'hab))));
                    end
                  else
                    begin
                      reg1000 <= {$signed($unsigned($unsigned(reg990)))};
                    end
                end
              reg1004 <= $signed((^(-(reg1003 ? reg989 : reg1001))));
              if (forvar1008)
                begin
                  for (forvar1005 = (1'h0); (forvar1005 < (1'h0)); forvar1005 = (forvar1005 + (1'h1)))
                    begin
                      reg1006 <= ({(wire984 ^ (reg1013 ?
                              forvar1003 : reg999))} ^~ reg1005);
                    end
                  for (forvar1007 = (1'h0); (forvar1007 < (2'h2)); forvar1007 = (forvar1007 + (1'h1)))
                    begin
                      reg1008 <= $unsigned(($unsigned(reg997) << forvar988));
                      reg1009 <= ((!{(^reg991)}) ?
                          $signed({$unsigned(reg992)}) : reg999);
                      reg1010 <= $signed($unsigned(((&reg1006) ?
                          (reg998 ? (8'hb2) : reg997) : reg990)));
                    end
                end
              else
                begin
                  if (((~|({(8'hb7)} >>> (|(8'hb7)))) * (forvar1008 ?
                      ((reg1012 <<< reg1003) < $signed(reg1012)) : forvar995)))
                    begin
                      reg1005 <= $signed((forvar989 != $signed($signed(reg993))));
                      reg1006 <= $signed({$signed((~^reg1007))});
                      reg1007 <= (^$signed($signed(reg1006[(3'h6):(1'h0)])));
                    end
                  else
                    begin
                      reg1005 <= (!forvar990);
                      reg1006 <= forvar989;
                      reg1007 <= $signed(reg1004[(4'he):(4'he)]);
                      reg1008 <= (reg1002 + forvar1005[(3'h5):(2'h2)]);
                    end
                end
              if ((8'hac))
                begin
                  for (forvar1011 = (1'h0); (forvar1011 < (1'h1)); forvar1011 = (forvar1011 + (1'h1)))
                    begin
                      reg1012 <= $signed($signed($unsigned(wire986[(3'h4):(1'h0)])));
                      reg1013 <= (((8'h9e) <= (reg990 ~^ reg1003)) < forvar989);
                      reg1014 <= $signed(forvar1007);
                      reg1015 <= (~(({forvar1008} ^~ $unsigned(wire981)) ?
                          (~(&reg1001)) : $unsigned((^(8'ha8)))));
                    end
                end
              else
                begin
                  if (((|((^(8'ha3)) || reg1015)) >= ($signed((~forvar1007)) ?
                      {(&forvar1008)} : wire982)))
                    begin
                      reg1011 <= reg999[(3'h4):(2'h2)];
                      reg1012 <= reg999[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1011 <= {(((&reg1015) ?
                              (reg989 ^~ reg994) : ((8'hb5) ?
                                  forvar988 : (8'haa))) * ((forvar994 != (8'hb3)) ?
                              wire984 : $signed(reg998)))};
                      reg1012 <= (forvar1011 ?
                          $signed({$unsigned(wire984)}) : reg1009[(3'h4):(3'h4)]);
                      reg1013 <= {$unsigned(wire983)};
                      reg1014 <= forvar1008;
                    end
                  for (forvar1015 = (1'h0); (forvar1015 < (1'h0)); forvar1015 = (forvar1015 + (1'h1)))
                    begin
                      reg1016 <= reg1015;
                      reg1017 <= {(+(8'hb7))};
                      reg1018 <= reg1012[(1'h1):(1'h0)];
                      reg1019 <= {{((8'h9c) >> (reg1009 ? (8'ha0) : (8'had)))}};
                    end
                  for (forvar1020 = (1'h0); (forvar1020 < (1'h1)); forvar1020 = (forvar1020 + (1'h1)))
                    begin
                      reg1021 <= {$unsigned(($signed(reg993) ?
                              wire982[(3'h6):(1'h0)] : forvar994[(3'h7):(3'h5)]))};
                      reg1022 <= reg1007;
                      reg1023 <= reg989;
                    end
                  for (forvar1024 = (1'h0); (forvar1024 < (1'h1)); forvar1024 = (forvar1024 + (1'h1)))
                    begin
                      reg1025 <= (~|(reg1002 ?
                          (reg1023 ^ $signed(forvar1001)) : ((8'hb3) >> $unsigned(forvar1007))));
                      reg1026 <= $unsigned(reg1013);
                    end
                end
            end
          if (reg1022)
            begin
              for (forvar1027 = (1'h0); (forvar1027 < (2'h2)); forvar1027 = (forvar1027 + (1'h1)))
                begin
                  reg1028 <= reg1019[(2'h3):(2'h2)];
                  for (forvar1029 = (1'h0); (forvar1029 < (1'h0)); forvar1029 = (forvar1029 + (1'h1)))
                    begin
                      reg1030 <= reg1021[(2'h2):(2'h2)];
                    end
                end
              for (forvar1031 = (1'h0); (forvar1031 < (2'h2)); forvar1031 = (forvar1031 + (1'h1)))
                begin
                  for (forvar1032 = (1'h0); (forvar1032 < (1'h0)); forvar1032 = (forvar1032 + (1'h1)))
                    begin
                      reg1033 <= (8'hb2);
                      reg1034 <= reg1006;
                      reg1035 <= reg1003[(3'h7):(1'h1)];
                      reg1036 <= reg1018;
                    end
                  if ($signed((8'ha5)))
                    begin
                      reg1037 <= reg1003;
                    end
                  else
                    begin
                      reg1037 <= reg991[(1'h1):(1'h1)];
                      reg1038 <= ((-$unsigned({reg1033})) ?
                          (|{((8'haa) ~^ reg991)}) : (((reg991 + wire982) <= (reg1035 ^ reg1010)) ?
                              (reg993 ?
                                  (reg999 && reg1036) : $unsigned(reg1016)) : (~$unsigned(reg1011))));
                    end
                  if ($unsigned({$signed($signed(reg1019))}))
                    begin
                      reg1039 <= (8'hb3);
                      reg1040 <= (reg1033 >= $signed($unsigned(forvar995[(2'h2):(2'h2)])));
                      reg1041 <= (reg1003 ^~ reg1035[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1039 <= reg1007[(2'h2):(1'h1)];
                      reg1040 <= (^~($signed(reg1014[(2'h3):(1'h0)]) | $unsigned($signed(reg1007))));
                      reg1041 <= reg1000;
                      reg1042 <= forvar988;
                    end
                  for (forvar1043 = (1'h0); (forvar1043 < (2'h3)); forvar1043 = (forvar1043 + (1'h1)))
                    begin
                      reg1044 <= reg1006;
                      reg1045 <= $signed($signed(forvar1020));
                    end
                end
              for (forvar1046 = (1'h0); (forvar1046 < (2'h2)); forvar1046 = (forvar1046 + (1'h1)))
                begin
                  for (forvar1047 = (1'h0); (forvar1047 < (1'h0)); forvar1047 = (forvar1047 + (1'h1)))
                    begin
                      reg1048 <= (8'hb2);
                      reg1049 <= wire983[(3'h4):(1'h0)];
                      reg1050 <= (~|(-(|forvar990)));
                      reg1051 <= (|forvar988);
                    end
                  if ($unsigned($unsigned($signed((8'had)))))
                    begin
                      reg1052 <= reg1041[(1'h0):(1'h0)];
                      reg1053 <= $unsigned(forvar1008[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg1052 <= reg1030;
                      reg1053 <= reg989[(2'h3):(2'h3)];
                      reg1054 <= ($signed(wire983) ~^ {(8'hae)});
                    end
                end
            end
          else
            begin
              reg1027 <= $unsigned((^{reg1000}));
            end
          if (($unsigned(((reg1008 <= reg1001) <= reg1000[(2'h3):(1'h0)])) || (8'hb4)))
            begin
              if ((!$unsigned(wire982)))
                begin
                  for (forvar1055 = (1'h0); (forvar1055 < (1'h1)); forvar1055 = (forvar1055 + (1'h1)))
                    begin
                      reg1056 <= reg1018;
                      reg1057 <= ($signed($signed(reg998)) >>> (reg1006[(2'h3):(2'h3)] && (!forvar1020[(2'h2):(1'h1)])));
                    end
                end
              else
                begin
                  for (forvar1055 = (1'h0); (forvar1055 < (2'h3)); forvar1055 = (forvar1055 + (1'h1)))
                    begin
                      reg1056 <= (reg1036[(1'h0):(1'h0)] || (({(8'h9e)} ?
                          (forvar1027 >> forvar1032) : $signed(forvar988)) || wire984[(1'h0):(1'h0)]));
                    end
                end
              if (reg1033)
                begin
                  for (forvar1058 = (1'h0); (forvar1058 < (1'h1)); forvar1058 = (forvar1058 + (1'h1)))
                    begin
                      reg1059 <= $signed(reg989);
                    end
                  if ((reg1023[(2'h3):(1'h1)] ~^ $unsigned(reg1052[(2'h3):(1'h1)])))
                    begin
                      reg1060 <= reg1041[(1'h0):(1'h0)];
                      reg1061 <= wire982;
                      reg1062 <= (-reg1038[(2'h3):(2'h2)]);
                      reg1063 <= ((~$signed((reg1030 >> reg1060))) >>> reg1042[(4'h8):(4'h8)]);
                    end
                  else
                    begin
                      reg1060 <= ($signed((8'hb3)) ?
                          $signed((8'ha7)) : (reg998[(1'h1):(1'h0)] ?
                              ((reg1057 ? forvar1047 : reg1027) ?
                                  ((8'h9f) && reg992) : $signed(forvar1003)) : $signed((reg989 ?
                                  forvar1055 : reg1013))));
                    end
                  for (forvar1064 = (1'h0); (forvar1064 < (2'h3)); forvar1064 = (forvar1064 + (1'h1)))
                    begin
                      reg1065 <= (8'hac);
                      reg1066 <= (~^forvar1007);
                      reg1067 <= $unsigned($signed(reg1019[(4'he):(2'h2)]));
                      reg1068 <= {(!$unsigned($unsigned(reg1034)))};
                    end
                  for (forvar1069 = (1'h0); (forvar1069 < (1'h1)); forvar1069 = (forvar1069 + (1'h1)))
                    begin
                      reg1070 <= $unsigned($unsigned(reg995[(2'h2):(1'h0)]));
                    end
                end
              else
                begin
                  reg1058 <= reg1050;
                end
              for (forvar1071 = (1'h0); (forvar1071 < (2'h2)); forvar1071 = (forvar1071 + (1'h1)))
                begin
                  reg1072 <= reg1038;
                  for (forvar1073 = (1'h0); (forvar1073 < (2'h2)); forvar1073 = (forvar1073 + (1'h1)))
                    begin
                      reg1074 <= ($signed((+(!wire985))) & (forvar1046 ^~ $signed(reg1010)));
                      reg1075 <= reg998;
                      reg1076 <= reg1049[(3'h7):(3'h4)];
                    end
                  if ($unsigned(($signed($signed(forvar1069)) == ((forvar1064 ?
                      forvar988 : reg1023) ^ (~(8'ha0))))))
                    begin
                      reg1077 <= (^forvar1055);
                      reg1078 <= ($signed({reg1022[(1'h1):(1'h0)]}) ?
                          reg1056 : (~|$signed($signed(reg1063))));
                    end
                  else
                    begin
                      reg1077 <= (~(($unsigned(reg1013) ^~ (reg1051 ~^ reg1018)) ?
                          {$unsigned(reg1022)} : ($signed(reg1014) ?
                              {(8'ha3)} : (reg1021 <= (8'hb4)))));
                      reg1078 <= reg992[(2'h2):(1'h1)];
                    end
                end
            end
          else
            begin
              for (forvar1055 = (1'h0); (forvar1055 < (2'h2)); forvar1055 = (forvar1055 + (1'h1)))
                begin
                  if (($signed({forvar1031}) && (((reg1028 >>> (8'ha7)) || (reg1008 >> forvar995)) ?
                      reg1074 : reg1038)))
                    begin
                      reg1056 <= $signed($signed({forvar988[(1'h0):(1'h0)]}));
                      reg1057 <= reg1054;
                    end
                  else
                    begin
                      reg1056 <= $signed($signed(({reg1030} ?
                          ((8'h9f) << reg1005) : (reg1037 * reg1015))));
                      reg1057 <= (-(!$unsigned(reg1037[(2'h2):(1'h1)])));
                      reg1058 <= wire986;
                    end
                end
              for (forvar1059 = (1'h0); (forvar1059 < (1'h0)); forvar1059 = (forvar1059 + (1'h1)))
                begin
                  if ({$signed($signed((&forvar1047)))})
                    begin
                      reg1060 <= $signed(reg1061);
                    end
                  else
                    begin
                      reg1060 <= $signed({(^~$signed(reg1050))});
                    end
                  for (forvar1061 = (1'h0); (forvar1061 < (2'h2)); forvar1061 = (forvar1061 + (1'h1)))
                    begin
                      reg1062 <= reg997;
                    end
                  for (forvar1063 = (1'h0); (forvar1063 < (2'h2)); forvar1063 = (forvar1063 + (1'h1)))
                    begin
                      reg1064 <= (+(^~reg995[(1'h0):(1'h0)]));
                    end
                  reg1065 <= ($signed($signed($signed((8'hae)))) ?
                      $unsigned(forvar1003[(2'h3):(2'h2)]) : reg1018[(2'h2):(1'h1)]);
                end
            end
          for (forvar1079 = (1'h0); (forvar1079 < (2'h3)); forvar1079 = (forvar1079 + (1'h1)))
            begin
              if ((^~(8'ha8)))
                begin
                  reg1080 <= $unsigned($unsigned({(reg1035 - (8'hb7))}));
                  for (forvar1081 = (1'h0); (forvar1081 < (1'h1)); forvar1081 = (forvar1081 + (1'h1)))
                    begin
                      reg1082 <= forvar1063;
                      reg1083 <= $signed(({(~^forvar1073)} ?
                          $signed({reg1019}) : {forvar1011[(3'h4):(2'h3)]}));
                    end
                  for (forvar1084 = (1'h0); (forvar1084 < (1'h0)); forvar1084 = (forvar1084 + (1'h1)))
                    begin
                      reg1085 <= $unsigned(forvar1071);
                      reg1086 <= (+(~^forvar1043[(4'hc):(2'h2)]));
                      reg1087 <= ($unsigned((^~(forvar1032 ?
                              reg1061 : forvar1024))) ?
                          ($signed((8'ha3)) & (~&(reg1063 ~^ (8'hba)))) : $unsigned($unsigned((reg1060 >= reg1051))));
                    end
                  if ($signed((($signed(forvar1031) ?
                      (reg1085 ?
                          reg1060 : reg1062) : ((8'hb7) << reg1061)) <= $unsigned((|reg1026)))))
                    begin
                      reg1088 <= $unsigned(((&reg1005[(3'h7):(2'h3)]) * $unsigned({reg989})));
                    end
                  else
                    begin
                      reg1088 <= (forvar1046 ? (8'haa) : reg1044);
                    end
                end
              else
                begin
                  if (reg1033)
                    begin
                      reg1080 <= {(($unsigned(reg1007) ^ $unsigned(forvar1061)) ?
                              ((8'ha6) ?
                                  (reg1037 && reg1011) : $unsigned(reg1054)) : (^(8'haf)))};
                      reg1081 <= reg1087;
                    end
                  else
                    begin
                      reg1080 <= $unsigned(forvar1001[(5'h10):(4'h9)]);
                      reg1081 <= $unsigned((&((reg1050 * reg1085) ?
                          (8'hb7) : $unsigned((8'h9c)))));
                      reg1082 <= $signed(reg1023[(2'h2):(1'h1)]);
                      reg1083 <= (^~{(reg1056 ? $signed(reg999) : forvar1071)});
                    end
                end
              reg1089 <= ($unsigned((~(reg1037 ? reg1082 : reg1019))) ?
                  $signed(reg1050[(3'h4):(1'h1)]) : $unsigned(((&forvar1079) ?
                      $unsigned(reg1030) : $unsigned(reg1077))));
            end
        end
      if ($signed((8'hb7)))
        begin
          for (forvar1090 = (1'h0); (forvar1090 < (2'h3)); forvar1090 = (forvar1090 + (1'h1)))
            begin
              reg1091 <= {reg1052[(1'h1):(1'h0)]};
              for (forvar1092 = (1'h0); (forvar1092 < (2'h2)); forvar1092 = (forvar1092 + (1'h1)))
                begin
                  if ((8'hb3))
                    begin
                      reg1093 <= $unsigned(((wire982 && $unsigned(reg1039)) ?
                          (-reg992) : (~|reg1013[(3'h5):(3'h4)])));
                      reg1094 <= (reg992[(2'h3):(2'h3)] ?
                          $unsigned(($signed(reg1034) ?
                              (forvar1032 ?
                                  forvar1011 : reg1057) : (&reg1041))) : (((forvar1003 ?
                                      reg1081 : forvar1020) ?
                                  $unsigned(reg1080) : (reg1067 ?
                                      (8'hb3) : reg1048)) ?
                              reg994[(1'h1):(1'h1)] : {reg1048[(3'h4):(1'h1)]}));
                      reg1095 <= reg1025[(4'h9):(4'h9)];
                    end
                  else
                    begin
                      reg1093 <= {(|reg1004[(4'hb):(4'hb)])};
                      reg1094 <= $signed($unsigned($unsigned((forvar1031 == reg1013))));
                      reg1095 <= (((~&$signed(wire984)) <<< forvar1061) & $unsigned(reg997[(3'h4):(3'h4)]));
                      reg1096 <= reg997[(2'h3):(1'h1)];
                    end
                  for (forvar1097 = (1'h0); (forvar1097 < (1'h1)); forvar1097 = (forvar1097 + (1'h1)))
                    begin
                      reg1098 <= $signed((($signed((8'ha8)) ?
                              $signed((8'h9e)) : ((8'hac) ?
                                  reg1044 : forvar1092)) ?
                          ((reg1057 ? reg1008 : reg1056) ?
                              forvar1024 : (~|reg1063)) : (~^$signed(reg991))));
                      reg1099 <= (^(^~(!(~&reg1064))));
                      reg1100 <= ((reg1050[(4'h8):(4'h8)] || {reg1027}) - $signed($signed(reg1095)));
                      reg1101 <= $signed(wire983[(1'h0):(1'h0)]);
                    end
                end
            end
          if (reg1002)
            begin
              for (forvar1102 = (1'h0); (forvar1102 < (2'h2)); forvar1102 = (forvar1102 + (1'h1)))
                begin
                  if ($unsigned($signed($signed((reg1037 >> forvar1011)))))
                    begin
                      reg1103 <= (reg995 ?
                          (^(~&(reg989 ?
                              reg1044 : reg1100))) : forvar1001[(3'h7):(3'h4)]);
                    end
                  else
                    begin
                      reg1103 <= ($unsigned(reg996[(2'h3):(2'h2)]) ?
                          (($unsigned(forvar1032) ?
                                  reg1006[(3'h4):(2'h2)] : reg1066) ?
                              $unsigned(((8'hab) >> reg1033)) : $signed(((8'haf) < reg1022))) : reg1010[(4'hb):(3'h4)]);
                    end
                  if (forvar1069[(3'h4):(1'h0)])
                    begin
                      reg1104 <= ($unsigned(((forvar988 * reg1100) <<< reg1064)) ?
                          $signed($unsigned($signed(reg1025))) : forvar1102);
                      reg1105 <= ((8'hb8) && reg1089[(4'hc):(3'h5)]);
                      reg1106 <= (+(|(~^(reg1101 ? reg1041 : reg998))));
                      reg1107 <= forvar989[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg1104 <= reg1064;
                      reg1105 <= $signed(reg1016[(4'ha):(4'h8)]);
                      reg1106 <= (8'ha4);
                      reg1107 <= forvar990[(3'h6):(2'h3)];
                    end
                end
            end
          else
            begin
              reg1102 <= reg996;
            end
          if (reg1082)
            begin
              reg1108 <= forvar990;
              reg1109 <= forvar988;
              for (forvar1110 = (1'h0); (forvar1110 < (1'h0)); forvar1110 = (forvar1110 + (1'h1)))
                begin
                  for (forvar1111 = (1'h0); (forvar1111 < (1'h1)); forvar1111 = (forvar1111 + (1'h1)))
                    begin
                      reg1112 <= (|$unsigned((+(forvar1058 ?
                          forvar995 : forvar1043))));
                      reg1113 <= (reg1004 == reg1061[(3'h5):(2'h3)]);
                      reg1114 <= reg1014;
                    end
                  for (forvar1115 = (1'h0); (forvar1115 < (2'h2)); forvar1115 = (forvar1115 + (1'h1)))
                    begin
                      reg1116 <= (^reg995[(2'h3):(2'h3)]);
                    end
                  reg1117 <= (~forvar1097[(3'h7):(3'h7)]);
                end
            end
          else
            begin
              for (forvar1108 = (1'h0); (forvar1108 < (1'h0)); forvar1108 = (forvar1108 + (1'h1)))
                begin
                  for (forvar1109 = (1'h0); (forvar1109 < (2'h3)); forvar1109 = (forvar1109 + (1'h1)))
                    begin
                      reg1110 <= reg998[(2'h2):(2'h2)];
                      reg1111 <= reg1013[(3'h7):(3'h7)];
                    end
                  if ((reg1076[(2'h3):(2'h2)] ^ $signed(forvar1073[(3'h6):(3'h5)])))
                    begin
                      reg1112 <= {{((!reg1096) ? (+reg1005) : (!(8'ha9)))}};
                    end
                  else
                    begin
                      reg1112 <= forvar1102;
                      reg1113 <= $unsigned($signed({(~forvar994)}));
                    end
                  reg1114 <= forvar1055;
                  if (({(-(-reg1010))} << (reg1012 ?
                      (^~(reg1117 ~^ reg1117)) : (^((8'ha4) <<< (8'ha0))))))
                    begin
                      reg1115 <= $unsigned(reg1062[(3'h4):(2'h2)]);
                      reg1116 <= (8'hb4);
                      reg1117 <= {forvar1071[(5'h10):(4'h9)]};
                      reg1118 <= forvar1079;
                    end
                  else
                    begin
                      reg1115 <= ((~reg1095[(3'h5):(3'h4)]) ?
                          forvar1108[(2'h3):(2'h2)] : {reg1057});
                      reg1116 <= reg1056;
                      reg1117 <= forvar1081;
                      reg1118 <= reg1049[(4'h8):(3'h6)];
                    end
                end
              reg1119 <= (^(^~((~&reg1009) > reg1053[(2'h2):(1'h0)])));
            end
          for (forvar1120 = (1'h0); (forvar1120 < (1'h1)); forvar1120 = (forvar1120 + (1'h1)))
            begin
              if ((&(-$signed($unsigned(reg1117)))))
                begin
                  if (reg1088[(3'h5):(3'h5)])
                    begin
                      reg1121 <= (&($signed((8'had)) <= (~^reg1107[(1'h1):(1'h1)])));
                      reg1122 <= ($signed($unsigned(reg1018)) >> $unsigned($unsigned((8'hb3))));
                    end
                  else
                    begin
                      reg1121 <= (8'ha6);
                    end
                  if ($unsigned($signed((reg1000 ?
                      (~^reg997) : (reg996 ? (8'ha2) : forvar1110)))))
                    begin
                      reg1123 <= ($signed((&$signed(reg997))) << $unsigned(reg998));
                    end
                  else
                    begin
                      reg1123 <= $signed({(!((8'hb5) ? reg1028 : forvar1108))});
                      reg1124 <= {$signed(reg1095)};
                      reg1125 <= {((~^(~|reg998)) ?
                              {reg1075} : ((+reg1100) & {reg1054}))};
                      reg1126 <= reg1044[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  if ((&{((!forvar1047) ? forvar1081 : $unsigned((8'hac)))}))
                    begin
                      reg1121 <= (reg1003 || (($unsigned(reg1066) ?
                              forvar1115[(2'h2):(1'h0)] : (reg1067 >= reg1023)) ?
                          $unsigned(reg1042) : reg1006));
                    end
                  else
                    begin
                      reg1121 <= (reg997 > $signed(reg1056[(1'h1):(1'h0)]));
                      reg1122 <= {(~reg999)};
                      reg1123 <= forvar1102;
                    end
                end
              if ($signed($unsigned((~^{reg1113}))))
                begin
                  for (forvar1127 = (1'h0); (forvar1127 < (1'h1)); forvar1127 = (forvar1127 + (1'h1)))
                    begin
                      reg1128 <= forvar1011[(4'ha):(3'h6)];
                      reg1129 <= reg1033;
                      reg1130 <= (~|$unsigned($signed(reg1067[(4'h9):(3'h5)])));
                    end
                  for (forvar1131 = (1'h0); (forvar1131 < (1'h0)); forvar1131 = (forvar1131 + (1'h1)))
                    begin
                      reg1132 <= $signed((^~$signed($signed((8'hae)))));
                    end
                end
              else
                begin
                  if (($unsigned((8'hb5)) ?
                      (reg1066[(2'h2):(1'h0)] ?
                          ($unsigned(reg1081) ?
                              (reg1121 ~^ reg1105) : (reg1027 ?
                                  reg1010 : reg1039)) : reg1123[(2'h3):(2'h3)]) : $signed((~&reg1062))))
                    begin
                      reg1127 <= $unsigned(reg998[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1127 <= {($unsigned((~forvar1109)) ?
                              (&wire986) : ($signed((8'ha6)) ~^ reg1051))};
                    end
                  if ($unsigned(reg1118))
                    begin
                      reg1128 <= ($signed($signed((reg1061 ?
                          reg1014 : reg1107))) << (reg1003 ?
                          forvar1081[(1'h0):(1'h0)] : reg1080[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg1128 <= $signed({(reg1114 ?
                              (reg1100 ? forvar1131 : reg1123) : {reg1105})});
                    end
                  for (forvar1129 = (1'h0); (forvar1129 < (1'h1)); forvar1129 = (forvar1129 + (1'h1)))
                    begin
                      reg1130 <= ($unsigned((8'hb0)) ?
                          $unsigned(((reg1039 ? reg1044 : reg1002) ?
                              $signed(forvar1127) : reg1081)) : ({reg1118} >>> reg1054[(3'h7):(3'h5)]));
                      reg1131 <= $unsigned({((forvar1127 > reg1091) ?
                              (|forvar1120) : reg1042[(4'hd):(4'hb)])});
                    end
                  if (reg1026)
                    begin
                      reg1132 <= $unsigned(reg1076[(3'h4):(3'h4)]);
                      reg1133 <= $unsigned((({reg1003} ?
                          (reg1050 == reg991) : $unsigned(reg989)) ~^ $signed($signed(forvar1029))));
                    end
                  else
                    begin
                      reg1132 <= $signed(reg1132);
                      reg1133 <= {forvar988};
                      reg1134 <= (reg1076[(4'h8):(2'h3)] ?
                          (~((forvar1015 ?
                              (8'hba) : (8'hb2)) & reg1018)) : (reg993 >> forvar1079[(1'h1):(1'h1)]));
                      reg1135 <= reg1077[(3'h4):(2'h2)];
                    end
                end
              for (forvar1136 = (1'h0); (forvar1136 < (1'h0)); forvar1136 = (forvar1136 + (1'h1)))
                begin
                  if ((^$signed($signed($signed(forvar1058)))))
                    begin
                      reg1137 <= (8'hba);
                      reg1138 <= reg1056;
                      reg1139 <= $unsigned($signed(reg1133));
                    end
                  else
                    begin
                      reg1137 <= reg993;
                    end
                end
              for (forvar1140 = (1'h0); (forvar1140 < (1'h0)); forvar1140 = (forvar1140 + (1'h1)))
                begin
                  if ($signed((($signed(reg1080) ?
                          $unsigned(reg1086) : reg1019) ?
                      $unsigned((+forvar994)) : reg1082)))
                    begin
                      reg1141 <= ($signed(((8'ha4) || reg1050)) ?
                          reg1062 : (!forvar1059[(2'h3):(1'h1)]));
                      reg1142 <= reg994[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1141 <= reg1103;
                      reg1142 <= $signed($unsigned((((8'h9d) >>> reg1040) ?
                          ((8'hb2) & forvar1129) : reg1139)));
                      reg1143 <= reg1070[(2'h2):(1'h1)];
                    end
                  reg1144 <= {$signed($signed((reg1012 ? reg1083 : reg1042)))};
                  if ($signed(forvar1136[(1'h1):(1'h1)]))
                    begin
                      reg1145 <= (8'hb9);
                    end
                  else
                    begin
                      reg1145 <= reg1014[(1'h1):(1'h0)];
                    end
                end
            end
        end
      else
        begin
          reg1090 <= forvar1064;
          for (forvar1091 = (1'h0); (forvar1091 < (1'h0)); forvar1091 = (forvar1091 + (1'h1)))
            begin
              for (forvar1092 = (1'h0); (forvar1092 < (1'h0)); forvar1092 = (forvar1092 + (1'h1)))
                begin
                  reg1093 <= (forvar1027 ?
                      $signed(reg1110[(3'h4):(1'h1)]) : $signed((8'hb6)));
                  if ($unsigned(($unsigned($signed(reg995)) ?
                      {(reg1014 | forvar1071)} : reg1012[(2'h2):(1'h0)])))
                    begin
                      reg1094 <= {reg1070[(2'h2):(1'h0)]};
                      reg1095 <= (reg1042[(3'h4):(1'h0)] & (^reg1044[(2'h2):(2'h2)]));
                      reg1096 <= (~|(!$signed(((8'h9f) || (8'hb4)))));
                      reg1097 <= {(-(~&$signed(reg1109)))};
                    end
                  else
                    begin
                      reg1094 <= $signed(forvar1097[(4'h8):(3'h4)]);
                      reg1095 <= ((-reg1122) == (~|((8'hb4) ?
                          (reg1099 << reg997) : $signed(reg1083))));
                    end
                end
              reg1098 <= forvar1061;
            end
          for (forvar1099 = (1'h0); (forvar1099 < (2'h2)); forvar1099 = (forvar1099 + (1'h1)))
            begin
              for (forvar1100 = (1'h0); (forvar1100 < (2'h3)); forvar1100 = (forvar1100 + (1'h1)))
                begin
                  for (forvar1101 = (1'h0); (forvar1101 < (2'h3)); forvar1101 = (forvar1101 + (1'h1)))
                    begin
                      reg1102 <= ((~|{(8'hb1)}) ?
                          $signed((^~(~&reg1044))) : $signed({reg1002}));
                    end
                  reg1103 <= ($signed($signed((reg1123 * reg1138))) ~^ $signed(reg1131));
                  for (forvar1104 = (1'h0); (forvar1104 < (1'h1)); forvar1104 = (forvar1104 + (1'h1)))
                    begin
                      reg1105 <= $unsigned((forvar1007[(4'h9):(3'h6)] >= {$unsigned(reg1061)}));
                      reg1106 <= (((8'haa) & ((forvar994 <= reg1056) ?
                              (reg1061 ?
                                  reg1001 : forvar1092) : (reg1066 << reg1021))) ?
                          ((reg1053 ?
                              reg1058 : (^reg1144)) <<< $signed(reg1131[(1'h1):(1'h0)])) : (^(reg1097[(4'ha):(3'h5)] ?
                              wire985 : $unsigned(forvar1001))));
                    end
                  for (forvar1107 = (1'h0); (forvar1107 < (1'h1)); forvar1107 = (forvar1107 + (1'h1)))
                    begin
                      reg1108 <= $unsigned(wire981[(1'h1):(1'h0)]);
                      reg1109 <= (^~(|$unsigned((reg1128 ?
                          reg1089 : forvar1058))));
                      reg1110 <= forvar1059;
                      reg1111 <= (!$unsigned($unsigned((reg1113 ~^ reg1003))));
                    end
                end
            end
        end
    end
  assign wire1146 = (~|(reg1023 & {((8'h9f) * reg1059)}));
  assign wire1147 = $signed(($unsigned((reg1016 > reg1083)) ?
                        {reg1065} : (wire986 != (~reg1006))));
  module1148 #() modinst1659 (.y(wire1658), .wire1153(reg1070), .wire1151(reg1038), .wire1149(wire1147), .wire1150(reg1091), .wire1152(reg1097), .clk(clk));
  always
    @(posedge clk) begin
      reg1660 <= reg1040;
      if (((((reg1067 && reg1126) * {reg1037}) ?
          reg1012[(2'h2):(1'h0)] : $signed(reg1087[(3'h6):(2'h3)])) - ((reg1052[(1'h0):(1'h0)] && $unsigned(reg1110)) ~^ ({reg1099} ?
          $unsigned((8'hb6)) : (reg1112 ? reg1058 : (8'ha5))))))
        begin
          if (reg1038)
            begin
              for (forvar1661 = (1'h0); (forvar1661 < (1'h1)); forvar1661 = (forvar1661 + (1'h1)))
                begin
                  if (($unsigned(($unsigned(reg1137) == (reg1119 ?
                          wire1658 : reg1019))) ?
                      reg1036 : ($unsigned($signed(reg1119)) + (|((8'hba) >>> wire982)))))
                    begin
                      reg1662 <= $unsigned((&$unsigned(reg1028)));
                      reg1663 <= reg1119;
                    end
                  else
                    begin
                      reg1662 <= ((~reg1048[(1'h0):(1'h0)]) ?
                          (reg1124[(2'h2):(1'h1)] - (wire1147 <= (reg1076 ?
                              reg1087 : reg1143))) : (&reg1078[(3'h7):(1'h0)]));
                    end
                  if (reg1133[(2'h2):(1'h1)])
                    begin
                      reg1664 <= (($unsigned((reg1037 > reg1005)) ?
                              ((reg1027 >= reg1082) && (~|(8'had))) : $unsigned(reg1122)) ?
                          wire1146 : $signed((^reg1138[(2'h2):(1'h1)])));
                    end
                  else
                    begin
                      reg1664 <= ((reg1042[(4'hc):(2'h3)] ?
                          (~|$signed((8'hb2))) : ($unsigned((8'ha4)) ^~ (reg1106 ?
                              reg1049 : (8'haa)))) ^ reg1143[(4'h8):(3'h4)]);
                      reg1665 <= $signed((reg1085 ?
                          $unsigned($unsigned(reg1009)) : reg989[(1'h1):(1'h0)]));
                    end
                end
            end
          else
            begin
              for (forvar1661 = (1'h0); (forvar1661 < (2'h2)); forvar1661 = (forvar1661 + (1'h1)))
                begin
                  for (forvar1662 = (1'h0); (forvar1662 < (1'h1)); forvar1662 = (forvar1662 + (1'h1)))
                    begin
                      reg1663 <= (($unsigned((reg1117 == reg1132)) ?
                              (|{reg998}) : reg1065) ?
                          $unsigned(($signed(wire983) ^ (reg1016 && reg1025))) : (($signed(forvar1661) ?
                                  reg1076[(3'h4):(1'h0)] : $signed(reg1086)) ?
                              reg1091 : reg1068));
                      reg1664 <= $unsigned(reg1111[(3'h6):(1'h0)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar1661 = (1'h0); (forvar1661 < (1'h0)); forvar1661 = (forvar1661 + (1'h1)))
            begin
              for (forvar1662 = (1'h0); (forvar1662 < (2'h2)); forvar1662 = (forvar1662 + (1'h1)))
                begin
                  if ((-$unsigned($signed(reg1035[(1'h1):(1'h0)]))))
                    begin
                      reg1663 <= (~|$signed(((reg1038 ? (8'hb1) : reg1106) ?
                          $signed((8'ha3)) : (reg1011 < reg1027))));
                    end
                  else
                    begin
                      reg1663 <= reg1127[(3'h4):(2'h2)];
                    end
                end
            end
          reg1664 <= reg1058;
        end
      if ((^~$unsigned(reg1037[(1'h0):(1'h0)])))
        begin
          for (forvar1666 = (1'h0); (forvar1666 < (2'h3)); forvar1666 = (forvar1666 + (1'h1)))
            begin
              if ($signed(reg1109))
                begin
                  for (forvar1667 = (1'h0); (forvar1667 < (1'h0)); forvar1667 = (forvar1667 + (1'h1)))
                    begin
                      reg1668 <= (^~reg1095);
                    end
                  if (reg989[(1'h0):(1'h0)])
                    begin
                      reg1669 <= reg990[(3'h4):(2'h3)];
                      reg1670 <= reg1051[(2'h2):(2'h2)];
                      reg1671 <= $signed(reg1056[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1669 <= reg1038;
                      reg1670 <= (|(($unsigned((8'hb9)) == {reg1671}) ^~ $signed((~^reg1057))));
                      reg1671 <= ($unsigned($unsigned(reg1145)) ?
                          (+$unsigned($signed(reg1127))) : $signed((~(reg1022 ?
                              (8'ha3) : reg1040))));
                    end
                  for (forvar1672 = (1'h0); (forvar1672 < (1'h1)); forvar1672 = (forvar1672 + (1'h1)))
                    begin
                      reg1673 <= {((((8'hab) ?
                              (8'hb6) : reg1057) || {reg1007}) * $unsigned($unsigned(forvar1672)))};
                    end
                end
              else
                begin
                  for (forvar1667 = (1'h0); (forvar1667 < (2'h2)); forvar1667 = (forvar1667 + (1'h1)))
                    begin
                      reg1668 <= (reg1057 ?
                          $signed($signed($unsigned(reg1051))) : $unsigned($unsigned(reg1045[(2'h2):(1'h1)])));
                      reg1669 <= (~^($signed($signed(reg1027)) ?
                          (8'hb3) : reg994[(1'h0):(1'h0)]));
                      reg1670 <= $unsigned((((~^reg1673) ?
                              {reg1091} : $unsigned(reg1011)) ?
                          $unsigned((!reg1673)) : {reg1080}));
                      reg1671 <= {(|reg1111)};
                    end
                end
            end
          for (forvar1674 = (1'h0); (forvar1674 < (2'h2)); forvar1674 = (forvar1674 + (1'h1)))
            begin
              if ((|(({reg1013} ?
                  (reg1135 ?
                      reg1028 : reg1077) : {(8'h9f)}) - reg1090[(3'h4):(1'h1)])))
                begin
                  if ($signed(((&(reg1080 ? (8'ha2) : reg1035)) * reg1128)))
                    begin
                      reg1675 <= (((reg1035 ?
                          $signed(reg1014) : reg1010[(3'h5):(1'h1)]) > (forvar1672[(4'he):(4'h9)] ?
                          $unsigned(reg1082) : (reg1101 ^ reg1145))) * $unsigned(reg1039[(2'h3):(1'h1)]));
                      reg1676 <= $unsigned(($unsigned(reg1670) - {(~|reg1028)}));
                      reg1677 <= ($signed($signed({reg1052})) ?
                          wire981 : (reg1108 ?
                              ($signed(reg1005) ?
                                  {reg1015} : reg1067) : {$unsigned(reg1056)}));
                      reg1678 <= (((-$unsigned(reg1673)) & (8'h9f)) ?
                          (^((reg1663 ? reg1122 : reg1066) ?
                              (~reg1121) : $unsigned(reg1072))) : $unsigned((reg1015 ?
                              reg1677 : (reg1064 >= reg1115))));
                    end
                  else
                    begin
                      reg1675 <= wire987;
                      reg1676 <= forvar1662;
                    end
                end
              else
                begin
                  for (forvar1675 = (1'h0); (forvar1675 < (1'h1)); forvar1675 = (forvar1675 + (1'h1)))
                    begin
                      reg1676 <= (reg1670 ?
                          $unsigned($signed((reg1138 ?
                              reg996 : reg1135))) : (^~(+(reg993 + (8'ha0)))));
                    end
                  for (forvar1677 = (1'h0); (forvar1677 < (2'h3)); forvar1677 = (forvar1677 + (1'h1)))
                    begin
                      reg1678 <= (~$signed(reg994[(2'h2):(2'h2)]));
                      reg1679 <= (~^$signed(reg1039));
                    end
                  if ($signed($unsigned(reg1007[(4'h8):(2'h3)])))
                    begin
                      reg1680 <= $unsigned(((|{reg1086}) ?
                          (|{reg995}) : ($unsigned(reg1111) ?
                              ((8'hab) >= reg1110) : (reg1011 ?
                                  (8'hab) : (8'hb9)))));
                    end
                  else
                    begin
                      reg1680 <= (reg1126[(1'h0):(1'h0)] ?
                          ({{reg1017}} >> $unsigned(reg1665)) : {$signed((^forvar1666))});
                    end
                  for (forvar1681 = (1'h0); (forvar1681 < (2'h2)); forvar1681 = (forvar1681 + (1'h1)))
                    begin
                      reg1682 <= reg1094;
                      reg1683 <= reg1026[(2'h3):(1'h1)];
                      reg1684 <= ((!(|(-reg1134))) < (reg1017[(2'h3):(1'h0)] ?
                          (-(~&reg1124)) : (~|(reg1090 << reg1066))));
                      reg1685 <= (+reg1101[(2'h3):(2'h2)]);
                    end
                end
            end
        end
      else
        begin
          reg1666 <= $signed(reg999);
        end
      for (forvar1686 = (1'h0); (forvar1686 < (2'h2)); forvar1686 = (forvar1686 + (1'h1)))
        begin
          for (forvar1687 = (1'h0); (forvar1687 < (2'h3)); forvar1687 = (forvar1687 + (1'h1)))
            begin
              for (forvar1688 = (1'h0); (forvar1688 < (1'h1)); forvar1688 = (forvar1688 + (1'h1)))
                begin
                  for (forvar1689 = (1'h0); (forvar1689 < (1'h1)); forvar1689 = (forvar1689 + (1'h1)))
                    begin
                      reg1690 <= (^reg1058);
                      reg1691 <= $signed((($unsigned(reg1670) ?
                          $signed(reg1034) : (&reg1116)) << $unsigned((8'ha0))));
                      reg1692 <= $unsigned({reg1118[(2'h3):(2'h2)]});
                      reg1693 <= reg1013[(1'h1):(1'h0)];
                    end
                  for (forvar1694 = (1'h0); (forvar1694 < (2'h3)); forvar1694 = (forvar1694 + (1'h1)))
                    begin
                      reg1695 <= ((~$unsigned($signed((8'hb9)))) ?
                          ((reg1075[(3'h7):(2'h3)] ?
                              (!reg1144) : $signed(reg1097)) > $signed((reg1119 ?
                              reg1039 : reg1142))) : (($unsigned(reg1673) - ((8'ha1) <<< reg1144)) <<< $signed($signed(reg1104))));
                    end
                end
              for (forvar1696 = (1'h0); (forvar1696 < (1'h0)); forvar1696 = (forvar1696 + (1'h1)))
                begin
                  reg1697 <= reg1134;
                  for (forvar1698 = (1'h0); (forvar1698 < (2'h3)); forvar1698 = (forvar1698 + (1'h1)))
                    begin
                      reg1699 <= (^~reg1070[(2'h2):(1'h1)]);
                      reg1700 <= (^wire982[(4'h8):(3'h5)]);
                      reg1701 <= (reg1103[(2'h2):(1'h0)] ?
                          reg1118 : (reg1042 == $unsigned((~(8'h9f)))));
                    end
                  reg1702 <= reg1130[(4'h8):(3'h6)];
                  reg1703 <= (^reg1690[(4'h8):(2'h3)]);
                end
            end
          reg1704 <= reg1108[(2'h2):(2'h2)];
        end
    end
  assign wire1705 = {(|{reg1118[(1'h0):(1'h0)]})};
  always
    @(posedge clk) begin
      if ({$unsigned(((|reg1056) < $signed(wire986)))})
        begin
          reg1706 <= reg1039;
          for (forvar1707 = (1'h0); (forvar1707 < (1'h1)); forvar1707 = (forvar1707 + (1'h1)))
            begin
              for (forvar1708 = (1'h0); (forvar1708 < (2'h3)); forvar1708 = (forvar1708 + (1'h1)))
                begin
                  reg1709 <= reg995;
                  if ($unsigned($signed((8'hb4))))
                    begin
                      reg1710 <= $signed(reg1675[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg1710 <= $signed((8'haf));
                      reg1711 <= (~^reg1125);
                    end
                  if ((reg1080[(1'h0):(1'h0)] ^ forvar1708))
                    begin
                      reg1712 <= (8'ha5);
                      reg1713 <= reg1003;
                    end
                  else
                    begin
                      reg1712 <= {((+$signed((8'h9c))) ?
                              $signed({reg1095}) : $unsigned(wire982))};
                    end
                  reg1714 <= reg1014[(1'h1):(1'h0)];
                end
            end
          if ($unsigned({reg1038}))
            begin
              if ((-reg1702))
                begin
                  for (forvar1715 = (1'h0); (forvar1715 < (2'h3)); forvar1715 = (forvar1715 + (1'h1)))
                    begin
                      reg1716 <= ($unsigned(reg1142) && (reg1025[(4'hd):(1'h1)] ?
                          reg1018[(3'h4):(3'h4)] : reg1027[(4'hd):(4'hd)]));
                      reg1717 <= $signed(wire982[(3'h6):(2'h2)]);
                      reg1718 <= ($signed($unsigned(reg1007)) ?
                          reg1057[(3'h5):(2'h2)] : (((~reg1006) ?
                                  (+(8'h9c)) : reg1679[(3'h4):(1'h1)]) ?
                              $unsigned(reg1098[(1'h1):(1'h1)]) : reg1144[(2'h3):(1'h1)]));
                      reg1719 <= ((!wire1146) != $unsigned((~|(8'hb9))));
                    end
                end
              else
                begin
                  reg1715 <= $unsigned((reg1666 ?
                      (~^(~|reg1027)) : (reg1051 ?
                          $unsigned(reg1123) : reg1704)));
                  if ($signed(reg1666))
                    begin
                      reg1716 <= $signed(reg989[(1'h0):(1'h0)]);
                      reg1717 <= (((-reg1714) <<< reg1098[(1'h1):(1'h0)]) ~^ ({(|reg1715)} ?
                          {((8'ha5) ?
                                  reg1037 : wire984)} : $unsigned($signed(reg1059))));
                    end
                  else
                    begin
                      reg1716 <= (reg1036 ?
                          ($signed($signed(reg1142)) - reg1091) : $unsigned($unsigned(reg1693[(1'h1):(1'h0)])));
                    end
                  for (forvar1718 = (1'h0); (forvar1718 < (2'h3)); forvar1718 = (forvar1718 + (1'h1)))
                    begin
                      reg1719 <= (8'h9f);
                      reg1720 <= reg1063;
                      reg1721 <= $signed($signed($signed((&reg1101))));
                      reg1722 <= (reg1135[(4'ha):(3'h4)] ?
                          (reg1666 << (&(reg1036 == reg1134))) : reg1714[(2'h3):(1'h0)]);
                    end
                  for (forvar1723 = (1'h0); (forvar1723 < (2'h3)); forvar1723 = (forvar1723 + (1'h1)))
                    begin
                      reg1724 <= (reg990[(3'h6):(1'h1)] & reg1090);
                      reg1725 <= ($signed(reg1717) ?
                          ((reg1677 ?
                                  $signed(reg1045) : ((8'h9e) ?
                                      reg990 : (8'ha5))) ?
                              forvar1707 : ((reg1039 < reg1005) ?
                                  {reg1719} : (reg989 > reg1056))) : $unsigned((8'ha4)));
                    end
                end
              if ((reg1041[(1'h0):(1'h0)] ? (!$signed((-reg1096))) : wire1658))
                begin
                  for (forvar1726 = (1'h0); (forvar1726 < (1'h1)); forvar1726 = (forvar1726 + (1'h1)))
                    begin
                      reg1727 <= forvar1718[(4'ha):(3'h7)];
                      reg1728 <= ($signed({$signed(reg1144)}) ?
                          reg1013 : {(~^((8'ha8) ? reg1015 : reg1135))});
                      reg1729 <= (^($unsigned(reg1670) <<< reg1030));
                      reg1730 <= reg1129;
                    end
                  for (forvar1731 = (1'h0); (forvar1731 < (1'h1)); forvar1731 = (forvar1731 + (1'h1)))
                    begin
                      reg1732 <= reg1126;
                      reg1733 <= wire1146[(2'h2):(1'h1)];
                      reg1734 <= $unsigned((^(8'hb4)));
                      reg1735 <= reg1096[(3'h4):(2'h3)];
                    end
                  reg1736 <= $signed(reg1676[(3'h4):(3'h4)]);
                  for (forvar1737 = (1'h0); (forvar1737 < (1'h1)); forvar1737 = (forvar1737 + (1'h1)))
                    begin
                      reg1738 <= ($signed($signed($signed(reg1003))) ?
                          reg1068[(3'h4):(3'h4)] : wire1147);
                    end
                end
              else
                begin
                  if ((&$unsigned((((8'hba) ?
                      reg1077 : forvar1731) < reg1009))))
                    begin
                      reg1726 <= (|$signed($unsigned($signed((8'haa)))));
                    end
                  else
                    begin
                      reg1726 <= reg1717;
                      reg1727 <= $signed($signed(reg1041[(2'h2):(1'h1)]));
                      reg1728 <= $unsigned(reg1703);
                      reg1729 <= (!$signed((reg992[(1'h1):(1'h1)] != (reg1113 ?
                          reg994 : reg990))));
                    end
                  reg1730 <= (((~|((8'hb0) ? reg1065 : reg1016)) ?
                      ((~reg1704) ?
                          (reg1016 | reg1036) : reg1700) : ({reg1716} <= {(8'ha4)})) < $unsigned($unsigned((reg1668 == reg1018))));
                  if (reg1697)
                    begin
                      reg1731 <= ((^~((^~reg1673) + reg1077[(2'h3):(1'h1)])) > {($unsigned((8'ha2)) < {reg1662})});
                      reg1732 <= $signed((~reg1735[(4'hc):(3'h4)]));
                      reg1733 <= (reg1715 ?
                          (^~$unsigned(reg1126[(2'h2):(1'h1)])) : ($unsigned((reg1712 ?
                              reg1082 : reg994)) >> $unsigned($signed((8'h9f)))));
                    end
                  else
                    begin
                      reg1731 <= (+$signed(reg1666));
                      reg1732 <= reg1014[(3'h4):(2'h3)];
                      reg1733 <= ((reg1138 >= reg1110) ?
                          reg1014[(2'h2):(1'h1)] : {{{reg1129}}});
                      reg1734 <= $unsigned({$signed(reg997[(1'h1):(1'h0)])});
                    end
                  if (reg1065[(3'h5):(2'h2)])
                    begin
                      reg1735 <= $unsigned({(^~$signed(reg1690))});
                    end
                  else
                    begin
                      reg1735 <= (reg1112[(4'h9):(4'h8)] == (8'ha0));
                    end
                end
              for (forvar1739 = (1'h0); (forvar1739 < (1'h0)); forvar1739 = (forvar1739 + (1'h1)))
                begin
                  reg1740 <= reg1059[(2'h2):(2'h2)];
                  if ((^reg1035))
                    begin
                      reg1741 <= (^~reg1030);
                    end
                  else
                    begin
                      reg1741 <= $signed((($signed(reg1127) + (wire983 - reg996)) ?
                          $signed((reg1060 ?
                              reg1733 : reg1729)) : ((~|forvar1739) ?
                              (reg1740 && reg1725) : $signed(reg1711))));
                      reg1742 <= (8'hac);
                      reg1743 <= (reg1062[(1'h1):(1'h1)] >= ({(reg1740 ?
                              reg1664 : reg1015)} + reg1129[(4'ha):(2'h3)]));
                    end
                  if (($signed($signed($signed((8'h9d)))) && $signed((reg1137[(3'h5):(3'h5)] > {reg1108}))))
                    begin
                      reg1744 <= $signed(({reg1074} * (^(reg1051 ?
                          (8'ha6) : reg1081))));
                    end
                  else
                    begin
                      reg1744 <= $signed($unsigned((~&$unsigned(reg1732))));
                      reg1745 <= reg1732[(3'h6):(1'h0)];
                    end
                end
              for (forvar1746 = (1'h0); (forvar1746 < (1'h1)); forvar1746 = (forvar1746 + (1'h1)))
                begin
                  for (forvar1747 = (1'h0); (forvar1747 < (1'h1)); forvar1747 = (forvar1747 + (1'h1)))
                    begin
                      reg1748 <= forvar1707[(2'h2):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar1715 = (1'h0); (forvar1715 < (1'h0)); forvar1715 = (forvar1715 + (1'h1)))
                begin
                  for (forvar1716 = (1'h0); (forvar1716 < (2'h3)); forvar1716 = (forvar1716 + (1'h1)))
                    begin
                      reg1717 <= $unsigned((!((reg1052 ?
                          wire1658 : reg995) | (reg1013 ? reg1041 : reg1045))));
                      reg1718 <= reg1058[(4'h9):(4'h8)];
                      reg1719 <= ({((reg1025 ?
                                  reg1139 : reg1097) ^~ reg1733[(2'h3):(2'h3)])} ?
                          ({reg1736} ?
                              ((8'hb4) + {(8'haa)}) : $signed((reg1001 ^ wire981))) : $unsigned(($signed(forvar1708) && {forvar1718})));
                      reg1720 <= $signed(reg1074[(1'h0):(1'h0)]);
                    end
                  for (forvar1721 = (1'h0); (forvar1721 < (2'h3)); forvar1721 = (forvar1721 + (1'h1)))
                    begin
                      reg1722 <= reg1103[(3'h5):(1'h1)];
                      reg1723 <= (reg1103[(2'h3):(2'h2)] || $signed((~|{wire1658})));
                    end
                  reg1724 <= (reg1680[(1'h0):(1'h0)] ?
                      $signed({$unsigned(reg1714)}) : (!reg1712[(4'h9):(4'h8)]));
                  reg1725 <= ({($signed(reg1132) ?
                          reg1137 : (reg1692 <= forvar1731))} ^~ $signed($signed({forvar1715})));
                end
              for (forvar1726 = (1'h0); (forvar1726 < (1'h1)); forvar1726 = (forvar1726 + (1'h1)))
                begin
                  reg1727 <= $unsigned(reg1077[(2'h3):(1'h1)]);
                  if ($signed((8'ha2)))
                    begin
                      reg1728 <= (reg1003[(3'h4):(1'h0)] << reg994[(1'h1):(1'h0)]);
                      reg1729 <= reg1083;
                      reg1730 <= ($unsigned((((8'hb5) ?
                              (8'haf) : reg1077) * reg1710[(1'h1):(1'h1)])) ?
                          $signed(forvar1731[(3'h5):(3'h4)]) : (reg1665[(4'ha):(2'h2)] & ((~&reg1735) ?
                              reg1703 : reg1022)));
                    end
                  else
                    begin
                      reg1728 <= ((reg1006[(4'h8):(4'h8)] ~^ (&{(8'hb9)})) ?
                          (reg1700[(1'h1):(1'h1)] ?
                              (-(~|reg1666)) : ((reg1015 ?
                                  reg1102 : reg1713) * (+reg1123))) : (~|reg1742[(1'h1):(1'h1)]));
                      reg1729 <= $unsigned(reg1040);
                      reg1730 <= (~(8'haa));
                      reg1731 <= $signed($unsigned($unsigned(reg1025)));
                    end
                  reg1732 <= ((~|(reg1113 ?
                          (reg1726 >= reg1129) : ((8'hb9) * reg1038))) ?
                      reg1022[(1'h0):(1'h0)] : {reg1103});
                  for (forvar1733 = (1'h0); (forvar1733 < (1'h0)); forvar1733 = (forvar1733 + (1'h1)))
                    begin
                      reg1734 <= $signed(($unsigned($unsigned((8'h9f))) | $unsigned($unsigned(reg1108))));
                      reg1735 <= $signed((8'haf));
                    end
                end
              for (forvar1736 = (1'h0); (forvar1736 < (1'h1)); forvar1736 = (forvar1736 + (1'h1)))
                begin
                  reg1737 <= {reg1663[(1'h0):(1'h0)]};
                  for (forvar1738 = (1'h0); (forvar1738 < (1'h1)); forvar1738 = (forvar1738 + (1'h1)))
                    begin
                      reg1739 <= forvar1737[(4'h9):(3'h7)];
                      reg1740 <= $signed($unsigned(($signed(reg1115) ?
                          (reg1052 ? reg1082 : wire985) : $signed((8'ha5)))));
                      reg1741 <= $signed($signed((8'hb0)));
                    end
                  for (forvar1742 = (1'h0); (forvar1742 < (2'h2)); forvar1742 = (forvar1742 + (1'h1)))
                    begin
                      reg1743 <= $unsigned($signed((8'hb0)));
                      reg1744 <= $unsigned((forvar1733[(4'hc):(4'hc)] || reg1068[(2'h2):(2'h2)]));
                      reg1745 <= reg1675[(3'h6):(1'h0)];
                    end
                  for (forvar1746 = (1'h0); (forvar1746 < (1'h1)); forvar1746 = (forvar1746 + (1'h1)))
                    begin
                      reg1747 <= {{reg1670[(4'h9):(4'h9)]}};
                      reg1748 <= $unsigned(((~|((8'hb3) | reg1722)) || {(reg1715 ?
                              reg1102 : reg1044)}));
                      reg1749 <= (8'hb4);
                      reg1750 <= reg1700;
                    end
                end
              for (forvar1751 = (1'h0); (forvar1751 < (1'h1)); forvar1751 = (forvar1751 + (1'h1)))
                begin
                  for (forvar1752 = (1'h0); (forvar1752 < (1'h0)); forvar1752 = (forvar1752 + (1'h1)))
                    begin
                      reg1753 <= ($unsigned(({wire1147} + (reg1117 ?
                          (8'hb7) : reg1091))) << reg1058[(4'hb):(1'h1)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar1706 = (1'h0); (forvar1706 < (2'h2)); forvar1706 = (forvar1706 + (1'h1)))
            begin
              for (forvar1707 = (1'h0); (forvar1707 < (1'h1)); forvar1707 = (forvar1707 + (1'h1)))
                begin
                  if ({$unsigned($signed($unsigned(reg1706)))})
                    begin
                      reg1708 <= ((8'ha7) ?
                          reg1037[(2'h2):(1'h1)] : (((-reg1144) | (^reg1693)) ?
                              reg1058[(1'h0):(1'h0)] : reg1012));
                    end
                  else
                    begin
                      reg1708 <= (~({(reg1715 <= (8'h9c))} ?
                          (~|(reg1070 ?
                              (8'ha9) : wire987)) : $signed({reg1052})));
                      reg1709 <= ({$unsigned((reg999 || reg1006))} + $signed(reg1716));
                      reg1710 <= ((($signed(forvar1706) || reg1662) || reg1749) != ((8'haa) ?
                          $unsigned(forvar1726[(4'h8):(4'h8)]) : reg1115));
                      reg1711 <= (($signed($signed(reg1099)) ?
                          $signed($unsigned(reg1131)) : reg1713) ^ (&(~$signed(reg1101))));
                    end
                  for (forvar1712 = (1'h0); (forvar1712 < (1'h1)); forvar1712 = (forvar1712 + (1'h1)))
                    begin
                      reg1713 <= $unsigned(reg1680[(2'h2):(1'h0)]);
                      reg1714 <= ((forvar1742[(3'h5):(1'h1)] << (reg1095[(1'h0):(1'h0)] < {reg1750})) ?
                          {reg1089} : reg1016);
                    end
                end
              for (forvar1715 = (1'h0); (forvar1715 < (2'h3)); forvar1715 = (forvar1715 + (1'h1)))
                begin
                  for (forvar1716 = (1'h0); (forvar1716 < (2'h3)); forvar1716 = (forvar1716 + (1'h1)))
                    begin
                      reg1717 <= ((($signed((8'haa)) ?
                          $unsigned(reg1131) : ((8'haf) & reg1025)) ^~ reg1050[(3'h5):(3'h5)]) | $unsigned($unsigned($unsigned(reg1126))));
                      reg1718 <= wire987[(2'h2):(2'h2)];
                    end
                  if (reg1003)
                    begin
                      reg1719 <= reg1040;
                      reg1720 <= ((!({reg1747} | reg1039[(1'h1):(1'h1)])) >>> (^(~|reg1736[(2'h2):(1'h1)])));
                    end
                  else
                    begin
                      reg1719 <= $signed((^~reg1066[(2'h2):(1'h0)]));
                      reg1720 <= (reg1089[(3'h4):(2'h2)] * (({reg1083} <= (reg1714 <<< reg1117)) ?
                          {(~|reg1141)} : reg1036[(1'h1):(1'h0)]));
                      reg1721 <= $signed($unsigned({reg1017[(3'h4):(1'h0)]}));
                      reg1722 <= reg1130;
                    end
                  for (forvar1723 = (1'h0); (forvar1723 < (2'h3)); forvar1723 = (forvar1723 + (1'h1)))
                    begin
                      reg1724 <= reg1695[(3'h4):(1'h0)];
                      reg1725 <= reg1729[(4'he):(2'h3)];
                      reg1726 <= $unsigned(reg1121[(4'ha):(1'h1)]);
                    end
                end
              reg1727 <= (~((!(reg1679 ?
                  reg1738 : reg1727)) | $signed($signed(reg1065))));
              for (forvar1728 = (1'h0); (forvar1728 < (1'h0)); forvar1728 = (forvar1728 + (1'h1)))
                begin
                  for (forvar1729 = (1'h0); (forvar1729 < (1'h0)); forvar1729 = (forvar1729 + (1'h1)))
                    begin
                      reg1730 <= (reg1115[(3'h4):(3'h4)] ?
                          ((~^(~reg1137)) ?
                              reg1044[(2'h2):(2'h2)] : ((reg1743 ?
                                  forvar1729 : reg1712) >>> $unsigned((8'ha2)))) : reg1726[(3'h7):(3'h7)]);
                    end
                  for (forvar1731 = (1'h0); (forvar1731 < (2'h2)); forvar1731 = (forvar1731 + (1'h1)))
                    begin
                      reg1732 <= {$unsigned(reg1108)};
                      reg1733 <= $unsigned((reg1057[(3'h6):(3'h6)] ?
                          reg1714[(1'h1):(1'h1)] : (~&reg1727[(4'ha):(3'h4)])));
                    end
                  for (forvar1734 = (1'h0); (forvar1734 < (1'h0)); forvar1734 = (forvar1734 + (1'h1)))
                    begin
                      reg1735 <= forvar1712[(1'h0):(1'h0)];
                      reg1736 <= $unsigned($signed(($signed(forvar1707) >>> forvar1715)));
                      reg1737 <= wire987;
                      reg1738 <= (|forvar1734);
                    end
                  if ($signed($unsigned(($signed(reg1111) ?
                      ((8'ha0) ? reg1064 : reg1023) : (8'hb3)))))
                    begin
                      reg1739 <= ({reg1054[(2'h3):(2'h3)]} ?
                          (~(-$unsigned(reg1675))) : (^~$unsigned($signed(reg1747))));
                    end
                  else
                    begin
                      reg1739 <= reg1082[(1'h0):(1'h0)];
                      reg1740 <= $unsigned((&((+reg1107) ?
                          (&reg993) : ((8'hb5) > reg1050))));
                    end
                end
            end
        end
      if ($signed((&(!(reg1731 && reg1118)))))
        begin
          reg1754 <= (reg1063 ?
              $unsigned((~|(forvar1739 >>> (8'h9e)))) : $unsigned($signed($unsigned(reg990))));
          reg1755 <= {reg1715[(1'h0):(1'h0)]};
          for (forvar1756 = (1'h0); (forvar1756 < (1'h1)); forvar1756 = (forvar1756 + (1'h1)))
            begin
              for (forvar1757 = (1'h0); (forvar1757 < (1'h0)); forvar1757 = (forvar1757 + (1'h1)))
                begin
                  for (forvar1758 = (1'h0); (forvar1758 < (1'h1)); forvar1758 = (forvar1758 + (1'h1)))
                    begin
                      reg1759 <= $unsigned(reg1042);
                      reg1760 <= ((reg1044[(1'h0):(1'h0)] * ($signed((8'hb4)) * $unsigned((8'ha6)))) >= reg1006[(2'h2):(1'h0)]);
                      reg1761 <= $unsigned(((~|$unsigned(reg1679)) ?
                          reg1119[(1'h0):(1'h0)] : (reg1016[(3'h4):(3'h4)] ?
                              reg1009 : $unsigned(reg1717))));
                    end
                  if ((^($unsigned(reg1021) ^ ({reg1011} | reg1724))))
                    begin
                      reg1762 <= reg1028[(1'h0):(1'h0)];
                      reg1763 <= (^reg1062[(3'h5):(3'h5)]);
                    end
                  else
                    begin
                      reg1762 <= (+($signed((reg1690 ? reg1706 : reg1734)) ?
                          ({reg1743} ? forvar1737 : forvar1758) : reg1119));
                      reg1763 <= (~^reg1103);
                    end
                  if ((8'hb6))
                    begin
                      reg1764 <= reg1058;
                      reg1765 <= $unsigned(((reg1712 ^~ (+reg1700)) & ($signed(reg1085) >= (~^reg1025))));
                    end
                  else
                    begin
                      reg1764 <= $signed((8'ha3));
                      reg1765 <= reg1042[(4'hf):(3'h6)];
                      reg1766 <= reg1019[(2'h2):(2'h2)];
                      reg1767 <= reg1124[(2'h2):(1'h1)];
                    end
                  if (reg1015[(4'hf):(4'hc)])
                    begin
                      reg1768 <= (~^($signed(reg1051) ?
                          reg1710 : ($unsigned(reg1119) ?
                              $signed(reg1713) : (+reg1141))));
                      reg1769 <= $signed(reg1028[(2'h2):(1'h1)]);
                      reg1770 <= reg1002;
                      reg1771 <= (((~&$signed(reg1670)) >>> (reg1683 ^ reg1709)) ?
                          $signed($signed((reg1089 - reg1028))) : {$signed({(8'hae)})});
                    end
                  else
                    begin
                      reg1768 <= ((~&$unsigned((reg1692 | reg1074))) && reg1738[(2'h2):(2'h2)]);
                      reg1769 <= ((~|((!reg1670) + reg1750[(3'h6):(3'h4)])) || $unsigned({(~^reg1001)}));
                      reg1770 <= (|{($signed(reg1693) ?
                              forvar1751 : reg1731[(4'hf):(3'h6)])});
                      reg1771 <= (^~($unsigned(forvar1707[(1'h0):(1'h0)]) ?
                          (reg1680[(3'h4):(3'h4)] ?
                              (&reg1091) : $unsigned(reg1006)) : reg1679));
                    end
                end
              for (forvar1772 = (1'h0); (forvar1772 < (2'h3)); forvar1772 = (forvar1772 + (1'h1)))
                begin
                  if (reg1741[(3'h4):(2'h2)])
                    begin
                      reg1773 <= reg1076[(3'h6):(3'h6)];
                      reg1774 <= (~|($unsigned($unsigned((8'ha0))) ?
                          $unsigned(reg1086[(4'h9):(1'h0)]) : forvar1739[(4'hb):(4'h9)]));
                    end
                  else
                    begin
                      reg1773 <= forvar1706[(2'h3):(2'h3)];
                      reg1774 <= wire987[(3'h6):(1'h1)];
                    end
                end
              for (forvar1775 = (1'h0); (forvar1775 < (1'h1)); forvar1775 = (forvar1775 + (1'h1)))
                begin
                  for (forvar1776 = (1'h0); (forvar1776 < (1'h1)); forvar1776 = (forvar1776 + (1'h1)))
                    begin
                      reg1777 <= ($unsigned($unsigned((!(8'h9d)))) ?
                          reg1724 : (~&$signed((reg1134 || (8'ha0)))));
                      reg1778 <= reg1122;
                      reg1779 <= {((reg999 != $unsigned((8'ha9))) ^ (((8'hb1) ?
                                  wire981 : reg1115) ?
                              (reg1769 ?
                                  reg1037 : reg1683) : reg1137[(3'h5):(3'h5)]))};
                      reg1780 <= (forvar1721[(1'h1):(1'h1)] && $unsigned(forvar1718[(3'h6):(1'h1)]));
                    end
                  if ($signed((reg1748[(4'h9):(1'h0)] ?
                      $unsigned((reg1143 * forvar1729)) : ((reg1139 ?
                              forvar1739 : (8'hb5)) ?
                          reg1770[(3'h7):(3'h7)] : reg1145))))
                    begin
                      reg1781 <= $signed(((-(reg1081 <<< (8'hba))) == (^~(reg1142 ?
                          reg1117 : reg1110))));
                      reg1782 <= ((reg1057[(1'h1):(1'h0)] ?
                          {(reg999 ?
                                  reg1111 : reg1058)} : (8'ha2)) ^~ (~^(forvar1706 ?
                          reg1699[(4'hd):(1'h0)] : reg1668)));
                      reg1783 <= $signed(forvar1738[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg1781 <= $unsigned((reg1697[(3'h4):(2'h3)] ?
                          (reg1125 ?
                              ((8'hb2) | reg1009) : {forvar1772}) : $unsigned($signed(reg1677))));
                      reg1782 <= reg1115;
                      reg1783 <= reg1678;
                      reg1784 <= $unsigned((!{(reg991 ? reg1728 : reg1002)}));
                    end
                  reg1785 <= (reg1026[(1'h1):(1'h1)] ~^ (~|reg1711));
                end
              reg1786 <= (^$unsigned((8'hb0)));
            end
        end
      else
        begin
          for (forvar1754 = (1'h0); (forvar1754 < (2'h2)); forvar1754 = (forvar1754 + (1'h1)))
            begin
              if (({(-reg1750[(3'h4):(2'h3)])} >= reg1678))
                begin
                  for (forvar1755 = (1'h0); (forvar1755 < (2'h3)); forvar1755 = (forvar1755 + (1'h1)))
                    begin
                      reg1756 <= (~^$unsigned(reg1764[(3'h5):(2'h2)]));
                      reg1757 <= (($signed((reg1036 ^ reg1119)) >>> reg1075) | $unsigned((reg1738[(4'hd):(4'ha)] + (8'hb6))));
                      reg1758 <= reg1110[(2'h2):(1'h1)];
                      reg1759 <= reg1709[(4'h8):(3'h5)];
                    end
                  for (forvar1760 = (1'h0); (forvar1760 < (1'h1)); forvar1760 = (forvar1760 + (1'h1)))
                    begin
                      reg1761 <= (reg1077 ?
                          forvar1757[(2'h3):(1'h1)] : ((~&(forvar1707 ?
                                  forvar1757 : reg1113)) ?
                              reg1726[(3'h7):(3'h4)] : $signed((reg1718 <= (8'hae)))));
                      reg1762 <= (8'ha2);
                    end
                  for (forvar1763 = (1'h0); (forvar1763 < (1'h1)); forvar1763 = (forvar1763 + (1'h1)))
                    begin
                      reg1764 <= {$unsigned($unsigned($unsigned(reg1093)))};
                      reg1765 <= $signed(reg1677);
                      reg1766 <= $signed($unsigned($signed(reg1008)));
                      reg1767 <= (&$unsigned($signed(wire986)));
                    end
                end
              else
                begin
                  for (forvar1755 = (1'h0); (forvar1755 < (1'h0)); forvar1755 = (forvar1755 + (1'h1)))
                    begin
                      reg1756 <= {$unsigned($signed($signed(reg1760)))};
                      reg1757 <= $signed({(((8'hab) ? reg1717 : reg1035) ?
                              (reg1118 ? reg1663 : (8'hba)) : (reg1734 ?
                                  reg1713 : reg1716))});
                    end
                  reg1758 <= ((((reg1663 ? reg1142 : reg1676) ?
                          reg1077[(2'h2):(1'h0)] : {reg1145}) ?
                      (reg1721[(2'h2):(1'h0)] ?
                          reg1075 : ((8'had) ?
                              reg1018 : reg1086)) : reg1088) ^~ $unsigned($unsigned((-reg1098))));
                end
              for (forvar1768 = (1'h0); (forvar1768 < (2'h3)); forvar1768 = (forvar1768 + (1'h1)))
                begin
                  for (forvar1769 = (1'h0); (forvar1769 < (1'h0)); forvar1769 = (forvar1769 + (1'h1)))
                    begin
                      reg1770 <= ((|((~(8'hb3)) <<< (reg1106 ?
                              reg1060 : reg1756))) ?
                          reg1101 : (reg1747 | $signed($signed((8'hba)))));
                      reg1771 <= (reg1763[(2'h3):(2'h2)] ?
                          (~^reg1098) : $unsigned((~|(~^forvar1731))));
                      reg1772 <= (^~$signed(reg1035));
                    end
                  for (forvar1773 = (1'h0); (forvar1773 < (2'h3)); forvar1773 = (forvar1773 + (1'h1)))
                    begin
                      reg1774 <= reg1039;
                      reg1775 <= reg1093[(2'h3):(2'h2)];
                    end
                end
              for (forvar1776 = (1'h0); (forvar1776 < (2'h2)); forvar1776 = (forvar1776 + (1'h1)))
                begin
                  if ((8'haa))
                    begin
                      reg1777 <= reg1064[(3'h6):(3'h5)];
                      reg1778 <= forvar1754;
                      reg1779 <= (^~(($unsigned((8'h9d)) < (8'ha8)) & reg1670[(4'he):(1'h1)]));
                    end
                  else
                    begin
                      reg1777 <= $unsigned({($unsigned(reg1692) ?
                              $unsigned((8'hb1)) : (reg1098 == reg1692))});
                      reg1778 <= $unsigned((&($unsigned(reg1782) ~^ (reg1774 ~^ forvar1715))));
                      reg1779 <= (({$signed((8'ha7))} ?
                              reg1721 : $unsigned(reg1775)) ?
                          ($signed(reg1058) ?
                              reg1669 : reg1018) : (($signed(reg1724) & forvar1755[(4'hc):(3'h6)]) * $signed(reg1065[(3'h5):(2'h2)])));
                      reg1780 <= $signed((8'hb9));
                    end
                end
            end
        end
      if ($signed(($signed(reg1722) ?
          (reg1771 == (forvar1708 ?
              reg1693 : reg1750)) : $signed($unsigned(reg1052)))))
        begin
          for (forvar1787 = (1'h0); (forvar1787 < (1'h1)); forvar1787 = (forvar1787 + (1'h1)))
            begin
              if (((($unsigned(reg1786) ?
                  {forvar1729} : (reg1671 && reg1671)) == $unsigned({forvar1746})) >= $unsigned(($signed(reg1033) ?
                  $unsigned(reg1075) : (reg1748 != reg1673)))))
                begin
                  reg1788 <= $signed(reg1034[(4'hb):(1'h0)]);
                  for (forvar1789 = (1'h0); (forvar1789 < (1'h0)); forvar1789 = (forvar1789 + (1'h1)))
                    begin
                      reg1790 <= $signed(((8'h9e) ?
                          (forvar1756[(4'hd):(4'h8)] ^ reg1700) : reg1059));
                      reg1791 <= reg1010[(1'h0):(1'h0)];
                      reg1792 <= reg1762[(3'h4):(3'h4)];
                      reg1793 <= reg1037[(2'h2):(1'h1)];
                    end
                  for (forvar1794 = (1'h0); (forvar1794 < (2'h2)); forvar1794 = (forvar1794 + (1'h1)))
                    begin
                      reg1795 <= reg1783[(2'h2):(1'h1)];
                      reg1796 <= reg1763[(2'h3):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar1788 = (1'h0); (forvar1788 < (2'h3)); forvar1788 = (forvar1788 + (1'h1)))
                    begin
                      reg1789 <= {$unsigned(reg1679)};
                      reg1790 <= forvar1723;
                    end
                end
              reg1797 <= reg1774;
            end
        end
      else
        begin
          for (forvar1787 = (1'h0); (forvar1787 < (1'h1)); forvar1787 = (forvar1787 + (1'h1)))
            begin
              for (forvar1788 = (1'h0); (forvar1788 < (2'h2)); forvar1788 = (forvar1788 + (1'h1)))
                begin
                  reg1789 <= (-reg1779[(3'h7):(3'h7)]);
                  if ((-((reg1036[(3'h6):(1'h1)] ?
                      reg1027 : reg1779[(1'h1):(1'h1)]) - forvar1789[(3'h4):(3'h4)])))
                    begin
                      reg1790 <= ((&(|(reg1766 ?
                          reg1078 : reg1102))) ^~ (reg1011[(3'h6):(2'h3)] ?
                          ({reg1018} && $unsigned(forvar1794)) : reg1791[(4'h8):(3'h6)]));
                      reg1791 <= {((~$unsigned(reg1684)) | {reg1753})};
                      reg1792 <= $signed($unsigned(reg1129[(4'h8):(4'h8)]));
                      reg1793 <= wire984[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg1790 <= reg1095[(3'h5):(1'h0)];
                      reg1791 <= $unsigned((forvar1707[(3'h4):(2'h3)] & (&(forvar1768 ~^ forvar1752))));
                      reg1792 <= reg1087;
                    end
                  if ($unsigned({({reg1030} ?
                          reg991[(3'h6):(1'h1)] : forvar1787)}))
                    begin
                      reg1794 <= (reg1093 ^~ ($unsigned(reg1769[(1'h0):(1'h0)]) <= ($unsigned(reg1119) ^~ $signed(wire986))));
                      reg1795 <= $signed($signed({reg1761}));
                      reg1796 <= (reg1118 ^ ({$unsigned((8'h9f))} ?
                          ($signed(reg1131) ^~ $unsigned(forvar1754)) : $signed(((8'haf) || reg1076))));
                      reg1797 <= $signed($unsigned(reg1730[(4'h8):(1'h0)]));
                    end
                  else
                    begin
                      reg1794 <= (~&$unsigned((8'ha7)));
                      reg1795 <= $signed((($signed(reg1775) && (&reg1756)) > reg1722[(4'ha):(4'ha)]));
                      reg1796 <= $signed($signed(reg1745));
                      reg1797 <= reg1088[(2'h3):(1'h1)];
                    end
                  if (($unsigned($unsigned({reg1722})) >= reg1108[(3'h6):(1'h0)]))
                    begin
                      reg1798 <= forvar1775;
                      reg1799 <= $unsigned(reg1011);
                      reg1800 <= $signed($unsigned(($unsigned(reg1045) ?
                          reg1083 : (reg1082 | reg1761))));
                      reg1801 <= (reg1796[(2'h3):(1'h0)] <<< {$unsigned(reg1117[(2'h3):(1'h1)])});
                    end
                  else
                    begin
                      reg1798 <= (($unsigned({forvar1751}) + {$signed(reg1008)}) * (8'haa));
                      reg1799 <= ((8'hb3) ^~ reg1695);
                      reg1800 <= (~$signed(reg1747[(1'h1):(1'h0)]));
                    end
                end
            end
          for (forvar1802 = (1'h0); (forvar1802 < (1'h0)); forvar1802 = (forvar1802 + (1'h1)))
            begin
              reg1803 <= reg1006;
              for (forvar1804 = (1'h0); (forvar1804 < (1'h1)); forvar1804 = (forvar1804 + (1'h1)))
                begin
                  for (forvar1805 = (1'h0); (forvar1805 < (1'h0)); forvar1805 = (forvar1805 + (1'h1)))
                    begin
                      reg1806 <= reg1783;
                      reg1807 <= reg1129;
                      reg1808 <= reg1010;
                      reg1809 <= ((~|($signed((8'hae)) ?
                              {forvar1716} : (&reg1132))) ?
                          $unsigned(reg1760[(3'h5):(2'h2)]) : (((reg994 << reg994) >= $signed((8'hb1))) | ((reg1128 >> reg1767) <= $unsigned((8'hba)))));
                    end
                end
              for (forvar1810 = (1'h0); (forvar1810 < (2'h3)); forvar1810 = (forvar1810 + (1'h1)))
                begin
                  for (forvar1811 = (1'h0); (forvar1811 < (2'h3)); forvar1811 = (forvar1811 + (1'h1)))
                    begin
                      reg1812 <= reg1013[(3'h7):(3'h6)];
                    end
                  reg1813 <= (~reg1058[(3'h6):(2'h2)]);
                  reg1814 <= $unsigned($signed(reg1711));
                  for (forvar1815 = (1'h0); (forvar1815 < (1'h1)); forvar1815 = (forvar1815 + (1'h1)))
                    begin
                      reg1816 <= $signed(reg991[(3'h5):(2'h3)]);
                      reg1817 <= $unsigned($unsigned($signed($signed(reg1076))));
                      reg1818 <= $unsigned((reg1008 ?
                          ($unsigned(wire1658) ?
                              reg1087[(3'h6):(2'h3)] : $unsigned(reg1715)) : reg1662[(4'h8):(3'h5)]));
                      reg1819 <= (8'haa);
                    end
                end
              for (forvar1820 = (1'h0); (forvar1820 < (1'h1)); forvar1820 = (forvar1820 + (1'h1)))
                begin
                  if (reg1103)
                    begin
                      reg1821 <= (|(^~$signed({(8'ha4)})));
                      reg1822 <= (!{(&{forvar1715})});
                      reg1823 <= (~reg992);
                      reg1824 <= reg1021[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1821 <= (reg1684[(3'h4):(2'h3)] > ((~^reg1033) + reg1779));
                      reg1822 <= reg1058[(3'h4):(2'h2)];
                    end
                end
            end
          for (forvar1825 = (1'h0); (forvar1825 < (2'h3)); forvar1825 = (forvar1825 + (1'h1)))
            begin
              for (forvar1826 = (1'h0); (forvar1826 < (1'h1)); forvar1826 = (forvar1826 + (1'h1)))
                begin
                  for (forvar1827 = (1'h0); (forvar1827 < (2'h3)); forvar1827 = (forvar1827 + (1'h1)))
                    begin
                      reg1828 <= ((reg1131[(2'h2):(2'h2)] ~^ reg1710[(1'h0):(1'h0)]) <<< (^$unsigned({reg1806})));
                      reg1829 <= forvar1775;
                      reg1830 <= $signed(((reg1813 ?
                          reg1021 : $unsigned(reg1790)) | ($signed(reg1747) ?
                          $unsigned(forvar1804) : (reg1036 ^~ (8'haa)))));
                    end
                  if ($signed(reg1830[(4'hd):(4'hc)]))
                    begin
                      reg1831 <= reg1830;
                      reg1832 <= $unsigned((!{(forvar1757 <<< reg1744)}));
                      reg1833 <= ($unsigned((^$signed(reg1831))) ?
                          (8'hae) : ((~|(^reg1803)) ?
                              (~^$signed(forvar1736)) : {reg1781[(1'h1):(1'h0)]}));
                    end
                  else
                    begin
                      reg1831 <= $unsigned(($unsigned($unsigned(reg1036)) ?
                          reg1747 : {(forvar1729 <<< reg990)}));
                      reg1832 <= $signed(reg1780[(1'h0):(1'h0)]);
                    end
                  if (reg1131[(1'h0):(1'h0)])
                    begin
                      reg1834 <= $unsigned((reg1088 | $signed(reg1693[(3'h4):(1'h1)])));
                      reg1835 <= $unsigned($signed(reg1801[(4'h9):(4'h9)]));
                      reg1836 <= ((&reg1765[(1'h1):(1'h0)]) ?
                          reg1135[(1'h1):(1'h0)] : forvar1729);
                    end
                  else
                    begin
                      reg1834 <= (~&reg1014[(2'h3):(2'h3)]);
                    end
                  for (forvar1837 = (1'h0); (forvar1837 < (2'h2)); forvar1837 = (forvar1837 + (1'h1)))
                    begin
                      reg1838 <= {(!reg1727[(4'h8):(3'h5)])};
                      reg1839 <= reg1835[(4'h9):(3'h6)];
                    end
                end
              for (forvar1840 = (1'h0); (forvar1840 < (2'h2)); forvar1840 = (forvar1840 + (1'h1)))
                begin
                  for (forvar1841 = (1'h0); (forvar1841 < (2'h2)); forvar1841 = (forvar1841 + (1'h1)))
                    begin
                      reg1842 <= forvar1718[(4'ha):(2'h3)];
                      reg1843 <= reg1111[(3'h7):(1'h1)];
                    end
                end
              if (($unsigned($unsigned(((8'hb0) | reg1130))) ?
                  (8'ha1) : reg1137[(4'h8):(1'h1)]))
                begin
                  reg1844 <= (~(-$unsigned((!reg1728))));
                  if ($signed((8'h9f)))
                    begin
                      reg1845 <= (~&reg1729);
                      reg1846 <= $signed($unsigned(((wire985 < reg1000) ?
                          (!reg1824) : (-reg1781))));
                      reg1847 <= ($unsigned(reg1671) ?
                          (&{(|forvar1706)}) : (^~(~^{reg1137})));
                      reg1848 <= ((reg1004[(4'he):(3'h6)] >= $unsigned($signed(forvar1715))) ?
                          ({$unsigned(reg1090)} ?
                              {(reg1144 > (8'h9d))} : (~$unsigned(reg1729))) : $signed(({forvar1805} ?
                              (-reg1830) : (reg1842 - reg1061))));
                    end
                  else
                    begin
                      reg1845 <= (reg1824 ?
                          (!$unsigned({(8'hb7)})) : (((forvar1768 <<< forvar1754) ?
                              forvar1756[(5'h10):(4'he)] : (forvar1737 && (8'h9c))) << (^~{forvar1811})));
                      reg1846 <= $signed({reg1662});
                      reg1847 <= reg1749[(3'h7):(3'h6)];
                    end
                  for (forvar1849 = (1'h0); (forvar1849 < (2'h3)); forvar1849 = (forvar1849 + (1'h1)))
                    begin
                      reg1850 <= ((reg1774 >>> {(reg1747 != (8'hb5))}) * wire984);
                      reg1851 <= $unsigned((!$unsigned(forvar1827)));
                    end
                end
              else
                begin
                  for (forvar1844 = (1'h0); (forvar1844 < (1'h1)); forvar1844 = (forvar1844 + (1'h1)))
                    begin
                      reg1845 <= reg1716;
                    end
                  reg1846 <= reg998;
                  if ((+(reg1016[(4'h8):(1'h1)] > $unsigned($unsigned(reg1144)))))
                    begin
                      reg1847 <= (reg1061 && {((reg1730 >= (8'ha4)) ?
                              (^~reg1683) : reg1127[(1'h0):(1'h0)])});
                      reg1848 <= $signed(reg1753);
                      reg1849 <= $signed((8'ha0));
                      reg1850 <= ((reg1132 ?
                              $signed((reg1813 <<< reg1704)) : {reg1721[(1'h0):(1'h0)]}) ?
                          reg1774[(3'h6):(2'h2)] : reg1839);
                    end
                  else
                    begin
                      reg1847 <= (!(|($unsigned(reg1101) * (^~(8'hba)))));
                    end
                  reg1851 <= (&(+(~&reg990)));
                end
              for (forvar1852 = (1'h0); (forvar1852 < (1'h1)); forvar1852 = (forvar1852 + (1'h1)))
                begin
                  for (forvar1853 = (1'h0); (forvar1853 < (1'h1)); forvar1853 = (forvar1853 + (1'h1)))
                    begin
                      reg1854 <= (~^$unsigned(reg1072[(4'hb):(4'hb)]));
                      reg1855 <= {(|({reg1110} > forvar1837))};
                    end
                  for (forvar1856 = (1'h0); (forvar1856 < (1'h1)); forvar1856 = (forvar1856 + (1'h1)))
                    begin
                      reg1857 <= $signed((!(&(~reg1728))));
                      reg1858 <= (+((&{reg1798}) ?
                          ($signed(reg1704) ?
                              (^~reg1720) : {reg1005}) : reg1022));
                      reg1859 <= (reg1106 && (8'hb1));
                      reg1860 <= $unsigned($signed(({reg1675} ?
                          (~wire1705) : (^~reg1101))));
                    end
                end
            end
        end
    end
  assign wire1861 = (($signed((reg1025 ? reg1770 : reg1670)) ?
                        (8'hac) : reg1062[(3'h7):(1'h0)]) * $signed({reg1660[(4'h8):(2'h3)]}));
  always
    @(posedge clk) begin
      for (forvar1862 = (1'h0); (forvar1862 < (1'h1)); forvar1862 = (forvar1862 + (1'h1)))
        begin
          reg1863 <= (($unsigned($unsigned((8'ha6))) != (-((8'ha0) == reg1844))) ?
              {reg1715[(1'h0):(1'h0)]} : $unsigned((reg1762 ?
                  (^reg1788) : $signed(reg1662))));
          for (forvar1864 = (1'h0); (forvar1864 < (2'h2)); forvar1864 = (forvar1864 + (1'h1)))
            begin
              for (forvar1865 = (1'h0); (forvar1865 < (1'h1)); forvar1865 = (forvar1865 + (1'h1)))
                begin
                  for (forvar1866 = (1'h0); (forvar1866 < (1'h0)); forvar1866 = (forvar1866 + (1'h1)))
                    begin
                      reg1867 <= ({reg1050} ?
                          $unsigned($signed(reg1790[(3'h5):(3'h4)])) : $signed($signed((8'had))));
                      reg1868 <= reg1141;
                      reg1869 <= (reg1027 ?
                          $signed(reg1690[(1'h1):(1'h1)]) : {($signed(reg1850) ?
                                  $signed(reg1763) : $signed(reg1044))});
                    end
                  reg1870 <= reg1064[(3'h6):(3'h5)];
                end
            end
          if ($unsigned((((wire1658 ?
              reg1077 : wire987) <= {reg1035}) | $unsigned((^~reg1061)))))
            begin
              if ((reg1018[(3'h4):(2'h3)] << (reg1676 ?
                  ($signed(reg1755) ~^ (reg1041 < (8'hb1))) : $signed($signed(reg1778)))))
                begin
                  for (forvar1871 = (1'h0); (forvar1871 < (1'h0)); forvar1871 = (forvar1871 + (1'h1)))
                    begin
                      reg1872 <= reg1062;
                      reg1873 <= reg1068[(4'h9):(3'h4)];
                    end
                  if (((reg1722[(4'hc):(2'h2)] ?
                          $unsigned((!forvar1865)) : reg1075) ?
                      reg1019[(4'he):(3'h5)] : reg1064))
                    begin
                      reg1874 <= ($signed(($unsigned((8'ha6)) ?
                              reg1684 : $signed(reg1054))) ?
                          $unsigned(((reg1760 ?
                              reg1025 : (8'ha1)) << $signed(reg1748))) : (reg991[(1'h1):(1'h0)] ^~ (reg1757 ?
                              reg1023[(3'h6):(2'h2)] : reg1836[(3'h5):(3'h4)])));
                      reg1875 <= reg1836[(3'h5):(2'h2)];
                      reg1876 <= (|(^(^reg1858)));
                      reg1877 <= $unsigned((|$signed({reg1748})));
                    end
                  else
                    begin
                      reg1874 <= ((8'hb4) != $unsigned($unsigned((reg1070 ?
                          reg1759 : reg1809))));
                      reg1875 <= $unsigned((reg1848[(3'h5):(2'h2)] >= reg1809[(4'hb):(3'h5)]));
                    end
                  for (forvar1878 = (1'h0); (forvar1878 < (2'h3)); forvar1878 = (forvar1878 + (1'h1)))
                    begin
                      reg1879 <= (reg1795 >> (~($unsigned((8'ha2)) ^ (^~reg1111))));
                      reg1880 <= (~^$unsigned((((8'ha5) ? reg1075 : reg1132) ?
                          $unsigned(reg1798) : (wire985 | reg1859))));
                      reg1881 <= $signed({reg1717});
                      reg1882 <= reg1112;
                    end
                end
              else
                begin
                  for (forvar1871 = (1'h0); (forvar1871 < (2'h2)); forvar1871 = (forvar1871 + (1'h1)))
                    begin
                      reg1872 <= {((~&$unsigned(reg1042)) ?
                              $unsigned((^~reg1772)) : {(8'hab)})};
                      reg1873 <= reg1023;
                    end
                  for (forvar1874 = (1'h0); (forvar1874 < (1'h0)); forvar1874 = (forvar1874 + (1'h1)))
                    begin
                      reg1875 <= (8'hb6);
                      reg1876 <= reg1085[(3'h4):(1'h0)];
                    end
                  for (forvar1877 = (1'h0); (forvar1877 < (2'h3)); forvar1877 = (forvar1877 + (1'h1)))
                    begin
                      reg1878 <= ($signed(reg1021[(2'h2):(1'h1)]) ?
                          reg1037[(2'h3):(2'h3)] : ({$unsigned(reg1834)} & reg1113));
                      reg1879 <= (~|({(reg1037 ? reg1068 : reg1075)} ?
                          reg1050 : (reg1834 >= $unsigned(reg1003))));
                      reg1880 <= reg989[(2'h2):(1'h1)];
                      reg1881 <= $signed(reg1089[(1'h1):(1'h0)]);
                    end
                end
              for (forvar1883 = (1'h0); (forvar1883 < (2'h2)); forvar1883 = (forvar1883 + (1'h1)))
                begin
                  for (forvar1884 = (1'h0); (forvar1884 < (2'h2)); forvar1884 = (forvar1884 + (1'h1)))
                    begin
                      reg1885 <= ((reg1007[(3'h4):(2'h3)] >> (&(~reg1774))) ?
                          (^~(!(reg1710 ^ reg991))) : $signed(reg1123));
                    end
                end
              reg1886 <= reg1690[(3'h6):(3'h6)];
              for (forvar1887 = (1'h0); (forvar1887 < (2'h3)); forvar1887 = (forvar1887 + (1'h1)))
                begin
                  for (forvar1888 = (1'h0); (forvar1888 < (1'h0)); forvar1888 = (forvar1888 + (1'h1)))
                    begin
                      reg1889 <= wire1658[(3'h5):(1'h1)];
                      reg1890 <= reg1671[(2'h3):(1'h1)];
                      reg1891 <= $unsigned($signed($unsigned(wire982)));
                      reg1892 <= $unsigned((!(reg1127[(2'h2):(1'h1)] ?
                          (|(8'hb2)) : $unsigned(reg1037))));
                    end
                  reg1893 <= reg1668;
                end
            end
          else
            begin
              if ((reg1797[(3'h6):(1'h0)] > {((+reg1018) ?
                      {reg1131} : (~^reg1091))}))
                begin
                  if (reg1117)
                    begin
                      reg1871 <= $signed({$unsigned(reg1126[(3'h4):(1'h1)])});
                      reg1872 <= reg1855;
                      reg1873 <= ((^$signed((-reg1023))) & $unsigned($signed(forvar1864)));
                    end
                  else
                    begin
                      reg1871 <= {reg1673};
                    end
                  for (forvar1874 = (1'h0); (forvar1874 < (1'h0)); forvar1874 = (forvar1874 + (1'h1)))
                    begin
                      reg1875 <= $signed({(~&(reg1048 ? (8'h9e) : (8'hb2)))});
                    end
                  if ((($unsigned((+(8'hb7))) ?
                      {$unsigned(reg1785)} : wire1861[(3'h6):(2'h3)]) >> reg1115))
                    begin
                      reg1876 <= reg1081;
                      reg1877 <= {$unsigned(reg1123[(1'h1):(1'h0)])};
                    end
                  else
                    begin
                      reg1876 <= {(&reg1718)};
                      reg1877 <= ($signed(((8'hb9) != (+wire983))) <= reg998[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  reg1871 <= (reg1877[(4'h8):(2'h2)] >= $unsigned((8'haf)));
                  for (forvar1872 = (1'h0); (forvar1872 < (1'h0)); forvar1872 = (forvar1872 + (1'h1)))
                    begin
                      reg1873 <= $signed(reg1700[(1'h0):(1'h0)]);
                      reg1874 <= $unsigned(reg1675[(3'h6):(1'h0)]);
                      reg1875 <= (^~$signed($unsigned((~&reg1103))));
                    end
                end
              for (forvar1878 = (1'h0); (forvar1878 < (1'h1)); forvar1878 = (forvar1878 + (1'h1)))
                begin
                  for (forvar1879 = (1'h0); (forvar1879 < (1'h1)); forvar1879 = (forvar1879 + (1'h1)))
                    begin
                      reg1880 <= (!reg1679[(1'h1):(1'h1)]);
                      reg1881 <= $unsigned((({(8'h9f)} ~^ $unsigned(forvar1883)) ?
                          (8'ha6) : reg1034[(4'hc):(4'hb)]));
                      reg1882 <= ($signed($signed((-reg998))) * reg1738);
                      reg1883 <= $signed($signed(($unsigned(reg991) ?
                          (+reg1101) : {reg1065})));
                    end
                  for (forvar1884 = (1'h0); (forvar1884 < (2'h3)); forvar1884 = (forvar1884 + (1'h1)))
                    begin
                      reg1885 <= reg1702[(4'h9):(3'h6)];
                      reg1886 <= $signed($unsigned((reg1858[(3'h5):(1'h0)] ~^ {(8'hb6)})));
                    end
                  if ($unsigned($unsigned(reg1809[(2'h2):(1'h1)])))
                    begin
                      reg1887 <= (-$signed((~|$signed(forvar1888))));
                      reg1888 <= $signed(reg1035);
                    end
                  else
                    begin
                      reg1887 <= $unsigned($unsigned((~^$signed(reg1844))));
                      reg1888 <= (((+reg1735[(1'h0):(1'h0)]) >= (~|reg1812)) < $signed((((8'hb7) >= reg1662) - $unsigned(reg1869))));
                    end
                  for (forvar1889 = (1'h0); (forvar1889 < (2'h3)); forvar1889 = (forvar1889 + (1'h1)))
                    begin
                      reg1890 <= (^~($signed(reg1879[(3'h7):(2'h2)]) * (reg1117[(3'h4):(2'h3)] ?
                          (reg1877 << reg1881) : (reg1757 ^ reg1769))));
                      reg1891 <= $signed($signed(wire986[(1'h1):(1'h1)]));
                    end
                end
              for (forvar1892 = (1'h0); (forvar1892 < (1'h1)); forvar1892 = (forvar1892 + (1'h1)))
                begin
                  for (forvar1893 = (1'h0); (forvar1893 < (2'h2)); forvar1893 = (forvar1893 + (1'h1)))
                    begin
                      reg1894 <= $unsigned((-$signed((~reg1110))));
                      reg1895 <= reg1015[(4'h9):(3'h5)];
                      reg1896 <= $unsigned({(reg1085[(4'h8):(1'h1)] ?
                              reg998[(2'h3):(2'h2)] : {reg1731})});
                      reg1897 <= ($signed(((reg1666 * reg1871) ?
                              $unsigned((8'ha1)) : {wire981})) ?
                          (($signed(reg1082) <<< $unsigned((8'hac))) ?
                              $signed((~reg1061)) : (~^$signed(reg1876))) : (^$signed((^reg1126))));
                    end
                  if ((reg1663[(1'h0):(1'h0)] != (&((reg1677 != reg1892) ?
                      reg1138 : $signed((8'hb6))))))
                    begin
                      reg1898 <= ({reg1075} ?
                          $unsigned((&$signed((8'hb0)))) : (-$signed(reg1050)));
                      reg1899 <= reg1129;
                      reg1900 <= ({$signed((~&reg1835))} <<< {((reg1842 ?
                                  reg1838 : reg1734) ?
                              (~reg1003) : $signed(reg1873))});
                      reg1901 <= ((reg1842[(3'h7):(1'h1)] << (8'ha8)) && (8'hb8));
                    end
                  else
                    begin
                      reg1898 <= $signed($unsigned($signed(reg1098[(3'h4):(3'h4)])));
                      reg1899 <= (wire986[(1'h0):(1'h0)] * (reg1673 + {reg1060[(1'h0):(1'h0)]}));
                      reg1900 <= (~&reg1818[(3'h7):(3'h6)]);
                      reg1901 <= $unsigned((~^{$unsigned(reg1014)}));
                    end
                  reg1902 <= ((|((reg1738 < reg1828) + $signed((8'ha9)))) ?
                      (((8'hb9) << ((8'h9c) <= reg1665)) ~^ (reg1900 ?
                          (reg1814 * reg1769) : $signed(reg1900))) : reg1014);
                  if (wire987)
                    begin
                      reg1903 <= ({(reg1110 ?
                              ((8'had) ?
                                  reg1022 : reg1037) : $unsigned(reg1708))} && reg1832);
                      reg1904 <= (^~{$unsigned(reg1819)});
                    end
                  else
                    begin
                      reg1903 <= $unsigned($signed({(|reg1085)}));
                      reg1904 <= (((forvar1874 ^ ((8'hae) <= reg1123)) ?
                          (&reg1761) : reg1063) || ((~^$signed(reg1836)) ?
                          ((forvar1884 ?
                              (8'ha8) : forvar1883) <= (8'ha3)) : ((reg1899 ?
                              reg1144 : reg1003) * reg1041[(1'h0):(1'h0)])));
                      reg1905 <= {reg1765};
                      reg1906 <= ({$signed((reg1135 ^ reg1839))} ?
                          $signed($unsigned(reg1886[(1'h1):(1'h0)])) : reg1144);
                    end
                end
            end
        end
    end
  assign wire1907 = ($unsigned(reg1125) && ((reg1145 ?
                        reg1093[(3'h6):(2'h2)] : (reg1706 | reg1130)) | $unsigned($signed((8'had)))));
  assign wire1908 = (({reg1765[(1'h1):(1'h1)]} <= $unsigned($unsigned(reg1760))) <<< ({((8'h9e) ?
                            reg1757 : (8'hab))} + ($unsigned(reg1754) ?
                        ((8'haa) == reg1679) : (reg1026 << (8'ha8)))));
  always
    @(posedge clk) begin
      for (forvar1909 = (1'h0); (forvar1909 < (2'h2)); forvar1909 = (forvar1909 + (1'h1)))
        begin
          reg1910 <= {(&reg1144[(2'h3):(2'h2)])};
        end
      reg1911 <= $unsigned(({reg1756} & reg1677));
      for (forvar1912 = (1'h0); (forvar1912 < (1'h1)); forvar1912 = (forvar1912 + (1'h1)))
        begin
          for (forvar1913 = (1'h0); (forvar1913 < (2'h2)); forvar1913 = (forvar1913 + (1'h1)))
            begin
              reg1914 <= (+reg1035[(1'h1):(1'h1)]);
            end
          if (($unsigned($unsigned(reg1733)) & (~&reg1706)))
            begin
              for (forvar1915 = (1'h0); (forvar1915 < (2'h3)); forvar1915 = (forvar1915 + (1'h1)))
                begin
                  if (reg1798[(4'h9):(4'h9)])
                    begin
                      reg1916 <= (reg1133 ^~ (8'hb2));
                    end
                  else
                    begin
                      reg1916 <= {{reg1090[(1'h0):(1'h0)]}};
                      reg1917 <= ($signed(reg1771) ?
                          {reg1129[(4'h9):(2'h2)]} : ({$unsigned((8'h9f))} >> {((8'had) << (8'haa))}));
                    end
                  for (forvar1918 = (1'h0); (forvar1918 < (1'h1)); forvar1918 = (forvar1918 + (1'h1)))
                    begin
                      reg1919 <= (^~$unsigned((reg1064[(2'h2):(1'h0)] >= $signed((8'ha8)))));
                      reg1920 <= (($signed(reg1066[(1'h0):(1'h0)]) ?
                              forvar1909[(4'h9):(3'h5)] : $unsigned((8'ha5))) ?
                          (($signed(reg1783) ?
                                  forvar1913 : reg989[(2'h3):(1'h1)]) ?
                              (-reg1730) : {$signed((8'hac))}) : wire985[(2'h3):(2'h3)]);
                    end
                  reg1921 <= (reg1910 <<< reg1010);
                end
            end
          else
            begin
              if (forvar1913)
                begin
                  for (forvar1915 = (1'h0); (forvar1915 < (2'h2)); forvar1915 = (forvar1915 + (1'h1)))
                    begin
                      reg1916 <= $unsigned({((reg989 ? (8'ha3) : reg1870) ?
                              (reg1025 != reg1745) : $signed(reg1130))});
                      reg1917 <= ($unsigned(reg1679) ^~ reg1760[(2'h3):(2'h3)]);
                      reg1918 <= (~(~^$unsigned((~(8'h9e)))));
                      reg1919 <= $signed((((reg1854 ? reg1124 : (8'hb1)) ?
                              (reg1854 & reg1090) : $signed(reg1724)) ?
                          {(~|reg1843)} : $unsigned({reg1115})));
                    end
                  if (reg1736)
                    begin
                      reg1920 <= (reg991[(3'h5):(2'h2)] <= forvar1918[(3'h5):(1'h1)]);
                      reg1921 <= reg1056;
                      reg1922 <= $unsigned((8'hab));
                      reg1923 <= {(wire986[(2'h2):(1'h1)] ?
                              $unsigned(reg1714) : $signed($unsigned(reg1902)))};
                    end
                  else
                    begin
                      reg1920 <= {$unsigned(reg1784)};
                    end
                  for (forvar1924 = (1'h0); (forvar1924 < (2'h3)); forvar1924 = (forvar1924 + (1'h1)))
                    begin
                      reg1925 <= reg1064[(3'h4):(1'h0)];
                      reg1926 <= $signed((^(reg1030 ?
                          $unsigned(reg1715) : $signed(reg1739))));
                    end
                end
              else
                begin
                  reg1915 <= ($signed(reg1018) ?
                      $signed({$signed(reg1738)}) : {reg1739});
                  for (forvar1916 = (1'h0); (forvar1916 < (1'h0)); forvar1916 = (forvar1916 + (1'h1)))
                    begin
                      reg1917 <= (((~(~reg1709)) ?
                          ((~|reg1716) ?
                              (reg1098 ?
                                  reg1796 : reg1718) : reg1008) : $signed($signed((8'hba)))) != (-((~wire1861) ^ $unsigned(reg1000))));
                      reg1918 <= (~&(&{reg1742[(3'h4):(3'h4)]}));
                      reg1919 <= reg1876[(3'h5):(2'h3)];
                      reg1920 <= $signed($signed(((8'hae) ~^ $unsigned(reg1747))));
                    end
                  for (forvar1921 = (1'h0); (forvar1921 < (1'h1)); forvar1921 = (forvar1921 + (1'h1)))
                    begin
                      reg1922 <= ($unsigned(($unsigned(reg1902) ?
                          reg1117[(3'h4):(2'h3)] : reg1054)) << ({reg1798[(4'h9):(3'h4)]} > (|reg1723)));
                    end
                end
              reg1927 <= wire1908[(2'h3):(1'h0)];
              for (forvar1928 = (1'h0); (forvar1928 < (1'h1)); forvar1928 = (forvar1928 + (1'h1)))
                begin
                  for (forvar1929 = (1'h0); (forvar1929 < (1'h1)); forvar1929 = (forvar1929 + (1'h1)))
                    begin
                      reg1930 <= reg1129;
                      reg1931 <= reg1741;
                      reg1932 <= ((forvar1929[(1'h0):(1'h0)] ?
                              (reg1757 ?
                                  $signed(reg1105) : ((8'ha4) ?
                                      reg1012 : (8'h9f))) : $unsigned($unsigned(reg1745))) ?
                          $unsigned($signed(reg1113[(4'h9):(2'h2)])) : $signed((^(reg1844 <<< reg990))));
                      reg1933 <= ((($signed(reg1773) || (reg1813 ?
                              (8'hb0) : (8'hb2))) << (^$unsigned(reg1737))) ?
                          $signed((~^$signed(reg1690))) : (+{(&reg1772)}));
                    end
                  for (forvar1934 = (1'h0); (forvar1934 < (1'h1)); forvar1934 = (forvar1934 + (1'h1)))
                    begin
                      reg1935 <= (reg1823[(4'ha):(2'h3)] <= $unsigned(({reg1051} & $unsigned(reg1011))));
                      reg1936 <= $unsigned({((!wire987) ?
                              {reg1104} : reg1108)});
                      reg1937 <= $unsigned(((^~$unsigned(reg1725)) ?
                          ($unsigned((8'hb3)) < $unsigned((8'ha3))) : $signed(reg1890[(3'h7):(3'h6)])));
                    end
                  for (forvar1938 = (1'h0); (forvar1938 < (1'h0)); forvar1938 = (forvar1938 + (1'h1)))
                    begin
                      reg1939 <= $signed((8'hb3));
                      reg1940 <= ((~^$signed((+reg1771))) & (((reg1760 ^~ reg1819) + $unsigned(reg1044)) ?
                          (^~$unsigned((8'hb6))) : $unsigned(reg1703[(4'h9):(2'h2)])));
                      reg1941 <= $signed((!$signed(reg1040[(3'h5):(3'h5)])));
                    end
                  for (forvar1942 = (1'h0); (forvar1942 < (2'h2)); forvar1942 = (forvar1942 + (1'h1)))
                    begin
                      reg1943 <= reg1670[(4'hc):(3'h5)];
                      reg1944 <= {{((reg1824 ?
                                  (8'haa) : reg1739) >>> (!reg1873))}};
                      reg1945 <= {$signed(((reg1096 ? reg1892 : forvar1918) ?
                              {forvar1912} : (~^reg1126)))};
                    end
                end
            end
          if ((reg1129[(4'ha):(3'h5)] ?
              reg1107 : ({reg1796[(1'h0):(1'h0)]} * ({reg1849} != reg1712[(3'h6):(3'h5)]))))
            begin
              if ((+(reg1063[(3'h4):(3'h4)] ?
                  $signed(reg1119[(3'h5):(1'h1)]) : ($unsigned(reg1664) | reg1009[(4'ha):(1'h0)]))))
                begin
                  for (forvar1946 = (1'h0); (forvar1946 < (2'h2)); forvar1946 = (forvar1946 + (1'h1)))
                    begin
                      reg1947 <= reg1091[(4'hf):(4'h9)];
                      reg1948 <= ($unsigned((~&$signed(reg1838))) ?
                          (~&(-reg1779)) : $signed(((reg1740 == reg1750) ?
                              (8'ha6) : $unsigned(reg1879))));
                    end
                  reg1949 <= ((|((reg1936 ? reg1859 : reg1048) ?
                          (reg1941 >>> reg1877) : (!reg1100))) ?
                      wire987 : $unsigned((~|$signed((8'haf)))));
                  for (forvar1950 = (1'h0); (forvar1950 < (1'h1)); forvar1950 = (forvar1950 + (1'h1)))
                    begin
                      reg1951 <= $signed((reg1712[(3'h4):(1'h1)] <= ($signed(reg1756) * $unsigned(wire1907))));
                      reg1952 <= $unsigned((($signed(reg1131) >= wire981[(4'h8):(3'h6)]) <= (!reg1117[(3'h5):(1'h1)])));
                      reg1953 <= reg1814;
                    end
                end
              else
                begin
                  if ({$signed((~&reg1806[(4'h8):(4'h8)]))})
                    begin
                      reg1946 <= reg1086[(2'h2):(1'h1)];
                      reg1947 <= reg1824;
                      reg1948 <= (+$unsigned({reg1670[(3'h4):(3'h4)]}));
                      reg1949 <= reg1851[(4'he):(4'hd)];
                    end
                  else
                    begin
                      reg1946 <= {(~|$signed((reg1953 ? reg1758 : reg1067)))};
                      reg1947 <= $unsigned((8'ha5));
                      reg1948 <= (^~reg1891[(1'h0):(1'h0)]);
                    end
                end
              if (reg1001)
                begin
                  if (((((reg1889 ? (8'h9d) : reg1822) ?
                          reg1764 : $unsigned(reg1880)) ^ wire987) ?
                      ($unsigned(reg995[(2'h2):(1'h0)]) ?
                          (~(-reg1935)) : $unsigned((reg1761 ?
                              reg1868 : reg1668))) : ((-$signed(reg1888)) ?
                          (reg1081 ~^ reg1768[(1'h1):(1'h0)]) : reg1105)))
                    begin
                      reg1954 <= ($signed(((reg1788 ? (8'hba) : (8'hb9)) ?
                              $unsigned(reg1139) : $signed(reg1911))) ?
                          (~&(reg1874 ?
                              $signed(reg1675) : $signed(reg1728))) : (8'had));
                    end
                  else
                    begin
                      reg1954 <= (|$signed((reg1729[(4'h9):(3'h7)] ?
                          (reg1874 ? reg1808 : reg1718) : (!reg1757))));
                      reg1955 <= reg1109[(1'h0):(1'h0)];
                    end
                  for (forvar1956 = (1'h0); (forvar1956 < (1'h0)); forvar1956 = (forvar1956 + (1'h1)))
                    begin
                      reg1957 <= $unsigned(reg1801[(4'ha):(2'h3)]);
                      reg1958 <= {$unsigned(($unsigned((8'hac)) ?
                              (^reg1834) : ((8'hb2) >= reg1754)))};
                      reg1959 <= $unsigned(($unsigned(reg1080[(3'h4):(1'h1)]) & (!(forvar1915 ?
                          reg1882 : reg992))));
                    end
                  reg1960 <= (!($signed((&reg1892)) != reg1011[(3'h5):(1'h0)]));
                  for (forvar1961 = (1'h0); (forvar1961 < (1'h1)); forvar1961 = (forvar1961 + (1'h1)))
                    begin
                      reg1962 <= ($unsigned($signed(reg1045)) ?
                          reg1104 : (~|{$unsigned((8'hae))}));
                      reg1963 <= ($signed(((reg1839 | reg1819) * $unsigned((8'ha3)))) ?
                          {({reg1692} >>> reg1107)} : ((8'ha4) + {(~|(8'ha7))}));
                      reg1964 <= reg1958[(1'h1):(1'h1)];
                      reg1965 <= $unsigned(reg1930);
                    end
                end
              else
                begin
                  reg1954 <= (reg1038[(4'h8):(3'h5)] << reg1783[(1'h0):(1'h0)]);
                end
              reg1966 <= reg1056[(1'h0):(1'h0)];
            end
          else
            begin
              if ($signed((~|((-reg1763) != {reg1730}))))
                begin
                  for (forvar1946 = (1'h0); (forvar1946 < (1'h1)); forvar1946 = (forvar1946 + (1'h1)))
                    begin
                      reg1947 <= $unsigned(((~|(reg1886 <<< reg1139)) ?
                          {reg1096[(3'h4):(2'h2)]} : $unsigned((reg1770 ?
                              reg1795 : reg1870))));
                    end
                  reg1948 <= reg1736;
                  reg1949 <= (^~($unsigned({reg1102}) - (^$unsigned(reg1100))));
                  if (($unsigned((&$signed((8'ha3)))) ?
                      reg1745[(2'h2):(1'h0)] : (8'hab)))
                    begin
                      reg1950 <= (reg1739[(3'h4):(1'h1)] ?
                          reg1838 : (($signed(reg1944) >>> {reg1809}) + {(reg1829 <<< reg1116)}));
                      reg1951 <= (~reg1786);
                      reg1952 <= {$unsigned($signed((-forvar1912)))};
                    end
                  else
                    begin
                      reg1950 <= reg1874[(4'h9):(3'h6)];
                      reg1951 <= (~|(reg1022 - reg1007[(3'h5):(1'h0)]));
                      reg1952 <= $unsigned($signed($unsigned(reg1001[(2'h2):(2'h2)])));
                      reg1953 <= (!reg1127[(2'h2):(1'h0)]);
                    end
                end
              else
                begin
                  if (reg1095[(4'hf):(4'hc)])
                    begin
                      reg1946 <= $unsigned($unsigned(((8'h9e) ?
                          {reg1888} : (reg1012 ? reg1829 : reg1880))));
                      reg1947 <= (+reg1108);
                      reg1948 <= reg1005;
                    end
                  else
                    begin
                      reg1946 <= ($unsigned($signed(((8'hba) * (8'hae)))) ?
                          ($unsigned((~|reg1133)) ?
                              reg1122[(4'he):(4'he)] : $unsigned($unsigned(reg1833))) : reg1813);
                      reg1947 <= reg1715[(2'h2):(1'h1)];
                    end
                end
            end
        end
    end
  assign wire1967 = {{reg1822[(1'h0):(1'h0)]}};
  assign wire1968 = reg1860[(1'h1):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1148
#(parameter param1657 = (((&{(8'h9f)}) ? (((8'ha0) ? (8'hb3) : (8'h9d)) ? (&(8'hb8)) : {(8'h9f)}) : (&((8'ha8) ? (8'hb8) : (8'hb1)))) ? (({(8'haa)} ? ((8'h9e) << (8'ha7)) : (^~(8'hb1))) ? ((-(8'hb9)) >= (~^(8'ha8))) : (^{(8'ha0)})) : (((~|(8'had)) ? ((8'h9f) < (8'h9d)) : {(8'ha1)}) + {((8'h9f) ~^ (8'h9d))})))
(y, clk, wire1153, wire1152, wire1151, wire1150, wire1149);
  output wire [(32'h143e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire1153;
  input wire signed [(4'hf):(1'h0)] wire1152;
  input wire signed [(3'h7):(1'h0)] wire1151;
  input wire [(4'hd):(1'h0)] wire1150;
  input wire [(4'hf):(1'h0)] wire1149;
  wire signed [(4'hd):(1'h0)] wire1656;
  wire signed [(4'hc):(1'h0)] wire1655;
  wire [(4'hb):(1'h0)] wire1464;
  wire signed [(2'h2):(1'h0)] wire1255;
  wire [(4'h9):(1'h0)] wire1254;
  wire [(4'ha):(1'h0)] wire1159;
  wire signed [(4'h9):(1'h0)] wire1158;
  wire [(4'hd):(1'h0)] wire1157;
  wire [(4'hc):(1'h0)] wire1156;
  wire [(4'hd):(1'h0)] wire1155;
  wire [(4'hc):(1'h0)] wire1154;
  reg signed [(3'h6):(1'h0)] reg1633 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1626 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1625 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1654 = (1'h0);
  reg [(3'h7):(1'h0)] reg1652 = (1'h0);
  reg [(5'h10):(1'h0)] reg1651 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1650 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1649 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1648 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1647 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1646 = (1'h0);
  reg [(3'h5):(1'h0)] reg1645 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1643 = (1'h0);
  reg [(3'h5):(1'h0)] reg1642 = (1'h0);
  reg [(2'h2):(1'h0)] reg1641 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1637 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1635 = (1'h0);
  reg [(2'h3):(1'h0)] reg1640 = (1'h0);
  reg [(4'hf):(1'h0)] reg1639 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1638 = (1'h0);
  reg [(4'ha):(1'h0)] reg1636 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1634 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1632 = (1'h0);
  reg [(2'h3):(1'h0)] reg1631 = (1'h0);
  reg [(3'h6):(1'h0)] reg1630 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1629 = (1'h0);
  reg [(3'h4):(1'h0)] reg1628 = (1'h0);
  reg [(2'h2):(1'h0)] reg1627 = (1'h0);
  reg [(4'h9):(1'h0)] reg1624 = (1'h0);
  reg [(2'h2):(1'h0)] reg1623 = (1'h0);
  reg [(5'h10):(1'h0)] reg1622 = (1'h0);
  reg [(2'h3):(1'h0)] reg1565 = (1'h0);
  reg [(3'h5):(1'h0)] reg1564 = (1'h0);
  reg [(4'hb):(1'h0)] reg1559 = (1'h0);
  reg [(3'h7):(1'h0)] reg1558 = (1'h0);
  reg [(3'h5):(1'h0)] reg1549 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1545 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1542 = (1'h0);
  reg [(4'hf):(1'h0)] reg1539 = (1'h0);
  reg [(3'h6):(1'h0)] reg1530 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1619 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1618 = (1'h0);
  reg [(3'h4):(1'h0)] reg1616 = (1'h0);
  reg [(4'he):(1'h0)] reg1615 = (1'h0);
  reg [(4'he):(1'h0)] reg1614 = (1'h0);
  reg [(4'h9):(1'h0)] reg1613 = (1'h0);
  reg [(4'hb):(1'h0)] reg1611 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1610 = (1'h0);
  reg [(5'h10):(1'h0)] reg1609 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1608 = (1'h0);
  reg [(2'h3):(1'h0)] reg1607 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1606 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1605 = (1'h0);
  reg [(4'h9):(1'h0)] reg1602 = (1'h0);
  reg [(2'h2):(1'h0)] reg1601 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1604 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1603 = (1'h0);
  reg [(4'hc):(1'h0)] reg1600 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1599 = (1'h0);
  reg [(3'h7):(1'h0)] reg1598 = (1'h0);
  reg [(2'h3):(1'h0)] reg1597 = (1'h0);
  reg [(4'hb):(1'h0)] reg1595 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1594 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1593 = (1'h0);
  reg [(4'hb):(1'h0)] reg1592 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1590 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1589 = (1'h0);
  reg [(3'h4):(1'h0)] reg1588 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1586 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1585 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1584 = (1'h0);
  reg [(3'h6):(1'h0)] reg1583 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1582 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1581 = (1'h0);
  reg [(3'h5):(1'h0)] reg1579 = (1'h0);
  reg [(4'hb):(1'h0)] reg1578 = (1'h0);
  reg [(2'h3):(1'h0)] reg1577 = (1'h0);
  reg [(2'h2):(1'h0)] reg1576 = (1'h0);
  reg [(4'h9):(1'h0)] reg1573 = (1'h0);
  reg [(4'hd):(1'h0)] reg1572 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1570 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1569 = (1'h0);
  reg [(3'h5):(1'h0)] reg1568 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1567 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1566 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1563 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1562 = (1'h0);
  reg [(4'hf):(1'h0)] reg1561 = (1'h0);
  reg [(3'h4):(1'h0)] reg1560 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1557 = (1'h0);
  reg [(4'hb):(1'h0)] reg1556 = (1'h0);
  reg [(2'h3):(1'h0)] reg1555 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1554 = (1'h0);
  reg [(4'hd):(1'h0)] reg1553 = (1'h0);
  reg [(3'h7):(1'h0)] reg1552 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1551 = (1'h0);
  reg [(4'hf):(1'h0)] reg1550 = (1'h0);
  reg [(5'h10):(1'h0)] reg1548 = (1'h0);
  reg [(2'h3):(1'h0)] reg1547 = (1'h0);
  reg [(4'hb):(1'h0)] reg1544 = (1'h0);
  reg [(2'h2):(1'h0)] reg1543 = (1'h0);
  reg [(2'h2):(1'h0)] reg1541 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1540 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1538 = (1'h0);
  reg [(4'h9):(1'h0)] reg1537 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1536 = (1'h0);
  reg [(2'h2):(1'h0)] reg1535 = (1'h0);
  reg [(3'h4):(1'h0)] reg1534 = (1'h0);
  reg [(4'ha):(1'h0)] reg1533 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1532 = (1'h0);
  reg [(4'h8):(1'h0)] reg1531 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1529 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1503 = (1'h0);
  reg [(4'ha):(1'h0)] reg1527 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1526 = (1'h0);
  reg [(4'hc):(1'h0)] reg1525 = (1'h0);
  reg [(4'ha):(1'h0)] reg1524 = (1'h0);
  reg [(3'h4):(1'h0)] reg1523 = (1'h0);
  reg [(4'hc):(1'h0)] reg1520 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1519 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1518 = (1'h0);
  reg [(2'h3):(1'h0)] reg1514 = (1'h0);
  reg [(3'h5):(1'h0)] reg1508 = (1'h0);
  reg [(4'he):(1'h0)] reg1517 = (1'h0);
  reg [(4'h8):(1'h0)] reg1516 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1515 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1513 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1512 = (1'h0);
  reg [(3'h4):(1'h0)] reg1511 = (1'h0);
  reg [(2'h2):(1'h0)] reg1510 = (1'h0);
  reg [(4'hd):(1'h0)] reg1509 = (1'h0);
  reg [(3'h7):(1'h0)] reg1507 = (1'h0);
  reg [(4'h9):(1'h0)] reg1506 = (1'h0);
  reg [(4'hd):(1'h0)] reg1505 = (1'h0);
  reg [(3'h5):(1'h0)] reg1504 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1502 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1501 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1500 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1499 = (1'h0);
  reg [(2'h3):(1'h0)] reg1498 = (1'h0);
  reg [(4'ha):(1'h0)] reg1496 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1495 = (1'h0);
  reg [(3'h4):(1'h0)] reg1494 = (1'h0);
  reg [(3'h5):(1'h0)] reg1493 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1490 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1492 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1491 = (1'h0);
  reg [(4'h8):(1'h0)] reg1489 = (1'h0);
  reg [(3'h6):(1'h0)] reg1488 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1487 = (1'h0);
  reg [(4'h9):(1'h0)] reg1486 = (1'h0);
  reg [(4'hc):(1'h0)] reg1485 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1483 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1482 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1481 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1480 = (1'h0);
  reg [(4'h9):(1'h0)] reg1479 = (1'h0);
  reg [(3'h7):(1'h0)] reg1478 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1477 = (1'h0);
  reg [(4'he):(1'h0)] reg1476 = (1'h0);
  reg [(4'he):(1'h0)] reg1474 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1473 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1472 = (1'h0);
  reg [(4'h8):(1'h0)] reg1470 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1466 = (1'h0);
  reg [(3'h4):(1'h0)] reg1468 = (1'h0);
  reg [(2'h3):(1'h0)] reg1467 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1463 = (1'h0);
  reg [(4'hc):(1'h0)] reg1462 = (1'h0);
  reg [(4'hd):(1'h0)] reg1461 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1459 = (1'h0);
  reg [(4'h9):(1'h0)] reg1458 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1457 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1456 = (1'h0);
  reg [(4'hd):(1'h0)] reg1453 = (1'h0);
  reg [(4'ha):(1'h0)] reg1452 = (1'h0);
  reg [(3'h5):(1'h0)] reg1451 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1448 = (1'h0);
  reg [(4'he):(1'h0)] reg1447 = (1'h0);
  reg [(4'h9):(1'h0)] reg1446 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1445 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1444 = (1'h0);
  reg [(4'hd):(1'h0)] reg1442 = (1'h0);
  reg [(4'h8):(1'h0)] reg1441 = (1'h0);
  reg [(4'ha):(1'h0)] reg1440 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1438 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1425 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1434 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1432 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1431 = (1'h0);
  reg [(4'hc):(1'h0)] reg1430 = (1'h0);
  reg [(3'h5):(1'h0)] reg1429 = (1'h0);
  reg [(4'ha):(1'h0)] reg1428 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1426 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1424 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1423 = (1'h0);
  reg [(3'h6):(1'h0)] reg1422 = (1'h0);
  reg [(4'h8):(1'h0)] reg1421 = (1'h0);
  reg [(2'h3):(1'h0)] reg1419 = (1'h0);
  reg [(5'h10):(1'h0)] reg1418 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1417 = (1'h0);
  reg [(2'h3):(1'h0)] reg1415 = (1'h0);
  reg [(4'h8):(1'h0)] reg1414 = (1'h0);
  reg [(4'hd):(1'h0)] reg1413 = (1'h0);
  reg [(3'h6):(1'h0)] reg1409 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1412 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1411 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1410 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1408 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1407 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1406 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1405 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1404 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1403 = (1'h0);
  reg [(3'h5):(1'h0)] reg1401 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1400 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1399 = (1'h0);
  reg [(5'h10):(1'h0)] reg1398 = (1'h0);
  reg [(4'hd):(1'h0)] reg1397 = (1'h0);
  reg [(4'hf):(1'h0)] reg1396 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1394 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1386 = (1'h0);
  reg [(3'h6):(1'h0)] reg1391 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1390 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1389 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1388 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1387 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1385 = (1'h0);
  reg [(4'hc):(1'h0)] reg1384 = (1'h0);
  reg [(3'h4):(1'h0)] reg1383 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1382 = (1'h0);
  reg [(3'h4):(1'h0)] reg1381 = (1'h0);
  reg [(2'h2):(1'h0)] reg1380 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1379 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1378 = (1'h0);
  reg [(4'hd):(1'h0)] reg1377 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1375 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1374 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1373 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1371 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1370 = (1'h0);
  reg [(4'he):(1'h0)] reg1367 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1366 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1365 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1364 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1362 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1361 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1360 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1359 = (1'h0);
  reg [(3'h6):(1'h0)] reg1358 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1356 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1355 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1354 = (1'h0);
  reg [(2'h2):(1'h0)] reg1353 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1351 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1348 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1347 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1346 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1344 = (1'h0);
  reg [(3'h7):(1'h0)] reg1343 = (1'h0);
  reg [(4'hb):(1'h0)] reg1340 = (1'h0);
  reg [(4'hc):(1'h0)] reg1339 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1338 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1337 = (1'h0);
  reg [(4'hf):(1'h0)] reg1336 = (1'h0);
  reg [(5'h10):(1'h0)] reg1334 = (1'h0);
  reg [(4'hc):(1'h0)] reg1333 = (1'h0);
  reg [(2'h2):(1'h0)] reg1332 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1331 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1328 = (1'h0);
  reg [(4'he):(1'h0)] reg1327 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1326 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1325 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1324 = (1'h0);
  reg [(4'hb):(1'h0)] reg1323 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1322 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1321 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1319 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1318 = (1'h0);
  reg [(3'h7):(1'h0)] reg1317 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1316 = (1'h0);
  reg [(4'hf):(1'h0)] reg1314 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1313 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1312 = (1'h0);
  reg [(4'hb):(1'h0)] reg1311 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1308 = (1'h0);
  reg [(4'hc):(1'h0)] reg1307 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1306 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1305 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1303 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1301 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1300 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1296 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1295 = (1'h0);
  reg [(4'h8):(1'h0)] reg1294 = (1'h0);
  reg [(4'hb):(1'h0)] reg1293 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1292 = (1'h0);
  reg [(4'h9):(1'h0)] reg1291 = (1'h0);
  reg [(3'h6):(1'h0)] reg1289 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1288 = (1'h0);
  reg [(2'h3):(1'h0)] reg1284 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1283 = (1'h0);
  reg [(2'h2):(1'h0)] reg1281 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1279 = (1'h0);
  reg [(4'ha):(1'h0)] reg1278 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1277 = (1'h0);
  reg [(2'h2):(1'h0)] reg1276 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1275 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1274 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1273 = (1'h0);
  reg [(2'h2):(1'h0)] reg1272 = (1'h0);
  reg [(4'h9):(1'h0)] reg1270 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1269 = (1'h0);
  reg [(4'ha):(1'h0)] reg1267 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1266 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1265 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1264 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1262 = (1'h0);
  reg [(3'h4):(1'h0)] reg1261 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1260 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1259 = (1'h0);
  reg [(4'h8):(1'h0)] reg1253 = (1'h0);
  reg [(3'h5):(1'h0)] reg1252 = (1'h0);
  reg [(2'h2):(1'h0)] reg1251 = (1'h0);
  reg [(4'hd):(1'h0)] reg1250 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1248 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1247 = (1'h0);
  reg [(3'h7):(1'h0)] reg1246 = (1'h0);
  reg [(4'hc):(1'h0)] reg1245 = (1'h0);
  reg [(3'h6):(1'h0)] reg1244 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1243 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1242 = (1'h0);
  reg [(2'h3):(1'h0)] reg1241 = (1'h0);
  reg [(2'h3):(1'h0)] reg1240 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1239 = (1'h0);
  reg [(4'h8):(1'h0)] reg1238 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1236 = (1'h0);
  reg [(4'hd):(1'h0)] reg1234 = (1'h0);
  reg [(4'hb):(1'h0)] reg1233 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1232 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1227 = (1'h0);
  reg [(3'h5):(1'h0)] reg1218 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1229 = (1'h0);
  reg [(4'h8):(1'h0)] reg1228 = (1'h0);
  reg [(2'h3):(1'h0)] reg1226 = (1'h0);
  reg [(3'h4):(1'h0)] reg1225 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1224 = (1'h0);
  reg [(3'h6):(1'h0)] reg1223 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1222 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1221 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1220 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1219 = (1'h0);
  reg [(4'hf):(1'h0)] reg1203 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1200 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1199 = (1'h0);
  reg [(3'h5):(1'h0)] reg1182 = (1'h0);
  reg [(2'h2):(1'h0)] reg1211 = (1'h0);
  reg [(4'he):(1'h0)] reg1215 = (1'h0);
  reg [(4'hc):(1'h0)] reg1214 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1213 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1212 = (1'h0);
  reg [(4'hf):(1'h0)] reg1210 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1193 = (1'h0);
  reg [(4'hc):(1'h0)] reg1208 = (1'h0);
  reg [(2'h2):(1'h0)] reg1206 = (1'h0);
  reg [(4'h8):(1'h0)] reg1205 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1204 = (1'h0);
  reg [(2'h2):(1'h0)] reg1202 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1201 = (1'h0);
  reg [(4'hc):(1'h0)] reg1198 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1197 = (1'h0);
  reg [(4'he):(1'h0)] reg1196 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1195 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1194 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1192 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1191 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1190 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1189 = (1'h0);
  reg [(4'ha):(1'h0)] reg1186 = (1'h0);
  reg [(4'hf):(1'h0)] reg1180 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1178 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1188 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1187 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1185 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1184 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1183 = (1'h0);
  reg [(4'h9):(1'h0)] reg1181 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1179 = (1'h0);
  reg [(5'h10):(1'h0)] reg1177 = (1'h0);
  reg [(5'h10):(1'h0)] reg1176 = (1'h0);
  reg [(4'hb):(1'h0)] reg1175 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1174 = (1'h0);
  reg [(5'h10):(1'h0)] reg1173 = (1'h0);
  reg [(2'h3):(1'h0)] reg1172 = (1'h0);
  reg [(2'h3):(1'h0)] reg1171 = (1'h0);
  reg [(3'h5):(1'h0)] reg1170 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1169 = (1'h0);
  reg [(4'hc):(1'h0)] reg1161 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1168 = (1'h0);
  reg [(3'h6):(1'h0)] reg1167 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1166 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1165 = (1'h0);
  reg [(4'h9):(1'h0)] reg1164 = (1'h0);
  reg [(4'hf):(1'h0)] reg1163 = (1'h0);
  reg [(2'h2):(1'h0)] reg1162 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1160 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1636 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1627 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1653 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1644 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1640 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1638 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1637 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1635 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1633 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1626 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1625 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1621 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1620 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1563 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1562 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1557 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1552 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1550 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1547 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1536 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1541 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1538 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1534 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1529 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1617 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1612 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1603 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1602 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1601 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1596 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1591 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1587 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1580 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1575 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1574 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1571 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1565 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1564 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1559 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1558 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1549 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1546 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1545 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1542 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1539 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1530 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1528 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1511 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1505 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1522 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1521 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1517 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1512 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1507 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1514 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1508 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1503 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1497 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1490 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1484 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1475 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1471 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1467 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1466 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1465 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1460 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1455 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1454 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1450 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1449 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1443 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1439 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1437 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1436 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1435 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1433 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1429 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1427 = (1'h0);
  reg [(4'he):(1'h0)] forvar1425 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1420 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1416 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1411 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1410 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1404 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1409 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1402 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1395 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1393 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1392 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1386 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1377 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1376 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1372 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1369 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1368 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1363 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1357 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1352 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1350 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1349 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1343 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1345 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1342 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1341 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1335 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1330 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1329 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1320 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1315 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1310 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1309 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1304 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1302 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1299 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1298 = (1'h0);
  reg [(4'he):(1'h0)] forvar1297 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1290 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1287 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1286 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1285 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1282 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1280 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1271 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1268 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1263 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1258 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1257 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1256 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1249 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1237 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1235 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1231 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1230 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1223 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1227 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1218 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1217 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1216 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1201 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1198 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1197 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1196 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1188 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1177 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1176 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1160 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1210 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1211 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1209 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1207 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1203 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1200 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1199 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1193 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1183 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1179 = (1'h0);
  reg [(4'he):(1'h0)] forvar1175 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1166 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1162 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1186 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1182 = (1'h0);
  reg [(4'he):(1'h0)] forvar1180 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1178 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1170 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1161 = (1'h0);
  assign y = {wire1656,
                 wire1655,
                 wire1464,
                 wire1255,
                 wire1254,
                 wire1159,
                 wire1158,
                 wire1157,
                 wire1156,
                 wire1155,
                 wire1154,
                 reg1633,
                 reg1626,
                 reg1625,
                 reg1654,
                 reg1652,
                 reg1651,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1647,
                 reg1646,
                 reg1645,
                 reg1643,
                 reg1642,
                 reg1641,
                 reg1637,
                 reg1635,
                 reg1640,
                 reg1639,
                 reg1638,
                 reg1636,
                 reg1634,
                 reg1632,
                 reg1631,
                 reg1630,
                 reg1629,
                 reg1628,
                 reg1627,
                 reg1624,
                 reg1623,
                 reg1622,
                 reg1565,
                 reg1564,
                 reg1559,
                 reg1558,
                 reg1549,
                 reg1545,
                 reg1542,
                 reg1539,
                 reg1530,
                 reg1619,
                 reg1618,
                 reg1616,
                 reg1615,
                 reg1614,
                 reg1613,
                 reg1611,
                 reg1610,
                 reg1609,
                 reg1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1602,
                 reg1601,
                 reg1604,
                 reg1603,
                 reg1600,
                 reg1599,
                 reg1598,
                 reg1597,
                 reg1595,
                 reg1594,
                 reg1593,
                 reg1592,
                 reg1590,
                 reg1589,
                 reg1588,
                 reg1586,
                 reg1585,
                 reg1584,
                 reg1583,
                 reg1582,
                 reg1581,
                 reg1579,
                 reg1578,
                 reg1577,
                 reg1576,
                 reg1573,
                 reg1572,
                 reg1570,
                 reg1569,
                 reg1568,
                 reg1567,
                 reg1566,
                 reg1563,
                 reg1562,
                 reg1561,
                 reg1560,
                 reg1557,
                 reg1556,
                 reg1555,
                 reg1554,
                 reg1553,
                 reg1552,
                 reg1551,
                 reg1550,
                 reg1548,
                 reg1547,
                 reg1544,
                 reg1543,
                 reg1541,
                 reg1540,
                 reg1538,
                 reg1537,
                 reg1536,
                 reg1535,
                 reg1534,
                 reg1533,
                 reg1532,
                 reg1531,
                 reg1529,
                 reg1503,
                 reg1527,
                 reg1526,
                 reg1525,
                 reg1524,
                 reg1523,
                 reg1520,
                 reg1519,
                 reg1518,
                 reg1514,
                 reg1508,
                 reg1517,
                 reg1516,
                 reg1515,
                 reg1513,
                 reg1512,
                 reg1511,
                 reg1510,
                 reg1509,
                 reg1507,
                 reg1506,
                 reg1505,
                 reg1504,
                 reg1502,
                 reg1501,
                 reg1500,
                 reg1499,
                 reg1498,
                 reg1496,
                 reg1495,
                 reg1494,
                 reg1493,
                 reg1490,
                 reg1492,
                 reg1491,
                 reg1489,
                 reg1488,
                 reg1487,
                 reg1486,
                 reg1485,
                 reg1483,
                 reg1482,
                 reg1481,
                 reg1480,
                 reg1479,
                 reg1478,
                 reg1477,
                 reg1476,
                 reg1474,
                 reg1473,
                 reg1472,
                 reg1470,
                 reg1469,
                 reg1466,
                 reg1468,
                 reg1467,
                 reg1463,
                 reg1462,
                 reg1461,
                 reg1459,
                 reg1458,
                 reg1457,
                 reg1456,
                 reg1453,
                 reg1452,
                 reg1451,
                 reg1448,
                 reg1447,
                 reg1446,
                 reg1445,
                 reg1444,
                 reg1442,
                 reg1441,
                 reg1440,
                 reg1438,
                 reg1425,
                 reg1434,
                 reg1432,
                 reg1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1426,
                 reg1424,
                 reg1423,
                 reg1422,
                 reg1421,
                 reg1419,
                 reg1418,
                 reg1417,
                 reg1415,
                 reg1414,
                 reg1413,
                 reg1409,
                 reg1412,
                 reg1411,
                 reg1410,
                 reg1408,
                 reg1407,
                 reg1406,
                 reg1405,
                 reg1404,
                 reg1403,
                 reg1401,
                 reg1400,
                 reg1399,
                 reg1398,
                 reg1397,
                 reg1396,
                 reg1394,
                 reg1386,
                 reg1391,
                 reg1390,
                 reg1389,
                 reg1388,
                 reg1387,
                 reg1385,
                 reg1384,
                 reg1383,
                 reg1382,
                 reg1381,
                 reg1380,
                 reg1379,
                 reg1378,
                 reg1377,
                 reg1375,
                 reg1374,
                 reg1373,
                 reg1371,
                 reg1370,
                 reg1367,
                 reg1366,
                 reg1365,
                 reg1364,
                 reg1362,
                 reg1361,
                 reg1360,
                 reg1359,
                 reg1358,
                 reg1356,
                 reg1355,
                 reg1354,
                 reg1353,
                 reg1351,
                 reg1348,
                 reg1347,
                 reg1346,
                 reg1344,
                 reg1343,
                 reg1340,
                 reg1339,
                 reg1338,
                 reg1337,
                 reg1336,
                 reg1334,
                 reg1333,
                 reg1332,
                 reg1331,
                 reg1328,
                 reg1327,
                 reg1326,
                 reg1325,
                 reg1324,
                 reg1323,
                 reg1322,
                 reg1321,
                 reg1319,
                 reg1318,
                 reg1317,
                 reg1316,
                 reg1314,
                 reg1313,
                 reg1312,
                 reg1311,
                 reg1308,
                 reg1307,
                 reg1306,
                 reg1305,
                 reg1303,
                 reg1301,
                 reg1300,
                 reg1296,
                 reg1295,
                 reg1294,
                 reg1293,
                 reg1292,
                 reg1291,
                 reg1289,
                 reg1288,
                 reg1284,
                 reg1283,
                 reg1281,
                 reg1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 reg1275,
                 reg1274,
                 reg1273,
                 reg1272,
                 reg1270,
                 reg1269,
                 reg1267,
                 reg1266,
                 reg1265,
                 reg1264,
                 reg1262,
                 reg1261,
                 reg1260,
                 reg1259,
                 reg1253,
                 reg1252,
                 reg1251,
                 reg1250,
                 reg1248,
                 reg1247,
                 reg1246,
                 reg1245,
                 reg1244,
                 reg1243,
                 reg1242,
                 reg1241,
                 reg1240,
                 reg1239,
                 reg1238,
                 reg1236,
                 reg1234,
                 reg1233,
                 reg1232,
                 reg1227,
                 reg1218,
                 reg1229,
                 reg1228,
                 reg1226,
                 reg1225,
                 reg1224,
                 reg1223,
                 reg1222,
                 reg1221,
                 reg1220,
                 reg1219,
                 reg1203,
                 reg1200,
                 reg1199,
                 reg1182,
                 reg1211,
                 reg1215,
                 reg1214,
                 reg1213,
                 reg1212,
                 reg1210,
                 reg1193,
                 reg1208,
                 reg1206,
                 reg1205,
                 reg1204,
                 reg1202,
                 reg1201,
                 reg1198,
                 reg1197,
                 reg1196,
                 reg1195,
                 reg1194,
                 reg1192,
                 reg1191,
                 reg1190,
                 reg1189,
                 reg1186,
                 reg1180,
                 reg1178,
                 reg1188,
                 reg1187,
                 reg1185,
                 reg1184,
                 reg1183,
                 reg1181,
                 reg1179,
                 reg1177,
                 reg1176,
                 reg1175,
                 reg1174,
                 reg1173,
                 reg1172,
                 reg1171,
                 reg1170,
                 reg1169,
                 reg1161,
                 reg1168,
                 reg1167,
                 reg1166,
                 reg1165,
                 reg1164,
                 reg1163,
                 reg1162,
                 reg1160,
                 forvar1636,
                 forvar1627,
                 forvar1653,
                 forvar1644,
                 forvar1640,
                 forvar1638,
                 forvar1637,
                 forvar1635,
                 forvar1633,
                 forvar1626,
                 forvar1625,
                 forvar1621,
                 forvar1620,
                 forvar1563,
                 forvar1562,
                 forvar1557,
                 forvar1552,
                 forvar1550,
                 forvar1547,
                 forvar1536,
                 forvar1541,
                 forvar1538,
                 forvar1534,
                 forvar1529,
                 forvar1617,
                 forvar1612,
                 forvar1603,
                 forvar1602,
                 forvar1601,
                 forvar1596,
                 forvar1591,
                 forvar1587,
                 forvar1580,
                 forvar1575,
                 forvar1574,
                 forvar1571,
                 forvar1565,
                 forvar1564,
                 forvar1559,
                 forvar1558,
                 forvar1549,
                 forvar1546,
                 forvar1545,
                 forvar1542,
                 forvar1539,
                 forvar1530,
                 forvar1528,
                 forvar1511,
                 forvar1505,
                 forvar1522,
                 forvar1521,
                 forvar1517,
                 forvar1512,
                 forvar1507,
                 forvar1514,
                 forvar1508,
                 forvar1503,
                 forvar1497,
                 forvar1490,
                 forvar1484,
                 forvar1475,
                 forvar1471,
                 forvar1467,
                 forvar1466,
                 forvar1465,
                 forvar1460,
                 forvar1455,
                 forvar1454,
                 forvar1450,
                 forvar1449,
                 forvar1443,
                 forvar1439,
                 forvar1437,
                 forvar1436,
                 forvar1435,
                 forvar1433,
                 forvar1429,
                 forvar1427,
                 forvar1425,
                 forvar1420,
                 forvar1416,
                 forvar1411,
                 forvar1410,
                 forvar1404,
                 forvar1409,
                 forvar1402,
                 forvar1395,
                 forvar1393,
                 forvar1392,
                 forvar1386,
                 forvar1377,
                 forvar1376,
                 forvar1372,
                 forvar1369,
                 forvar1368,
                 forvar1363,
                 forvar1357,
                 forvar1352,
                 forvar1350,
                 forvar1349,
                 forvar1343,
                 forvar1345,
                 forvar1342,
                 forvar1341,
                 forvar1335,
                 forvar1330,
                 forvar1329,
                 forvar1320,
                 forvar1315,
                 forvar1310,
                 forvar1309,
                 forvar1304,
                 forvar1302,
                 forvar1299,
                 forvar1298,
                 forvar1297,
                 forvar1290,
                 forvar1287,
                 forvar1286,
                 forvar1285,
                 forvar1282,
                 forvar1280,
                 forvar1271,
                 forvar1268,
                 forvar1263,
                 forvar1258,
                 forvar1257,
                 forvar1256,
                 forvar1249,
                 forvar1237,
                 forvar1235,
                 forvar1231,
                 forvar1230,
                 forvar1223,
                 forvar1227,
                 forvar1218,
                 forvar1217,
                 forvar1216,
                 forvar1201,
                 forvar1198,
                 forvar1197,
                 forvar1196,
                 forvar1188,
                 forvar1177,
                 forvar1176,
                 forvar1160,
                 forvar1210,
                 forvar1211,
                 forvar1209,
                 forvar1207,
                 forvar1203,
                 forvar1200,
                 forvar1199,
                 forvar1193,
                 forvar1183,
                 forvar1179,
                 forvar1175,
                 forvar1166,
                 forvar1162,
                 forvar1186,
                 forvar1182,
                 forvar1180,
                 forvar1178,
                 forvar1170,
                 forvar1161,
                 (1'h0)};
  assign wire1154 = {{$unsigned(wire1149[(1'h1):(1'h1)])}};
  assign wire1155 = wire1154[(1'h1):(1'h0)];
  assign wire1156 = $signed((8'h9e));
  assign wire1157 = ($unsigned({(wire1152 ? wire1151 : wire1153)}) ?
                        (($signed((8'ha2)) ?
                            $unsigned(wire1149) : wire1152[(4'h8):(3'h7)]) > (-((8'ha9) & wire1156))) : ((~&(wire1155 <= wire1150)) * wire1150));
  assign wire1158 = wire1151;
  assign wire1159 = $signed(({(wire1151 || wire1151)} != $signed(wire1157[(3'h5):(3'h4)])));
  always
    @(posedge clk) begin
      if ((8'hb2))
        begin
          reg1160 <= (|wire1150[(2'h3):(1'h0)]);
          if ($unsigned((~|$signed(wire1159))))
            begin
              if ((((!$unsigned(wire1154)) < {wire1155[(4'h9):(4'h9)]}) <<< ($signed({wire1156}) & $unsigned(wire1149))))
                begin
                  for (forvar1161 = (1'h0); (forvar1161 < (2'h2)); forvar1161 = (forvar1161 + (1'h1)))
                    begin
                      reg1162 <= (&forvar1161[(1'h0):(1'h0)]);
                      reg1163 <= (-$signed((((8'ha5) && (8'ha5)) & (wire1149 ?
                          (8'hba) : reg1160))));
                      reg1164 <= wire1153;
                    end
                  if ((wire1149 ?
                      wire1154[(4'h9):(2'h3)] : $signed($signed((^~reg1164)))))
                    begin
                      reg1165 <= ($signed($unsigned(wire1154)) ^~ $signed($unsigned(reg1160)));
                      reg1166 <= ((^~reg1160[(4'h8):(3'h6)]) || $unsigned((+$unsigned(wire1153))));
                    end
                  else
                    begin
                      reg1165 <= {($unsigned(wire1154[(1'h0):(1'h0)]) ?
                              wire1158[(3'h4):(2'h2)] : (^(wire1159 ?
                                  wire1156 : wire1149)))};
                      reg1166 <= $unsigned(($signed($unsigned(reg1160)) ?
                          (forvar1161 ?
                              reg1162[(1'h1):(1'h1)] : $unsigned((8'hb3))) : {(wire1151 << wire1155)}));
                      reg1167 <= (8'haf);
                    end
                  reg1168 <= reg1163[(4'hf):(4'hb)];
                end
              else
                begin
                  reg1161 <= (8'hb0);
                end
              reg1169 <= $signed($signed((~&(|wire1152))));
              if ((|$unsigned(wire1156[(4'h9):(1'h1)])))
                begin
                  if (reg1169)
                    begin
                      reg1170 <= ((wire1156[(3'h4):(2'h3)] && ((reg1168 >= (8'hac)) >>> $unsigned(wire1155))) ?
                          wire1159 : wire1157);
                    end
                  else
                    begin
                      reg1170 <= $unsigned((&$unsigned(((8'ha9) * wire1158))));
                      reg1171 <= ((wire1155[(3'h6):(3'h5)] ?
                          {(reg1160 ?
                                  wire1150 : wire1151)} : reg1163[(3'h6):(1'h0)]) < (^(^~$unsigned(wire1158))));
                    end
                  if (reg1161[(1'h1):(1'h1)])
                    begin
                      reg1172 <= ($signed($unsigned(((8'ha2) & (8'hba)))) << wire1153);
                      reg1173 <= $unsigned($signed($signed({wire1154})));
                      reg1174 <= $unsigned((reg1163 - $unsigned((reg1165 > (8'hb0)))));
                    end
                  else
                    begin
                      reg1172 <= $unsigned((8'ha7));
                      reg1173 <= ((wire1158[(3'h5):(2'h2)] < ($signed(reg1166) & reg1173[(4'h8):(4'h8)])) - $unsigned(((8'hb6) ?
                          $unsigned((8'hb8)) : reg1173)));
                      reg1174 <= ({($unsigned((8'hb5)) == (|wire1159))} ?
                          reg1165 : $signed(($unsigned(reg1169) ?
                              (~reg1164) : (reg1163 ? reg1171 : reg1166))));
                      reg1175 <= (~&$unsigned(({reg1169} ?
                          $signed(wire1156) : (wire1155 ? (8'hac) : reg1172))));
                    end
                end
              else
                begin
                  for (forvar1170 = (1'h0); (forvar1170 < (1'h0)); forvar1170 = (forvar1170 + (1'h1)))
                    begin
                      reg1171 <= {($signed($unsigned(reg1170)) - (8'ha7))};
                      reg1172 <= wire1154;
                      reg1173 <= (~^reg1165[(2'h3):(1'h1)]);
                    end
                  if ($signed(($unsigned($unsigned((8'ha9))) ?
                      (~^(reg1169 ?
                          wire1157 : (8'hb1))) : $unsigned(((8'hae) || wire1150)))))
                    begin
                      reg1174 <= reg1161;
                      reg1175 <= (~^(((wire1151 ? reg1171 : reg1160) ?
                          reg1173[(3'h5):(1'h1)] : reg1169) - ($signed(reg1169) * wire1158)));
                      reg1176 <= {(({reg1163} == (wire1159 ?
                              reg1173 : (8'hb5))) ~^ ($signed(wire1152) ?
                              $signed(reg1161) : reg1169))};
                      reg1177 <= (|$signed((+reg1162[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg1174 <= wire1154;
                      reg1175 <= $signed(forvar1170);
                      reg1176 <= reg1168;
                    end
                end
              for (forvar1178 = (1'h0); (forvar1178 < (1'h0)); forvar1178 = (forvar1178 + (1'h1)))
                begin
                  if (reg1166[(2'h2):(2'h2)])
                    begin
                      reg1179 <= (reg1168[(4'h8):(1'h1)] >= reg1174[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1179 <= $unsigned($unsigned((-wire1154)));
                    end
                  for (forvar1180 = (1'h0); (forvar1180 < (1'h1)); forvar1180 = (forvar1180 + (1'h1)))
                    begin
                      reg1181 <= reg1163[(4'hd):(3'h7)];
                    end
                  for (forvar1182 = (1'h0); (forvar1182 < (2'h3)); forvar1182 = (forvar1182 + (1'h1)))
                    begin
                      reg1183 <= (~&(reg1170[(1'h1):(1'h0)] ?
                          {(wire1151 | reg1162)} : (forvar1170[(2'h2):(2'h2)] > $unsigned(reg1170))));
                      reg1184 <= wire1156;
                      reg1185 <= $signed({($unsigned((8'hb6)) && (8'hb2))});
                    end
                  for (forvar1186 = (1'h0); (forvar1186 < (1'h1)); forvar1186 = (forvar1186 + (1'h1)))
                    begin
                      reg1187 <= reg1172[(1'h0):(1'h0)];
                      reg1188 <= ($signed($unsigned($unsigned(reg1167))) ^~ wire1153[(2'h3):(2'h3)]);
                    end
                end
            end
          else
            begin
              for (forvar1161 = (1'h0); (forvar1161 < (2'h2)); forvar1161 = (forvar1161 + (1'h1)))
                begin
                  for (forvar1162 = (1'h0); (forvar1162 < (1'h1)); forvar1162 = (forvar1162 + (1'h1)))
                    begin
                      reg1163 <= ($signed(wire1152) - reg1176[(3'h5):(1'h0)]);
                      reg1164 <= (^(8'h9d));
                      reg1165 <= ($signed((reg1172[(1'h0):(1'h0)] << (+(8'ha7)))) ~^ $signed((|(reg1165 ?
                          wire1154 : reg1160))));
                    end
                  for (forvar1166 = (1'h0); (forvar1166 < (2'h2)); forvar1166 = (forvar1166 + (1'h1)))
                    begin
                      reg1167 <= reg1162[(1'h1):(1'h1)];
                    end
                  if ({{$signed((reg1183 != reg1162))}})
                    begin
                      reg1168 <= $unsigned(reg1162);
                    end
                  else
                    begin
                      reg1168 <= $unsigned((((^~wire1153) ?
                          $signed(reg1163) : (reg1183 ?
                              (8'hab) : wire1156)) | (^~((8'h9f) ~^ (8'ha5)))));
                    end
                  reg1169 <= (forvar1161[(2'h2):(1'h0)] ?
                      reg1168[(4'h8):(3'h5)] : (8'hb3));
                end
              reg1170 <= (reg1185[(3'h4):(3'h4)] >= reg1174);
              if ((|(($unsigned((8'h9c)) ?
                      $unsigned(wire1156) : $unsigned(reg1162)) ?
                  ({reg1162} ?
                      reg1163[(2'h3):(1'h1)] : $unsigned(forvar1182)) : reg1171[(1'h0):(1'h0)])))
                begin
                  if (reg1165)
                    begin
                      reg1171 <= ($unsigned((~$signed((8'hb4)))) ?
                          reg1164 : reg1174[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg1171 <= $unsigned(reg1187);
                    end
                end
              else
                begin
                  if (wire1155)
                    begin
                      reg1171 <= $signed(($unsigned((8'hae)) ?
                          wire1155 : reg1166[(1'h1):(1'h1)]));
                      reg1172 <= {((|(-reg1175)) < wire1154)};
                      reg1173 <= $signed(wire1157);
                      reg1174 <= (8'h9c);
                    end
                  else
                    begin
                      reg1171 <= $unsigned(reg1185);
                    end
                  for (forvar1175 = (1'h0); (forvar1175 < (2'h3)); forvar1175 = (forvar1175 + (1'h1)))
                    begin
                      reg1176 <= (((8'ha2) != (~&(forvar1166 ?
                          (8'had) : wire1154))) * ($signed($unsigned(reg1172)) ?
                          (!(+reg1164)) : ((!(8'hb3)) ?
                              (|forvar1175) : (forvar1175 ?
                                  (8'hb6) : forvar1162))));
                      reg1177 <= ($unsigned($unsigned(reg1162)) ?
                          wire1151[(2'h2):(2'h2)] : (^wire1151));
                      reg1178 <= ($signed(reg1177) ?
                          ((~&((8'hb8) + forvar1180)) && wire1159) : {forvar1186[(1'h1):(1'h1)]});
                    end
                  for (forvar1179 = (1'h0); (forvar1179 < (1'h1)); forvar1179 = (forvar1179 + (1'h1)))
                    begin
                      reg1180 <= (|($signed((forvar1166 ? reg1163 : reg1167)) ?
                          {reg1179[(4'h9):(4'h8)]} : forvar1178));
                      reg1181 <= forvar1166;
                    end
                end
              for (forvar1182 = (1'h0); (forvar1182 < (2'h2)); forvar1182 = (forvar1182 + (1'h1)))
                begin
                  for (forvar1183 = (1'h0); (forvar1183 < (1'h0)); forvar1183 = (forvar1183 + (1'h1)))
                    begin
                      reg1184 <= ($unsigned($signed(wire1152)) << (8'ha7));
                      reg1185 <= ($unsigned((~$signed(wire1150))) << reg1183[(1'h1):(1'h1)]);
                    end
                  if ($signed(reg1181))
                    begin
                      reg1186 <= (+$signed(wire1152[(2'h3):(2'h2)]));
                      reg1187 <= reg1181[(3'h5):(3'h4)];
                      reg1188 <= {$signed($signed((reg1176 ^~ wire1153)))};
                      reg1189 <= (-$unsigned((~|((8'h9f) + forvar1170))));
                    end
                  else
                    begin
                      reg1186 <= $signed({wire1152[(4'hc):(1'h0)]});
                      reg1187 <= forvar1170;
                    end
                  if (reg1177[(3'h4):(2'h3)])
                    begin
                      reg1190 <= ((forvar1170 ~^ (|wire1151[(2'h3):(1'h0)])) * $signed($signed((~reg1188))));
                      reg1191 <= (8'haf);
                      reg1192 <= (~&$unsigned($signed((reg1163 + reg1184))));
                    end
                  else
                    begin
                      reg1190 <= $unsigned(($signed({wire1151}) >> reg1170[(1'h0):(1'h0)]));
                      reg1191 <= $signed((~|reg1186));
                      reg1192 <= reg1162;
                    end
                end
            end
          if (reg1174[(1'h0):(1'h0)])
            begin
              for (forvar1193 = (1'h0); (forvar1193 < (2'h3)); forvar1193 = (forvar1193 + (1'h1)))
                begin
                  if ((+$signed(wire1157)))
                    begin
                      reg1194 <= (($signed((wire1149 >> forvar1162)) ^ (8'hb8)) == {$unsigned((wire1153 ?
                              reg1172 : wire1156))});
                      reg1195 <= reg1171;
                    end
                  else
                    begin
                      reg1194 <= {$signed(reg1194)};
                      reg1195 <= reg1175[(1'h0):(1'h0)];
                      reg1196 <= (($unsigned((reg1163 <= reg1189)) >= reg1185) ?
                          reg1175[(2'h2):(1'h1)] : (|(reg1165 <= reg1164)));
                      reg1197 <= ($signed(($unsigned((8'ha6)) * ((8'haa) && reg1162))) ?
                          ($unsigned((~|reg1174)) && (reg1173 << reg1181[(4'h9):(3'h7)])) : $signed({$unsigned(reg1185)}));
                    end
                end
              reg1198 <= ($signed({reg1180[(4'hc):(3'h6)]}) ?
                  reg1168[(2'h2):(1'h0)] : reg1196);
              for (forvar1199 = (1'h0); (forvar1199 < (2'h2)); forvar1199 = (forvar1199 + (1'h1)))
                begin
                  for (forvar1200 = (1'h0); (forvar1200 < (2'h3)); forvar1200 = (forvar1200 + (1'h1)))
                    begin
                      reg1201 <= (~|$signed((8'hab)));
                      reg1202 <= $unsigned(((~^forvar1193) << (8'ha1)));
                    end
                  for (forvar1203 = (1'h0); (forvar1203 < (1'h0)); forvar1203 = (forvar1203 + (1'h1)))
                    begin
                      reg1204 <= (reg1180 ? wire1156 : wire1159);
                      reg1205 <= (reg1170[(1'h1):(1'h0)] ?
                          $unsigned(forvar1200[(4'hd):(4'ha)]) : {(-(~^reg1174))});
                      reg1206 <= wire1149;
                    end
                end
              for (forvar1207 = (1'h0); (forvar1207 < (1'h1)); forvar1207 = (forvar1207 + (1'h1)))
                begin
                  if (reg1201)
                    begin
                      reg1208 <= (((reg1172[(1'h1):(1'h1)] & $signed(reg1174)) | {(reg1178 - (8'hac))}) <<< ((~&$signed(wire1155)) ?
                          (^(reg1181 ?
                              forvar1162 : wire1157)) : $unsigned({forvar1161})));
                    end
                  else
                    begin
                      reg1208 <= reg1180[(3'h6):(1'h1)];
                    end
                end
            end
          else
            begin
              reg1193 <= {(8'hb3)};
            end
          for (forvar1209 = (1'h0); (forvar1209 < (1'h1)); forvar1209 = (forvar1209 + (1'h1)))
            begin
              if ((($signed(reg1189[(4'hd):(4'hb)]) && reg1176[(4'hd):(4'ha)]) <<< (((-reg1170) ^~ $unsigned(forvar1186)) ?
                  reg1179 : (8'hb6))))
                begin
                  reg1210 <= (8'h9e);
                  for (forvar1211 = (1'h0); (forvar1211 < (2'h2)); forvar1211 = (forvar1211 + (1'h1)))
                    begin
                      reg1212 <= reg1187[(1'h0):(1'h0)];
                      reg1213 <= $signed(reg1162[(1'h1):(1'h1)]);
                      reg1214 <= (wire1157[(3'h5):(3'h4)] ?
                          ({{wire1152}} > $unsigned($unsigned(forvar1203))) : wire1151);
                      reg1215 <= $unsigned($unsigned($signed(wire1151)));
                    end
                end
              else
                begin
                  for (forvar1210 = (1'h0); (forvar1210 < (1'h1)); forvar1210 = (forvar1210 + (1'h1)))
                    begin
                      reg1211 <= ((({forvar1193} <= $signed(reg1185)) ?
                              reg1173[(4'hd):(4'hc)] : (wire1152[(3'h4):(1'h0)] ?
                                  ((8'hba) ?
                                      reg1176 : (8'hab)) : (wire1151 ^ forvar1161))) ?
                          ($unsigned((reg1188 ?
                              forvar1210 : forvar1210)) < (forvar1203[(1'h1):(1'h0)] ?
                              reg1170 : $signed(reg1176))) : reg1189[(2'h2):(1'h0)]);
                      reg1212 <= ({(+(-reg1189))} ?
                          reg1177[(1'h0):(1'h0)] : ($signed((forvar1175 >>> reg1213)) ^~ forvar1211[(1'h1):(1'h0)]));
                    end
                end
            end
        end
      else
        begin
          if ((8'ha3))
            begin
              reg1160 <= (^{wire1152[(3'h7):(3'h6)]});
            end
          else
            begin
              if ((^$signed((forvar1211[(4'h9):(3'h6)] >> (forvar1186 ?
                  (8'h9c) : (8'ha7))))))
                begin
                  for (forvar1160 = (1'h0); (forvar1160 < (2'h3)); forvar1160 = (forvar1160 + (1'h1)))
                    begin
                      reg1161 <= (8'hb5);
                    end
                end
              else
                begin
                  if (forvar1211[(4'hb):(4'h8)])
                    begin
                      reg1160 <= $signed(forvar1199[(2'h2):(1'h0)]);
                      reg1161 <= (8'hae);
                      reg1162 <= $unsigned((8'ha4));
                      reg1163 <= ($signed($unsigned(wire1159[(3'h7):(2'h2)])) ?
                          (^~{(wire1150 ? reg1179 : wire1151)}) : (~|(8'hb3)));
                    end
                  else
                    begin
                      reg1160 <= wire1155[(4'h9):(3'h4)];
                    end
                  if ((8'haa))
                    begin
                      reg1164 <= $signed($unsigned({$unsigned(reg1169)}));
                      reg1165 <= (+reg1190);
                      reg1166 <= forvar1203;
                      reg1167 <= $unsigned($unsigned($signed({forvar1161})));
                    end
                  else
                    begin
                      reg1164 <= $signed((reg1161 ^~ $signed($signed(reg1171))));
                      reg1165 <= ({({reg1196} ?
                                  {(8'ha5)} : reg1175[(4'h8):(1'h0)])} ?
                          $signed(reg1172[(2'h3):(1'h1)]) : reg1211);
                      reg1166 <= (^~({$unsigned(reg1187)} ?
                          wire1158[(4'h8):(2'h3)] : $unsigned(reg1163)));
                      reg1167 <= ((reg1166[(1'h0):(1'h0)] <<< (~^$unsigned((8'ha4)))) ?
                          (^~((+reg1190) ^ (+(8'ha6)))) : $unsigned(((reg1178 ?
                              reg1202 : wire1158) << $unsigned(wire1156))));
                    end
                  if ((($unsigned(forvar1210) | wire1153) ?
                      $signed((forvar1209 ?
                          ((8'ha2) ? reg1205 : reg1188) : reg1161)) : wire1152))
                    begin
                      reg1168 <= ((~&$unsigned($unsigned(reg1193))) <= reg1162[(1'h1):(1'h1)]);
                      reg1169 <= ($signed((^reg1172)) ?
                          (reg1176[(3'h6):(2'h3)] - $unsigned((reg1180 || reg1196))) : ((-(^(8'hb6))) != ($unsigned(forvar1209) || {forvar1160})));
                      reg1170 <= (~|$unsigned((reg1169 ?
                          (reg1168 != reg1214) : $unsigned(reg1190))));
                      reg1171 <= reg1162[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg1168 <= (~^{$unsigned((reg1213 ~^ (8'hb7)))});
                    end
                  if ((|{(((8'haa) ?
                          reg1172 : reg1170) <= forvar1170[(2'h2):(1'h0)])}))
                    begin
                      reg1172 <= (forvar1161[(1'h1):(1'h0)] ^ (($signed(reg1193) - {reg1188}) ?
                          (reg1161[(3'h4):(2'h2)] >= $unsigned(reg1163)) : reg1198));
                      reg1173 <= $unsigned((^({forvar1170} == (reg1178 ?
                          reg1162 : reg1178))));
                      reg1174 <= {$signed($unsigned((~^reg1192)))};
                      reg1175 <= $signed({$signed((&(8'ha5)))});
                    end
                  else
                    begin
                      reg1172 <= (reg1169[(3'h5):(1'h0)] << $unsigned({$unsigned(reg1188)}));
                      reg1173 <= $unsigned({(8'h9e)});
                      reg1174 <= (((|$unsigned(reg1194)) ?
                              reg1188[(2'h3):(1'h0)] : (wire1150 ?
                                  $signed(reg1212) : (-wire1156))) ?
                          ($signed($signed(reg1191)) ?
                              reg1176[(4'ha):(3'h7)] : (reg1193 ?
                                  $signed(wire1157) : $unsigned(reg1179))) : $unsigned({((8'ha9) ?
                                  (8'hb4) : reg1189)}));
                    end
                end
              for (forvar1176 = (1'h0); (forvar1176 < (1'h0)); forvar1176 = (forvar1176 + (1'h1)))
                begin
                  for (forvar1177 = (1'h0); (forvar1177 < (2'h2)); forvar1177 = (forvar1177 + (1'h1)))
                    begin
                      reg1178 <= (((!$unsigned(reg1179)) || (reg1172 <<< (^reg1179))) < (~($unsigned(forvar1182) ?
                          (~|wire1158) : {wire1158})));
                      reg1179 <= reg1181[(3'h7):(2'h2)];
                    end
                  if ($signed((^(&(wire1157 - wire1149)))))
                    begin
                      reg1180 <= wire1153;
                      reg1181 <= (wire1156[(3'h6):(3'h5)] >= (($unsigned(reg1205) ?
                              $unsigned((8'ha9)) : $signed(wire1157)) ?
                          forvar1175[(3'h6):(1'h1)] : (~|$unsigned(reg1188))));
                      reg1182 <= $signed(((8'ha7) && {reg1173}));
                      reg1183 <= {(8'ha8)};
                    end
                  else
                    begin
                      reg1180 <= (8'hb3);
                      reg1181 <= (((8'ha2) ^ forvar1207[(1'h0):(1'h0)]) ?
                          $signed($unsigned(wire1155)) : forvar1200);
                      reg1182 <= (-$unsigned((reg1178[(1'h1):(1'h0)] ?
                          (&wire1156) : (!reg1168))));
                    end
                  if ($unsigned(((forvar1210[(3'h6):(1'h1)] ?
                          $unsigned(forvar1193) : (~&forvar1160)) ?
                      {{reg1160}} : $signed((reg1166 - forvar1161)))))
                    begin
                      reg1184 <= (8'hba);
                    end
                  else
                    begin
                      reg1184 <= $unsigned(($signed((&reg1201)) | ({reg1201} ?
                          (forvar1209 != wire1149) : $unsigned(reg1205))));
                      reg1185 <= ({(-(wire1151 ?
                              reg1205 : reg1186))} >= reg1173);
                      reg1186 <= $unsigned((8'h9e));
                      reg1187 <= (reg1202[(1'h0):(1'h0)] ?
                          $unsigned(($signed(reg1177) ?
                              forvar1166 : (-reg1202))) : {wire1149});
                    end
                  for (forvar1188 = (1'h0); (forvar1188 < (2'h3)); forvar1188 = (forvar1188 + (1'h1)))
                    begin
                      reg1189 <= ((reg1213[(2'h2):(1'h1)] ?
                          $unsigned({reg1160}) : ((forvar1188 ?
                              forvar1207 : wire1154) ^ $unsigned(reg1202))) != $signed(forvar1166[(1'h0):(1'h0)]));
                      reg1190 <= (|$signed(((&(8'hae)) + (~&reg1181))));
                      reg1191 <= forvar1176;
                      reg1192 <= $unsigned(($signed((|reg1193)) ?
                          (reg1168[(3'h6):(3'h5)] ?
                              (reg1214 ?
                                  reg1188 : forvar1162) : reg1192) : forvar1193[(1'h0):(1'h0)]));
                    end
                end
              reg1193 <= ((&reg1185) << (~reg1185[(1'h0):(1'h0)]));
              reg1194 <= wire1158;
            end
          reg1195 <= {(($signed(wire1158) + (~reg1215)) ?
                  $signed(forvar1176[(2'h2):(1'h1)]) : forvar1200)};
          for (forvar1196 = (1'h0); (forvar1196 < (2'h2)); forvar1196 = (forvar1196 + (1'h1)))
            begin
              for (forvar1197 = (1'h0); (forvar1197 < (2'h3)); forvar1197 = (forvar1197 + (1'h1)))
                begin
                  for (forvar1198 = (1'h0); (forvar1198 < (2'h2)); forvar1198 = (forvar1198 + (1'h1)))
                    begin
                      reg1199 <= ({({reg1161} | reg1161)} ~^ {$signed((~|wire1156))});
                      reg1200 <= reg1205[(1'h1):(1'h1)];
                    end
                end
              for (forvar1201 = (1'h0); (forvar1201 < (2'h3)); forvar1201 = (forvar1201 + (1'h1)))
                begin
                  reg1202 <= $unsigned((~$unsigned(((8'hb6) ?
                      wire1155 : forvar1183))));
                end
              reg1203 <= forvar1179[(4'h8):(1'h0)];
            end
          reg1204 <= reg1202;
        end
      for (forvar1216 = (1'h0); (forvar1216 < (2'h2)); forvar1216 = (forvar1216 + (1'h1)))
        begin
          for (forvar1217 = (1'h0); (forvar1217 < (1'h0)); forvar1217 = (forvar1217 + (1'h1)))
            begin
              if ((^~reg1173[(3'h5):(1'h1)]))
                begin
                  for (forvar1218 = (1'h0); (forvar1218 < (1'h1)); forvar1218 = (forvar1218 + (1'h1)))
                    begin
                      reg1219 <= ((~{forvar1176}) & $unsigned(($unsigned(forvar1162) ?
                          (reg1212 ?
                              forvar1200 : reg1169) : reg1171[(2'h2):(1'h0)])));
                      reg1220 <= (-(($signed(forvar1186) && reg1203) ?
                          forvar1170 : (+(^forvar1177))));
                    end
                  if ((-$signed(($unsigned(reg1165) | (forvar1199 ?
                      (8'hb7) : forvar1176)))))
                    begin
                      reg1221 <= (reg1176[(4'hc):(4'h8)] << (reg1162 != forvar1197[(3'h5):(3'h5)]));
                      reg1222 <= $signed((8'hab));
                      reg1223 <= (forvar1210 ? reg1176 : {(8'ha4)});
                      reg1224 <= (forvar1180[(3'h6):(2'h3)] ?
                          (reg1201 ?
                              (~|$unsigned(reg1189)) : reg1194) : (reg1179 | reg1203));
                    end
                  else
                    begin
                      reg1221 <= ((!$signed((~&reg1192))) * reg1195[(1'h1):(1'h1)]);
                      reg1222 <= ($unsigned(reg1187[(2'h3):(1'h1)]) ?
                          forvar1177 : (reg1172[(1'h1):(1'h1)] ?
                              reg1171[(2'h3):(1'h1)] : $signed($signed(reg1178))));
                      reg1223 <= $unsigned((reg1200 * reg1203));
                      reg1224 <= reg1169;
                    end
                  if (($unsigned((^~$unsigned(reg1187))) ?
                      reg1172[(2'h2):(1'h1)] : $unsigned($signed((&reg1170)))))
                    begin
                      reg1225 <= ((((reg1222 || reg1160) ?
                          wire1154[(4'ha):(2'h3)] : reg1222[(2'h3):(2'h2)]) >= $signed(reg1194)) | (|forvar1211[(4'hf):(1'h1)]));
                    end
                  else
                    begin
                      reg1225 <= (~^$unsigned((^~reg1170[(2'h3):(1'h0)])));
                      reg1226 <= forvar1211[(4'hd):(4'hd)];
                    end
                  for (forvar1227 = (1'h0); (forvar1227 < (1'h1)); forvar1227 = (forvar1227 + (1'h1)))
                    begin
                      reg1228 <= $unsigned(reg1208);
                      reg1229 <= $unsigned(forvar1211);
                    end
                end
              else
                begin
                  if (forvar1176)
                    begin
                      reg1218 <= ($unsigned((~(&wire1154))) <<< $unsigned({forvar1201[(2'h3):(2'h3)]}));
                    end
                  else
                    begin
                      reg1218 <= ((+((forvar1198 ? forvar1207 : (8'hb8)) ?
                          reg1177[(4'h8):(1'h1)] : $signed(reg1224))) & reg1200[(4'he):(1'h1)]);
                      reg1219 <= $signed($signed({(forvar1193 ?
                              reg1171 : reg1182)}));
                      reg1220 <= $unsigned((+(8'hab)));
                      reg1221 <= (forvar1177[(2'h2):(1'h1)] >>> reg1187[(2'h2):(1'h0)]);
                    end
                  reg1222 <= wire1150[(4'h9):(3'h6)];
                  for (forvar1223 = (1'h0); (forvar1223 < (2'h3)); forvar1223 = (forvar1223 + (1'h1)))
                    begin
                      reg1224 <= $signed((+forvar1176));
                    end
                  if (reg1177[(4'he):(4'hd)])
                    begin
                      reg1225 <= {forvar1211};
                      reg1226 <= (~&(forvar1200[(3'h4):(2'h2)] ?
                          {(forvar1209 > reg1162)} : ($signed(reg1201) ?
                              $unsigned((8'ha8)) : (reg1184 != forvar1197))));
                      reg1227 <= $signed($signed((forvar1183 ?
                          (|wire1149) : $signed(reg1226))));
                      reg1228 <= {reg1178[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg1225 <= (-forvar1178);
                      reg1226 <= (reg1166[(1'h0):(1'h0)] + ((reg1227 & (-forvar1200)) & ((8'ha3) > (8'haf))));
                      reg1227 <= {(((~reg1169) ?
                                  reg1200[(4'hb):(4'h9)] : ((8'haa) <<< reg1215)) ?
                              (^reg1185) : reg1215)};
                    end
                end
              for (forvar1230 = (1'h0); (forvar1230 < (2'h2)); forvar1230 = (forvar1230 + (1'h1)))
                begin
                  for (forvar1231 = (1'h0); (forvar1231 < (1'h0)); forvar1231 = (forvar1231 + (1'h1)))
                    begin
                      reg1232 <= reg1211;
                      reg1233 <= forvar1227;
                      reg1234 <= $signed($signed((reg1211[(1'h0):(1'h0)] >>> reg1173[(2'h3):(2'h3)])));
                    end
                end
              for (forvar1235 = (1'h0); (forvar1235 < (2'h3)); forvar1235 = (forvar1235 + (1'h1)))
                begin
                  reg1236 <= reg1181[(1'h0):(1'h0)];
                end
              for (forvar1237 = (1'h0); (forvar1237 < (1'h1)); forvar1237 = (forvar1237 + (1'h1)))
                begin
                  if ($signed(($unsigned($signed(wire1150)) ?
                      (&{(8'ha0)}) : (!{(8'ha4)}))))
                    begin
                      reg1238 <= reg1232[(4'h8):(1'h0)];
                      reg1239 <= ($signed({reg1208[(1'h1):(1'h1)]}) ?
                          reg1211 : (($signed((8'ha5)) ^ forvar1162[(3'h4):(2'h2)]) ?
                              reg1171 : ((^~reg1220) ?
                                  forvar1201[(3'h4):(2'h3)] : {forvar1231})));
                      reg1240 <= $signed($unsigned(wire1151));
                      reg1241 <= $unsigned($unsigned((!$unsigned(reg1203))));
                    end
                  else
                    begin
                      reg1238 <= (~^((~(|(8'ha1))) ?
                          (+reg1236) : reg1185[(1'h1):(1'h0)]));
                      reg1239 <= $signed((~&$unsigned(forvar1231[(1'h1):(1'h1)])));
                      reg1240 <= reg1170[(1'h0):(1'h0)];
                    end
                  if ({((((8'hb1) >>> wire1150) ?
                              (&reg1198) : ((8'hb7) ? reg1233 : forvar1211)) ?
                          $unsigned($unsigned(reg1232)) : $unsigned(reg1233))})
                    begin
                      reg1242 <= ($signed(((+forvar1231) - (~|forvar1223))) & (((reg1163 > forvar1183) ?
                          $unsigned(wire1151) : reg1182) * $signed(reg1202[(1'h0):(1'h0)])));
                      reg1243 <= {forvar1183[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg1242 <= $signed($signed((^~(reg1185 > forvar1216))));
                      reg1243 <= $unsigned((forvar1199[(3'h5):(3'h4)] > (forvar1186[(1'h0):(1'h0)] ?
                          reg1199[(1'h1):(1'h1)] : (reg1160 ?
                              wire1155 : reg1178))));
                      reg1244 <= (reg1183 ?
                          ((~|(reg1221 != forvar1197)) <= (&$signed(reg1193))) : (reg1229 ?
                              wire1158[(1'h1):(1'h1)] : reg1176));
                      reg1245 <= ((&(^~(!forvar1176))) ?
                          ($signed((reg1167 ?
                              forvar1197 : wire1152)) << reg1206) : $unsigned({(|reg1173)}));
                    end
                  if ((-reg1225[(2'h2):(2'h2)]))
                    begin
                      reg1246 <= {({$unsigned(reg1225)} ?
                              $unsigned((-(8'hb5))) : $signed((~&reg1188)))};
                      reg1247 <= $signed(reg1168[(4'h8):(2'h2)]);
                      reg1248 <= reg1220[(4'hd):(4'hb)];
                    end
                  else
                    begin
                      reg1246 <= forvar1211[(1'h1):(1'h0)];
                    end
                  for (forvar1249 = (1'h0); (forvar1249 < (2'h3)); forvar1249 = (forvar1249 + (1'h1)))
                    begin
                      reg1250 <= {{$signed((+reg1192))}};
                    end
                end
            end
          reg1251 <= (8'ha8);
        end
      reg1252 <= $unsigned($signed($signed((reg1174 >= wire1151))));
      reg1253 <= (^~$signed(($unsigned(forvar1249) ?
          forvar1217[(3'h5):(3'h5)] : reg1196[(1'h0):(1'h0)])));
    end
  assign wire1254 = reg1167;
  assign wire1255 = $unsigned({((reg1180 * wire1152) ? (~|reg1204) : reg1163)});
  always
    @(posedge clk) begin
      for (forvar1256 = (1'h0); (forvar1256 < (1'h1)); forvar1256 = (forvar1256 + (1'h1)))
        begin
          for (forvar1257 = (1'h0); (forvar1257 < (1'h0)); forvar1257 = (forvar1257 + (1'h1)))
            begin
              for (forvar1258 = (1'h0); (forvar1258 < (1'h0)); forvar1258 = (forvar1258 + (1'h1)))
                begin
                  if ({wire1255})
                    begin
                      reg1259 <= $signed((-forvar1256));
                      reg1260 <= reg1244[(1'h0):(1'h0)];
                      reg1261 <= ((&$unsigned((reg1180 >> wire1151))) ?
                          reg1205[(3'h6):(1'h1)] : $signed($unsigned($signed(reg1238))));
                    end
                  else
                    begin
                      reg1259 <= reg1189;
                      reg1260 <= $unsigned($unsigned(reg1213[(3'h7):(2'h3)]));
                      reg1261 <= reg1179[(4'hd):(3'h7)];
                      reg1262 <= reg1219[(3'h4):(3'h4)];
                    end
                  for (forvar1263 = (1'h0); (forvar1263 < (2'h2)); forvar1263 = (forvar1263 + (1'h1)))
                    begin
                      reg1264 <= ({$unsigned($unsigned(reg1243))} == reg1212);
                      reg1265 <= (+reg1214);
                      reg1266 <= reg1170;
                      reg1267 <= (!reg1227);
                    end
                  for (forvar1268 = (1'h0); (forvar1268 < (1'h0)); forvar1268 = (forvar1268 + (1'h1)))
                    begin
                      reg1269 <= reg1239;
                      reg1270 <= {(8'hba)};
                    end
                end
              for (forvar1271 = (1'h0); (forvar1271 < (2'h3)); forvar1271 = (forvar1271 + (1'h1)))
                begin
                  if (((-{$unsigned(reg1220)}) && ($unsigned((reg1220 ?
                          reg1225 : reg1238)) ?
                      $signed((reg1252 | reg1250)) : $signed((reg1197 ?
                          wire1154 : forvar1268)))))
                    begin
                      reg1272 <= {(&((8'ha7) ? (-reg1183) : (-reg1171)))};
                      reg1273 <= reg1272;
                    end
                  else
                    begin
                      reg1272 <= (((reg1188 >= $signed(reg1218)) == reg1169[(3'h5):(1'h1)]) >= ((^~$signed(reg1165)) << ((!reg1195) < $signed(reg1186))));
                      reg1273 <= reg1161[(4'h9):(1'h0)];
                      reg1274 <= wire1255;
                      reg1275 <= $unsigned($unsigned((reg1224 ?
                          (reg1194 ~^ (8'hab)) : ((8'h9e) ?
                              (8'hac) : reg1166))));
                    end
                  if ($signed((&reg1161)))
                    begin
                      reg1276 <= $unsigned($signed(($signed(wire1157) | $unsigned(reg1241))));
                      reg1277 <= ((-$signed($unsigned((8'ha1)))) ?
                          $signed(reg1198) : reg1187[(4'hb):(3'h5)]);
                      reg1278 <= ((((reg1266 ?
                          reg1240 : forvar1258) >= wire1255[(1'h0):(1'h0)]) >> $unsigned((reg1170 ?
                          reg1196 : reg1208))) * ($signed((|forvar1271)) ?
                          (!(reg1213 >>> (8'hb5))) : (~&reg1167)));
                      reg1279 <= $unsigned((forvar1263[(1'h1):(1'h0)] * (~{reg1175})));
                    end
                  else
                    begin
                      reg1276 <= (~reg1183[(2'h3):(2'h3)]);
                    end
                  for (forvar1280 = (1'h0); (forvar1280 < (2'h3)); forvar1280 = (forvar1280 + (1'h1)))
                    begin
                      reg1281 <= $unsigned(reg1275[(5'h10):(3'h6)]);
                    end
                  for (forvar1282 = (1'h0); (forvar1282 < (1'h1)); forvar1282 = (forvar1282 + (1'h1)))
                    begin
                      reg1283 <= (($signed(wire1255) ?
                              $signed((reg1177 == reg1279)) : ($unsigned((8'ha5)) <= (!reg1281))) ?
                          $unsigned(wire1152[(4'h8):(2'h2)]) : reg1277[(4'hd):(3'h7)]);
                      reg1284 <= reg1266[(3'h4):(1'h0)];
                    end
                end
            end
          for (forvar1285 = (1'h0); (forvar1285 < (2'h2)); forvar1285 = (forvar1285 + (1'h1)))
            begin
              for (forvar1286 = (1'h0); (forvar1286 < (1'h0)); forvar1286 = (forvar1286 + (1'h1)))
                begin
                  for (forvar1287 = (1'h0); (forvar1287 < (1'h1)); forvar1287 = (forvar1287 + (1'h1)))
                    begin
                      reg1288 <= {$signed($signed((wire1156 ?
                              (8'hb7) : reg1172)))};
                      reg1289 <= $unsigned(reg1181[(2'h2):(1'h1)]);
                    end
                  for (forvar1290 = (1'h0); (forvar1290 < (1'h1)); forvar1290 = (forvar1290 + (1'h1)))
                    begin
                      reg1291 <= (({((8'h9f) ?
                              reg1181 : reg1281)} >= $signed((~reg1190))) * (&$signed($signed(wire1149))));
                      reg1292 <= $signed({((reg1183 ?
                              forvar1256 : reg1233) >>> $signed((8'ha4)))});
                      reg1293 <= (8'hba);
                      reg1294 <= $signed(reg1196[(1'h1):(1'h0)]);
                    end
                  reg1295 <= $unsigned($unsigned($unsigned((reg1179 ?
                      reg1177 : reg1164))));
                end
              reg1296 <= (~(-$signed({reg1228})));
            end
          for (forvar1297 = (1'h0); (forvar1297 < (2'h2)); forvar1297 = (forvar1297 + (1'h1)))
            begin
              for (forvar1298 = (1'h0); (forvar1298 < (1'h0)); forvar1298 = (forvar1298 + (1'h1)))
                begin
                  for (forvar1299 = (1'h0); (forvar1299 < (1'h1)); forvar1299 = (forvar1299 + (1'h1)))
                    begin
                      reg1300 <= $unsigned(((8'hac) ?
                          reg1266 : $unsigned($signed(reg1265))));
                      reg1301 <= $unsigned({reg1190[(3'h4):(1'h0)]});
                    end
                  for (forvar1302 = (1'h0); (forvar1302 < (1'h1)); forvar1302 = (forvar1302 + (1'h1)))
                    begin
                      reg1303 <= reg1233;
                    end
                  for (forvar1304 = (1'h0); (forvar1304 < (2'h3)); forvar1304 = (forvar1304 + (1'h1)))
                    begin
                      reg1305 <= {$signed(reg1166)};
                      reg1306 <= wire1155[(3'h6):(3'h6)];
                      reg1307 <= $signed((8'hb6));
                      reg1308 <= reg1261;
                    end
                end
              for (forvar1309 = (1'h0); (forvar1309 < (1'h1)); forvar1309 = (forvar1309 + (1'h1)))
                begin
                  for (forvar1310 = (1'h0); (forvar1310 < (2'h3)); forvar1310 = (forvar1310 + (1'h1)))
                    begin
                      reg1311 <= wire1158;
                      reg1312 <= (+$signed(($unsigned(forvar1257) << (forvar1287 ?
                          reg1238 : (8'hb6)))));
                      reg1313 <= $unsigned(reg1170[(1'h1):(1'h0)]);
                    end
                  reg1314 <= reg1234[(3'h4):(3'h4)];
                end
              for (forvar1315 = (1'h0); (forvar1315 < (2'h2)); forvar1315 = (forvar1315 + (1'h1)))
                begin
                  reg1316 <= reg1197[(1'h1):(1'h1)];
                  if (reg1191)
                    begin
                      reg1317 <= reg1221;
                      reg1318 <= reg1276[(1'h1):(1'h0)];
                      reg1319 <= ($unsigned(forvar1287[(3'h5):(3'h5)]) ?
                          forvar1271[(1'h0):(1'h0)] : wire1155[(4'ha):(4'h9)]);
                    end
                  else
                    begin
                      reg1317 <= {($unsigned((forvar1268 ?
                              (8'ha6) : reg1176)) ^ (wire1151[(3'h7):(3'h4)] ?
                              ((8'ha1) <= (8'had)) : $unsigned(reg1276)))};
                      reg1318 <= ($signed($signed($signed((8'hb4)))) << reg1292);
                      reg1319 <= wire1158[(4'h9):(3'h5)];
                    end
                  for (forvar1320 = (1'h0); (forvar1320 < (2'h2)); forvar1320 = (forvar1320 + (1'h1)))
                    begin
                      reg1321 <= ({((forvar1302 <= reg1178) >= reg1242[(1'h0):(1'h0)])} ?
                          {(reg1219 >>> $signed(wire1153))} : $signed(wire1158));
                      reg1322 <= reg1296[(3'h6):(1'h1)];
                      reg1323 <= (-$signed(((+(8'ha4)) >> ((8'hb5) - reg1232))));
                      reg1324 <= $unsigned((8'hb2));
                    end
                  if (forvar1256)
                    begin
                      reg1325 <= wire1254;
                      reg1326 <= $signed(reg1251);
                      reg1327 <= {(reg1260[(2'h3):(1'h0)] ?
                              ((reg1316 == reg1294) ?
                                  (reg1261 ?
                                      reg1272 : reg1206) : reg1184) : reg1194)};
                      reg1328 <= ($unsigned(($unsigned((8'h9f)) <= (reg1191 ^~ reg1238))) ~^ ($signed(reg1229[(4'h8):(3'h7)]) ?
                          (wire1157[(2'h3):(1'h0)] && ((8'h9d) ?
                              (8'hb7) : (8'hb0))) : forvar1282[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg1325 <= ((^$unsigned((&reg1222))) <<< (reg1328 & forvar1280[(3'h4):(2'h3)]));
                      reg1326 <= (~|(~^(~|(~|reg1198))));
                      reg1327 <= ((8'hb2) ?
                          $unsigned((~|(~&reg1171))) : (reg1192 == ($unsigned(reg1192) > (reg1180 ?
                              reg1205 : (8'hb6)))));
                    end
                end
              for (forvar1329 = (1'h0); (forvar1329 < (1'h1)); forvar1329 = (forvar1329 + (1'h1)))
                begin
                  for (forvar1330 = (1'h0); (forvar1330 < (1'h0)); forvar1330 = (forvar1330 + (1'h1)))
                    begin
                      reg1331 <= {((+wire1156[(1'h1):(1'h1)]) != $signed((reg1192 | reg1176)))};
                      reg1332 <= $signed({(~^$signed(wire1159))});
                      reg1333 <= {(forvar1309 != {{reg1224}})};
                      reg1334 <= $signed(($unsigned(reg1331[(3'h5):(1'h1)]) ?
                          ((reg1331 | reg1322) ?
                              $signed((8'ha5)) : {reg1288}) : (reg1215 || (wire1157 ?
                              reg1191 : forvar1330))));
                    end
                  for (forvar1335 = (1'h0); (forvar1335 < (1'h0)); forvar1335 = (forvar1335 + (1'h1)))
                    begin
                      reg1336 <= $signed($unsigned($signed($signed(reg1177))));
                    end
                  reg1337 <= ($unsigned($unsigned(((8'haf) ?
                      reg1241 : reg1334))) - $signed(reg1292[(3'h6):(1'h1)]));
                  if ($signed($unsigned($signed((reg1200 ?
                      reg1200 : reg1253)))))
                    begin
                      reg1338 <= reg1279;
                      reg1339 <= $signed(($unsigned((forvar1263 >>> reg1167)) << ($unsigned(reg1316) ?
                          reg1308 : (^reg1178))));
                    end
                  else
                    begin
                      reg1338 <= {($unsigned((reg1182 << reg1307)) - reg1262[(3'h7):(2'h3)])};
                      reg1339 <= $unsigned(($signed($signed(reg1171)) > (^reg1245)));
                      reg1340 <= (!{(reg1208[(1'h1):(1'h0)] != reg1300)});
                    end
                end
            end
        end
      for (forvar1341 = (1'h0); (forvar1341 < (2'h3)); forvar1341 = (forvar1341 + (1'h1)))
        begin
          for (forvar1342 = (1'h0); (forvar1342 < (1'h1)); forvar1342 = (forvar1342 + (1'h1)))
            begin
              if (reg1246)
                begin
                  reg1343 <= ($signed((8'ha8)) ? (+reg1269) : reg1182);
                  if (reg1284[(2'h2):(2'h2)])
                    begin
                      reg1344 <= ($unsigned(((reg1172 <<< reg1189) ^~ $unsigned(reg1168))) ?
                          (forvar1342[(1'h0):(1'h0)] ?
                              ($signed(forvar1329) ?
                                  {reg1241} : $signed(reg1169)) : reg1252[(1'h0):(1'h0)]) : (((reg1164 & reg1312) - (forvar1315 ^~ reg1278)) == (~|{(8'h9f)})));
                    end
                  else
                    begin
                      reg1344 <= ({{$unsigned(reg1184)}} + (^~($unsigned(forvar1286) != (~reg1198))));
                    end
                  for (forvar1345 = (1'h0); (forvar1345 < (1'h1)); forvar1345 = (forvar1345 + (1'h1)))
                    begin
                      reg1346 <= $signed({($signed(reg1322) ~^ (&reg1340))});
                      reg1347 <= (reg1170[(1'h0):(1'h0)] ^~ (~^$signed(reg1180)));
                      reg1348 <= ($signed(reg1316) ?
                          $signed(forvar1309[(3'h7):(1'h1)]) : (wire1255[(2'h2):(1'h0)] ?
                              (!$unsigned(wire1159)) : wire1156[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar1343 = (1'h0); (forvar1343 < (2'h3)); forvar1343 = (forvar1343 + (1'h1)))
                    begin
                      reg1344 <= $signed(reg1208);
                    end
                end
              for (forvar1349 = (1'h0); (forvar1349 < (2'h2)); forvar1349 = (forvar1349 + (1'h1)))
                begin
                  for (forvar1350 = (1'h0); (forvar1350 < (2'h2)); forvar1350 = (forvar1350 + (1'h1)))
                    begin
                      reg1351 <= ($unsigned((|reg1277)) ?
                          (reg1273[(3'h7):(3'h6)] ?
                              reg1251 : ((~|reg1164) ?
                                  (forvar1258 ?
                                      reg1205 : reg1162) : reg1277[(1'h0):(1'h0)])) : reg1174);
                    end
                  for (forvar1352 = (1'h0); (forvar1352 < (1'h1)); forvar1352 = (forvar1352 + (1'h1)))
                    begin
                      reg1353 <= (|{{(~&(8'ha4))}});
                      reg1354 <= ($unsigned($signed($unsigned(reg1294))) | ($signed(((8'ha6) ?
                          reg1188 : (8'hb8))) * reg1190));
                      reg1355 <= forvar1257[(1'h1):(1'h1)];
                    end
                  reg1356 <= reg1245;
                end
            end
          for (forvar1357 = (1'h0); (forvar1357 < (2'h2)); forvar1357 = (forvar1357 + (1'h1)))
            begin
              if ((((forvar1290 ^~ (reg1244 + reg1273)) <= $unsigned(reg1292)) >= ($signed((|reg1354)) ?
                  (-reg1259) : (&(reg1220 + reg1222)))))
                begin
                  if (reg1317)
                    begin
                      reg1358 <= ((~{(forvar1287 <<< wire1156)}) & reg1317[(3'h5):(3'h4)]);
                      reg1359 <= (((~|reg1356[(2'h2):(2'h2)]) > $unsigned(reg1294[(1'h1):(1'h0)])) ~^ reg1220[(3'h6):(3'h4)]);
                    end
                  else
                    begin
                      reg1358 <= ($signed(forvar1341) ?
                          (reg1250 == ($signed(reg1200) ?
                              (reg1262 << reg1321) : reg1272)) : (&reg1300[(3'h6):(2'h2)]));
                      reg1359 <= reg1229[(2'h2):(2'h2)];
                    end
                end
              else
                begin
                  if (($signed($unsigned((reg1162 >> reg1193))) != (~{reg1321[(3'h6):(1'h0)]})))
                    begin
                      reg1358 <= forvar1263;
                      reg1359 <= $signed({$signed($unsigned(reg1266))});
                      reg1360 <= $unsigned((reg1327 ?
                          $unsigned((^(8'ha5))) : ((!reg1265) ?
                              (~wire1153) : $unsigned((8'ha8)))));
                      reg1361 <= $unsigned($signed({reg1317}));
                    end
                  else
                    begin
                      reg1358 <= $unsigned(((-wire1254) || (+(reg1262 ?
                          (8'h9e) : (8'ha6)))));
                      reg1359 <= {reg1203};
                      reg1360 <= (reg1292[(1'h1):(1'h1)] ?
                          $signed((^((8'ha2) >>> reg1323))) : $signed($unsigned(reg1293)));
                      reg1361 <= {$unsigned($unsigned(reg1241))};
                    end
                  reg1362 <= (forvar1320[(1'h1):(1'h1)] - (((reg1220 ?
                      (8'ha7) : reg1283) | (reg1294 ?
                      reg1196 : (8'ha7))) < reg1344));
                  for (forvar1363 = (1'h0); (forvar1363 < (1'h1)); forvar1363 = (forvar1363 + (1'h1)))
                    begin
                      reg1364 <= (!$unsigned((|(+reg1210))));
                      reg1365 <= $signed($signed((~&(reg1180 ^~ reg1179))));
                      reg1366 <= reg1272[(1'h0):(1'h0)];
                      reg1367 <= forvar1335;
                    end
                end
              for (forvar1368 = (1'h0); (forvar1368 < (1'h0)); forvar1368 = (forvar1368 + (1'h1)))
                begin
                  for (forvar1369 = (1'h0); (forvar1369 < (2'h3)); forvar1369 = (forvar1369 + (1'h1)))
                    begin
                      reg1370 <= ($unsigned(reg1246) > (!(~^(~|(8'ha8)))));
                    end
                  reg1371 <= ($unsigned($unsigned((reg1338 ?
                          reg1347 : reg1295))) ?
                      $signed(reg1358[(2'h2):(2'h2)]) : $signed($unsigned((8'h9f))));
                  for (forvar1372 = (1'h0); (forvar1372 < (1'h0)); forvar1372 = (forvar1372 + (1'h1)))
                    begin
                      reg1373 <= $unsigned(reg1333);
                      reg1374 <= $signed($unsigned(reg1227));
                    end
                  reg1375 <= ((^~{$unsigned(wire1150)}) ?
                      $signed(($signed(reg1218) >= {reg1270})) : reg1200);
                end
            end
          for (forvar1376 = (1'h0); (forvar1376 < (2'h2)); forvar1376 = (forvar1376 + (1'h1)))
            begin
              if ($unsigned($signed($signed({reg1360}))))
                begin
                  if ($signed(reg1301[(1'h0):(1'h0)]))
                    begin
                      reg1377 <= (reg1316 >>> ($signed(wire1150[(4'h9):(3'h7)]) ?
                          ((~^reg1337) ?
                              $unsigned(reg1278) : reg1267) : reg1178));
                      reg1378 <= reg1214;
                    end
                  else
                    begin
                      reg1377 <= (+(^$unsigned(reg1233[(4'hb):(2'h3)])));
                      reg1378 <= ($unsigned(reg1323[(1'h0):(1'h0)]) | $signed($unsigned((reg1291 == reg1247))));
                      reg1379 <= reg1219;
                    end
                  if (wire1152[(4'he):(4'he)])
                    begin
                      reg1380 <= (!(8'hba));
                    end
                  else
                    begin
                      reg1380 <= (forvar1258[(1'h1):(1'h0)] && reg1343[(2'h3):(1'h1)]);
                      reg1381 <= $unsigned({($unsigned((8'hae)) && $signed(reg1308))});
                    end
                  reg1382 <= reg1171[(1'h1):(1'h1)];
                  if ((^~{{$signed(reg1176)}}))
                    begin
                      reg1383 <= $unsigned(({forvar1298[(3'h5):(2'h3)]} - (reg1228[(2'h3):(1'h1)] ?
                          (forvar1329 ? reg1358 : forvar1368) : {reg1215})));
                      reg1384 <= reg1208[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg1383 <= ($unsigned(((8'ha7) ?
                          (8'ha4) : $signed(reg1186))) <= ($signed(reg1227[(1'h1):(1'h1)]) ?
                          (8'ha1) : reg1179));
                      reg1384 <= (reg1266[(4'h8):(2'h3)] == $signed(reg1338));
                      reg1385 <= $unsigned(((!$signed(reg1226)) << $signed(reg1168)));
                    end
                end
              else
                begin
                  for (forvar1377 = (1'h0); (forvar1377 < (2'h2)); forvar1377 = (forvar1377 + (1'h1)))
                    begin
                      reg1378 <= reg1174[(1'h1):(1'h0)];
                      reg1379 <= forvar1299;
                    end
                end
              if (reg1379[(3'h4):(2'h3)])
                begin
                  for (forvar1386 = (1'h0); (forvar1386 < (2'h3)); forvar1386 = (forvar1386 + (1'h1)))
                    begin
                      reg1387 <= ({$signed(reg1358[(3'h6):(2'h2)])} | reg1204[(1'h0):(1'h0)]);
                      reg1388 <= (&reg1294);
                      reg1389 <= ((8'hb1) & reg1229);
                      reg1390 <= $signed(({$signed(reg1236)} ?
                          (&forvar1297) : reg1324[(2'h2):(1'h1)]));
                    end
                  reg1391 <= reg1375[(2'h3):(2'h2)];
                end
              else
                begin
                  reg1386 <= $unsigned(reg1200[(2'h2):(2'h2)]);
                end
            end
        end
      for (forvar1392 = (1'h0); (forvar1392 < (2'h2)); forvar1392 = (forvar1392 + (1'h1)))
        begin
          for (forvar1393 = (1'h0); (forvar1393 < (2'h3)); forvar1393 = (forvar1393 + (1'h1)))
            begin
              reg1394 <= wire1255;
              if ((^(!$unsigned((~(8'hb8))))))
                begin
                  for (forvar1395 = (1'h0); (forvar1395 < (2'h2)); forvar1395 = (forvar1395 + (1'h1)))
                    begin
                      reg1396 <= reg1218[(3'h5):(3'h4)];
                      reg1397 <= reg1339;
                      reg1398 <= $unsigned($unsigned(($signed((8'ha8)) ?
                          $signed(reg1253) : $signed(reg1242))));
                      reg1399 <= (forvar1363 ?
                          forvar1290 : {((reg1305 >> forvar1304) ?
                                  forvar1257[(2'h2):(2'h2)] : reg1308[(2'h3):(1'h1)])});
                    end
                end
              else
                begin
                  for (forvar1395 = (1'h0); (forvar1395 < (2'h3)); forvar1395 = (forvar1395 + (1'h1)))
                    begin
                      reg1396 <= reg1204[(2'h3):(2'h3)];
                      reg1397 <= (8'hb2);
                      reg1398 <= $unsigned({((reg1187 | reg1193) | (reg1295 - reg1203))});
                    end
                  if (forvar1329[(1'h0):(1'h0)])
                    begin
                      reg1399 <= (reg1161[(4'ha):(4'ha)] >> forvar1287[(3'h5):(3'h5)]);
                    end
                  else
                    begin
                      reg1399 <= forvar1377;
                      reg1400 <= $unsigned(((reg1277 < reg1163[(3'h6):(2'h3)]) ?
                          $signed(reg1172) : reg1228[(4'h8):(3'h6)]));
                      reg1401 <= {forvar1345};
                    end
                end
            end
          if ($unsigned(reg1184))
            begin
              for (forvar1402 = (1'h0); (forvar1402 < (1'h0)); forvar1402 = (forvar1402 + (1'h1)))
                begin
                  if (forvar1309)
                    begin
                      reg1403 <= (~&(&reg1201[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg1403 <= $unsigned((~(((8'hb4) ?
                          reg1181 : wire1157) + $signed(reg1210))));
                      reg1404 <= $unsigned(forvar1287);
                      reg1405 <= ($signed(forvar1299[(1'h0):(1'h0)]) ?
                          reg1187[(4'ha):(3'h4)] : reg1388[(2'h2):(2'h2)]);
                    end
                  if (reg1326[(1'h0):(1'h0)])
                    begin
                      reg1406 <= wire1157[(4'hd):(4'hb)];
                      reg1407 <= $unsigned(reg1259[(3'h5):(2'h3)]);
                    end
                  else
                    begin
                      reg1406 <= ($signed($unsigned((reg1366 ?
                              reg1325 : reg1405))) ?
                          reg1161[(4'hc):(1'h1)] : $signed(((~^reg1199) != $unsigned(reg1301))));
                      reg1407 <= reg1365[(4'h9):(3'h7)];
                      reg1408 <= $signed({($unsigned(forvar1286) ?
                              (|reg1177) : {reg1210})});
                    end
                  for (forvar1409 = (1'h0); (forvar1409 < (1'h1)); forvar1409 = (forvar1409 + (1'h1)))
                    begin
                      reg1410 <= ((((|(8'hae)) - reg1398[(2'h3):(2'h2)]) | $unsigned(reg1292)) ^~ reg1293);
                      reg1411 <= reg1261;
                    end
                end
              reg1412 <= reg1405;
            end
          else
            begin
              for (forvar1402 = (1'h0); (forvar1402 < (2'h3)); forvar1402 = (forvar1402 + (1'h1)))
                begin
                  reg1403 <= {$unsigned($unsigned((reg1279 ?
                          (8'ha5) : reg1179)))};
                  for (forvar1404 = (1'h0); (forvar1404 < (2'h3)); forvar1404 = (forvar1404 + (1'h1)))
                    begin
                      reg1405 <= reg1322[(2'h3):(1'h1)];
                      reg1406 <= (~|(((reg1267 ~^ wire1156) != ((8'ha1) ?
                              reg1273 : reg1401)) ?
                          forvar1297 : $unsigned((8'hb4))));
                      reg1407 <= $unsigned((^$unsigned(reg1305)));
                    end
                  if ($signed((($signed(reg1398) ?
                          (reg1222 ? reg1198 : reg1305) : (8'hb9)) ?
                      reg1193[(3'h6):(3'h6)] : ($unsigned(reg1367) < (~^reg1224)))))
                    begin
                      reg1408 <= (|reg1384[(4'hb):(1'h1)]);
                    end
                  else
                    begin
                      reg1408 <= (($signed((reg1303 >> reg1343)) & {{reg1292}}) + $unsigned($unsigned($signed((8'hb9)))));
                      reg1409 <= forvar1268[(1'h1):(1'h0)];
                    end
                end
              for (forvar1410 = (1'h0); (forvar1410 < (1'h0)); forvar1410 = (forvar1410 + (1'h1)))
                begin
                  for (forvar1411 = (1'h0); (forvar1411 < (1'h0)); forvar1411 = (forvar1411 + (1'h1)))
                    begin
                      reg1412 <= wire1149;
                      reg1413 <= (^~(~reg1403[(2'h2):(1'h0)]));
                      reg1414 <= $unsigned((|reg1383[(1'h0):(1'h0)]));
                      reg1415 <= $signed(((^~$unsigned(reg1227)) ?
                          ((&forvar1392) ?
                              forvar1369[(4'hb):(4'ha)] : $unsigned((8'had))) : $unsigned($unsigned((8'hb2)))));
                    end
                  for (forvar1416 = (1'h0); (forvar1416 < (1'h1)); forvar1416 = (forvar1416 + (1'h1)))
                    begin
                      reg1417 <= reg1238;
                      reg1418 <= reg1186;
                      reg1419 <= $unsigned(reg1325[(2'h3):(2'h3)]);
                    end
                  for (forvar1420 = (1'h0); (forvar1420 < (1'h1)); forvar1420 = (forvar1420 + (1'h1)))
                    begin
                      reg1421 <= ((^(reg1239[(2'h2):(1'h0)] ?
                          {(8'hab)} : (^(8'hb9)))) ~^ forvar1393[(3'h7):(1'h1)]);
                      reg1422 <= (reg1400[(3'h4):(1'h0)] ?
                          $unsigned($signed(reg1317)) : $unsigned(forvar1410));
                    end
                end
              reg1423 <= reg1252;
              reg1424 <= ({(reg1292[(3'h6):(2'h2)] + reg1198[(4'h9):(1'h1)])} | ((reg1171[(2'h3):(1'h1)] ?
                  $unsigned(forvar1341) : (wire1155 ?
                      (8'hb7) : forvar1349)) - ((reg1405 ?
                  reg1160 : reg1303) >>> (reg1359 ? forvar1392 : reg1325))));
            end
          if ((((forvar1352[(2'h3):(1'h0)] ? reg1424 : $unsigned(forvar1345)) ?
                  $signed($signed((8'haa))) : ((reg1199 ?
                      reg1373 : forvar1376) == $unsigned(reg1380))) ?
              ($signed(reg1176) * (reg1198[(4'h8):(1'h0)] ?
                  $unsigned((8'ha2)) : reg1303)) : reg1181))
            begin
              for (forvar1425 = (1'h0); (forvar1425 < (1'h0)); forvar1425 = (forvar1425 + (1'h1)))
                begin
                  reg1426 <= reg1167;
                  for (forvar1427 = (1'h0); (forvar1427 < (1'h1)); forvar1427 = (forvar1427 + (1'h1)))
                    begin
                      reg1428 <= {({reg1346} ? (8'hba) : $signed((8'hb4)))};
                    end
                end
              if (wire1254)
                begin
                  reg1429 <= $signed((8'ha5));
                  reg1430 <= $signed((reg1398[(4'hb):(4'h9)] && {(reg1170 * reg1407)}));
                  if ((^~reg1281))
                    begin
                      reg1431 <= reg1288;
                    end
                  else
                    begin
                      reg1431 <= (&reg1274);
                    end
                end
              else
                begin
                  for (forvar1429 = (1'h0); (forvar1429 < (2'h3)); forvar1429 = (forvar1429 + (1'h1)))
                    begin
                      reg1430 <= ((reg1422[(2'h3):(2'h3)] ?
                              (reg1343 - (reg1166 || reg1196)) : (reg1303 & reg1371[(1'h1):(1'h1)])) ?
                          (($unsigned(forvar1372) || (reg1233 && reg1406)) ?
                              ($unsigned((8'haf)) > (8'hb4)) : ((reg1160 ?
                                      reg1344 : reg1172) ?
                                  $unsigned(reg1408) : (reg1412 <<< reg1178))) : reg1193[(3'h6):(1'h1)]);
                      reg1431 <= (8'hb5);
                    end
                  reg1432 <= (^~(8'ha3));
                  for (forvar1433 = (1'h0); (forvar1433 < (1'h0)); forvar1433 = (forvar1433 + (1'h1)))
                    begin
                      reg1434 <= $unsigned(reg1222[(3'h4):(3'h4)]);
                    end
                end
            end
          else
            begin
              reg1425 <= reg1192;
              reg1426 <= {(reg1267 ?
                      ($unsigned(reg1196) ?
                          (forvar1310 ?
                              wire1157 : (8'hba)) : $signed(forvar1393)) : ((~reg1289) > (+(8'ha9))))};
              for (forvar1427 = (1'h0); (forvar1427 < (2'h2)); forvar1427 = (forvar1427 + (1'h1)))
                begin
                  reg1428 <= reg1168;
                  for (forvar1429 = (1'h0); (forvar1429 < (1'h1)); forvar1429 = (forvar1429 + (1'h1)))
                    begin
                      reg1430 <= $signed(reg1316[(5'h10):(4'hb)]);
                    end
                  reg1431 <= (^$signed($signed((~&reg1407))));
                end
            end
        end
      for (forvar1435 = (1'h0); (forvar1435 < (2'h3)); forvar1435 = (forvar1435 + (1'h1)))
        begin
          for (forvar1436 = (1'h0); (forvar1436 < (1'h1)); forvar1436 = (forvar1436 + (1'h1)))
            begin
              for (forvar1437 = (1'h0); (forvar1437 < (2'h2)); forvar1437 = (forvar1437 + (1'h1)))
                begin
                  reg1438 <= (($signed(forvar1263[(1'h1):(1'h1)]) || (!reg1166)) ?
                      {reg1288} : reg1434[(4'h8):(3'h6)]);
                  for (forvar1439 = (1'h0); (forvar1439 < (2'h3)); forvar1439 = (forvar1439 + (1'h1)))
                    begin
                      reg1440 <= {reg1431};
                      reg1441 <= $unsigned(forvar1341);
                    end
                end
              reg1442 <= $signed(reg1306);
              for (forvar1443 = (1'h0); (forvar1443 < (1'h0)); forvar1443 = (forvar1443 + (1'h1)))
                begin
                  reg1444 <= (~|forvar1429);
                  if ($unsigned(($unsigned(forvar1357) >= reg1359[(3'h5):(1'h1)])))
                    begin
                      reg1445 <= {$unsigned({$unsigned(reg1316)})};
                      reg1446 <= $signed((8'ha8));
                      reg1447 <= (forvar1343 ?
                          reg1284[(1'h0):(1'h0)] : reg1167[(3'h4):(2'h2)]);
                      reg1448 <= reg1312[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg1445 <= forvar1350;
                      reg1446 <= (reg1223[(3'h5):(2'h3)] ?
                          $signed($unsigned((|reg1288))) : $unsigned(($signed(wire1150) != (reg1202 ?
                              forvar1436 : reg1410))));
                      reg1447 <= $signed(reg1390);
                      reg1448 <= ((((^~reg1226) ?
                              $signed(reg1164) : $unsigned(reg1444)) <= $unsigned(((8'haa) ?
                              reg1385 : reg1422))) ?
                          reg1358[(2'h2):(1'h1)] : (+$signed((reg1227 ?
                              reg1375 : reg1319))));
                    end
                end
            end
          for (forvar1449 = (1'h0); (forvar1449 < (1'h0)); forvar1449 = (forvar1449 + (1'h1)))
            begin
              for (forvar1450 = (1'h0); (forvar1450 < (1'h1)); forvar1450 = (forvar1450 + (1'h1)))
                begin
                  if ((~&$signed(forvar1345)))
                    begin
                      reg1451 <= reg1225;
                      reg1452 <= {$unsigned((((8'ha6) << (8'hb2)) || $signed(reg1430)))};
                      reg1453 <= {$signed({(reg1265 << reg1306)})};
                    end
                  else
                    begin
                      reg1451 <= (~&(8'h9c));
                      reg1452 <= reg1251;
                    end
                end
              for (forvar1454 = (1'h0); (forvar1454 < (1'h1)); forvar1454 = (forvar1454 + (1'h1)))
                begin
                  for (forvar1455 = (1'h0); (forvar1455 < (2'h3)); forvar1455 = (forvar1455 + (1'h1)))
                    begin
                      reg1456 <= $signed($signed(reg1233[(1'h1):(1'h1)]));
                    end
                  if ({(reg1407 ^ (8'ha7))})
                    begin
                      reg1457 <= reg1391;
                      reg1458 <= (((forvar1402 << (~^(8'had))) ?
                              reg1200 : (-reg1373[(3'h5):(2'h3)])) ?
                          ((~(^reg1197)) ?
                              ((~|reg1374) != $signed((8'hab))) : $signed(reg1340[(4'ha):(3'h4)])) : reg1381);
                      reg1459 <= wire1159;
                    end
                  else
                    begin
                      reg1457 <= reg1197[(1'h0):(1'h0)];
                    end
                  for (forvar1460 = (1'h0); (forvar1460 < (1'h1)); forvar1460 = (forvar1460 + (1'h1)))
                    begin
                      reg1461 <= (($unsigned((-reg1346)) != $signed($signed(forvar1280))) ?
                          {$unsigned({reg1318})} : ($signed($unsigned((8'hb9))) >= (8'hb6)));
                      reg1462 <= (^~$signed($unsigned(reg1226)));
                      reg1463 <= (($unsigned((|(8'ha1))) * $signed((reg1403 - forvar1411))) ?
                          (!(^~reg1458[(4'h9):(3'h6)])) : $signed((+(reg1397 ?
                              forvar1315 : forvar1268))));
                    end
                end
            end
        end
    end
  assign wire1464 = reg1198;
  always
    @(posedge clk) begin
      if ((~^reg1424[(2'h2):(1'h1)]))
        begin
          for (forvar1465 = (1'h0); (forvar1465 < (2'h2)); forvar1465 = (forvar1465 + (1'h1)))
            begin
              for (forvar1466 = (1'h0); (forvar1466 < (1'h0)); forvar1466 = (forvar1466 + (1'h1)))
                begin
                  reg1467 <= reg1314[(4'h8):(2'h2)];
                end
            end
          reg1468 <= reg1426;
        end
      else
        begin
          for (forvar1465 = (1'h0); (forvar1465 < (1'h1)); forvar1465 = (forvar1465 + (1'h1)))
            begin
              reg1466 <= $unsigned({{(8'haa)}});
              for (forvar1467 = (1'h0); (forvar1467 < (2'h2)); forvar1467 = (forvar1467 + (1'h1)))
                begin
                  if ($unsigned($signed((!$unsigned(reg1383)))))
                    begin
                      reg1468 <= reg1233[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1468 <= {(((reg1196 | reg1164) ?
                              $signed(reg1425) : reg1440) >> reg1390)};
                      reg1469 <= $signed((~^reg1305[(2'h2):(1'h0)]));
                      reg1470 <= ((($unsigned(reg1182) ?
                              (^reg1332) : (~^reg1452)) ^ (reg1211[(1'h0):(1'h0)] ?
                              (reg1165 != reg1311) : reg1283)) ?
                          $unsigned((^$unsigned(wire1159))) : $unsigned({(reg1394 ^ (8'hb4))}));
                    end
                  for (forvar1471 = (1'h0); (forvar1471 < (1'h0)); forvar1471 = (forvar1471 + (1'h1)))
                    begin
                      reg1472 <= $signed((^$unsigned(reg1348[(4'h9):(2'h3)])));
                      reg1473 <= ({((!wire1464) ? (~|reg1324) : reg1205)} ?
                          ($unsigned($unsigned(reg1243)) ~^ (reg1414[(2'h2):(1'h1)] ?
                              (reg1409 ?
                                  reg1314 : reg1266) : (reg1233 + (8'ha7)))) : (reg1452 ?
                              forvar1466[(2'h2):(2'h2)] : reg1328));
                      reg1474 <= $unsigned((reg1470[(3'h5):(1'h1)] ?
                          (&(reg1265 - reg1371)) : ($unsigned(reg1377) ~^ $unsigned(reg1351))));
                    end
                end
              if (reg1162[(1'h0):(1'h0)])
                begin
                  for (forvar1475 = (1'h0); (forvar1475 < (1'h0)); forvar1475 = (forvar1475 + (1'h1)))
                    begin
                      reg1476 <= (-(^$unsigned(wire1156[(2'h3):(2'h2)])));
                      reg1477 <= (!reg1334[(2'h2):(1'h1)]);
                      reg1478 <= (!{(&(+reg1462))});
                    end
                  if (reg1384)
                    begin
                      reg1479 <= ((-$signed({reg1434})) ?
                          (~|reg1233[(3'h4):(2'h3)]) : (8'ha4));
                      reg1480 <= (reg1318[(3'h4):(2'h2)] ?
                          ({reg1184} >>> reg1355) : $signed((reg1191[(1'h0):(1'h0)] * ((8'ha3) ?
                              reg1346 : reg1223))));
                      reg1481 <= ($signed((-reg1198)) ?
                          (reg1168 - (reg1252 >>> reg1407)) : ($unsigned($unsigned(reg1276)) ?
                              reg1480 : ((reg1178 ? reg1401 : reg1399) ?
                                  reg1371 : {(8'had)})));
                    end
                  else
                    begin
                      reg1479 <= $unsigned({$signed($signed(wire1154))});
                      reg1480 <= $unsigned((reg1367 ^~ (reg1343[(3'h6):(1'h0)] ?
                          $signed((8'had)) : {reg1300})));
                      reg1481 <= (|$unsigned((~^(reg1187 ~^ reg1472))));
                      reg1482 <= (^~($signed(reg1251[(2'h2):(1'h0)]) < (((8'hb4) ?
                          wire1151 : forvar1475) && $unsigned(reg1218))));
                    end
                end
              else
                begin
                  for (forvar1475 = (1'h0); (forvar1475 < (2'h2)); forvar1475 = (forvar1475 + (1'h1)))
                    begin
                      reg1476 <= reg1411;
                      reg1477 <= (~&(+$unsigned((reg1481 ?
                          reg1401 : reg1203))));
                      reg1478 <= $signed((8'had));
                      reg1479 <= $unsigned({((8'hab) ?
                              reg1417 : $signed(reg1468))});
                    end
                  if ($signed((wire1155[(3'h5):(3'h4)] ^~ reg1388[(4'he):(2'h2)])))
                    begin
                      reg1480 <= $signed($unsigned((8'hb0)));
                      reg1481 <= reg1331;
                      reg1482 <= ((((-reg1331) | $unsigned(reg1373)) ?
                          ((+reg1374) ?
                              reg1432 : wire1464[(4'h9):(3'h5)]) : ((^~reg1185) ?
                              (reg1424 | reg1278) : reg1459[(2'h3):(1'h0)])) * (8'ha4));
                      reg1483 <= {(reg1175 ?
                              $unsigned({(8'ha8)}) : $unsigned((reg1365 ?
                                  reg1343 : reg1233)))};
                    end
                  else
                    begin
                      reg1480 <= $unsigned(reg1483[(4'hb):(3'h4)]);
                      reg1481 <= {{(~|reg1346[(4'hb):(2'h2)])}};
                      reg1482 <= {$signed(((|reg1483) ?
                              $unsigned(reg1198) : reg1179))};
                      reg1483 <= $unsigned((&((wire1150 ? reg1326 : reg1379) ?
                          (reg1388 ^ reg1379) : $unsigned((8'ha6)))));
                    end
                  for (forvar1484 = (1'h0); (forvar1484 < (1'h1)); forvar1484 = (forvar1484 + (1'h1)))
                    begin
                      reg1485 <= ({(-reg1183[(2'h2):(1'h1)])} << $signed(reg1414[(4'h8):(4'h8)]));
                    end
                end
              if (((-((reg1319 ? reg1269 : (8'hb5)) ?
                  $signed(reg1189) : (reg1364 + reg1467))) <<< $unsigned((~|(|(8'haf))))))
                begin
                  reg1486 <= ((!(reg1396[(4'h8):(3'h6)] ?
                      {reg1267} : (reg1390 & reg1227))) > $unsigned(($unsigned(reg1424) ?
                      {reg1412} : reg1196[(3'h4):(1'h0)])));
                  if (reg1374)
                    begin
                      reg1487 <= $unsigned(reg1370);
                      reg1488 <= ($unsigned((~forvar1467[(1'h1):(1'h1)])) ?
                          reg1164[(2'h3):(2'h3)] : {((|reg1365) ?
                                  (reg1384 ~^ reg1353) : $unsigned(reg1238))});
                      reg1489 <= (8'hab);
                    end
                  else
                    begin
                      reg1487 <= $signed(reg1396[(3'h7):(1'h0)]);
                      reg1488 <= ((+reg1233) ?
                          (wire1150[(3'h7):(2'h3)] ?
                              $signed(reg1291[(3'h7):(3'h5)]) : $signed({reg1228})) : reg1219);
                      reg1489 <= {{(|reg1185)}};
                    end
                  for (forvar1490 = (1'h0); (forvar1490 < (2'h2)); forvar1490 = (forvar1490 + (1'h1)))
                    begin
                      reg1491 <= reg1165[(2'h2):(1'h1)];
                      reg1492 <= ($unsigned($unsigned(wire1254[(4'h8):(1'h1)])) >>> $unsigned((-$unsigned(reg1338))));
                    end
                end
              else
                begin
                  if ($unsigned((+(reg1347 >> reg1184))))
                    begin
                      reg1486 <= $signed((wire1156 ?
                          reg1211[(1'h1):(1'h1)] : $signed($signed(reg1206))));
                      reg1487 <= (~|reg1232);
                      reg1488 <= $unsigned(reg1245[(4'h9):(4'h8)]);
                      reg1489 <= (reg1405 != $signed(reg1488));
                    end
                  else
                    begin
                      reg1486 <= $signed(($unsigned((~(8'hb2))) ?
                          ((reg1218 ? (8'hb9) : reg1358) ?
                              (reg1314 || reg1456) : $signed((8'ha5))) : $unsigned(reg1404)));
                      reg1487 <= $signed((reg1328[(2'h2):(1'h0)] ?
                          $signed(reg1448[(4'ha):(2'h3)]) : (8'hb1)));
                    end
                  if ((+$signed(($unsigned(reg1250) & $unsigned(reg1438)))))
                    begin
                      reg1490 <= ((((reg1279 - reg1438) ^~ $signed(wire1158)) < (~$signed(reg1452))) ?
                          ($signed(reg1383[(2'h2):(2'h2)]) == $unsigned($signed(reg1379))) : (8'h9e));
                      reg1491 <= $signed(reg1283[(2'h2):(2'h2)]);
                      reg1492 <= ({((reg1453 ?
                              reg1170 : reg1406) ^~ reg1313)} <<< {reg1487});
                      reg1493 <= (~|(reg1165[(2'h2):(1'h1)] ?
                          {{reg1227}} : (-$unsigned(reg1404))));
                    end
                  else
                    begin
                      reg1490 <= $signed(((!$signed(reg1404)) || $unsigned((reg1384 && reg1225))));
                      reg1491 <= {(8'hb2)};
                      reg1492 <= $signed(((+$signed(reg1245)) >= ({reg1276} ?
                          (reg1348 >> reg1332) : reg1444)));
                      reg1493 <= reg1477;
                    end
                  if ((reg1196 > reg1431[(2'h2):(1'h1)]))
                    begin
                      reg1494 <= reg1184[(3'h4):(1'h1)];
                      reg1495 <= (~(reg1481[(1'h0):(1'h0)] && (reg1166 ?
                          (reg1259 && reg1456) : reg1338[(4'h9):(1'h0)])));
                    end
                  else
                    begin
                      reg1494 <= (~|(($unsigned(reg1186) ?
                          (reg1390 < wire1159) : reg1351[(1'h1):(1'h0)]) != ((reg1279 || reg1175) && $signed(reg1481))));
                      reg1495 <= (wire1154 ? {reg1245} : forvar1475);
                      reg1496 <= $unsigned(forvar1475[(3'h4):(2'h3)]);
                    end
                  for (forvar1497 = (1'h0); (forvar1497 < (1'h1)); forvar1497 = (forvar1497 + (1'h1)))
                    begin
                      reg1498 <= (forvar1484 ?
                          ((!reg1325) ?
                              $signed($signed(reg1228)) : {{reg1343}}) : (!$signed($signed(reg1496))));
                      reg1499 <= (&$signed($signed($unsigned(reg1267))));
                      reg1500 <= (wire1156 ?
                          {((reg1398 ? wire1159 : reg1366) ?
                                  (reg1442 ? reg1190 : reg1191) : (reg1221 ?
                                      reg1448 : reg1371))} : reg1232[(1'h1):(1'h1)]);
                      reg1501 <= reg1169;
                    end
                end
            end
          reg1502 <= (|reg1222[(2'h2):(1'h1)]);
          if ((reg1191 != (8'hb3)))
            begin
              if ({$unsigned(reg1301[(3'h7):(3'h4)])})
                begin
                  for (forvar1503 = (1'h0); (forvar1503 < (2'h3)); forvar1503 = (forvar1503 + (1'h1)))
                    begin
                      reg1504 <= ($unsigned(((~&(8'hb7)) ?
                              $unsigned(reg1289) : (reg1288 - reg1167))) ?
                          {reg1312} : (8'hb5));
                      reg1505 <= ($unsigned($unsigned($signed(reg1293))) ?
                          (!$unsigned((~&reg1466))) : {reg1266[(1'h1):(1'h1)]});
                      reg1506 <= reg1185[(3'h4):(2'h3)];
                      reg1507 <= {(~(8'haf))};
                    end
                  for (forvar1508 = (1'h0); (forvar1508 < (2'h2)); forvar1508 = (forvar1508 + (1'h1)))
                    begin
                      reg1509 <= (($unsigned($unsigned((8'h9e))) == $unsigned(reg1177)) ^~ reg1208);
                      reg1510 <= $signed(({(~^wire1157)} <<< $unsigned(reg1407)));
                      reg1511 <= reg1489[(2'h3):(2'h2)];
                      reg1512 <= reg1505[(3'h4):(3'h4)];
                    end
                  reg1513 <= $signed(reg1340[(1'h1):(1'h1)]);
                  for (forvar1514 = (1'h0); (forvar1514 < (2'h2)); forvar1514 = (forvar1514 + (1'h1)))
                    begin
                      reg1515 <= (((wire1156[(1'h0):(1'h0)] ?
                              (reg1164 ~^ reg1204) : $signed(reg1200)) ?
                          reg1378 : (&reg1374)) + reg1222);
                      reg1516 <= $unsigned(reg1259);
                      reg1517 <= (!(~&(&(reg1248 >= reg1214))));
                    end
                end
              else
                begin
                  for (forvar1503 = (1'h0); (forvar1503 < (1'h0)); forvar1503 = (forvar1503 + (1'h1)))
                    begin
                      reg1504 <= $unsigned($signed((!(reg1212 * reg1316))));
                      reg1505 <= $signed(reg1322);
                      reg1506 <= (reg1354 | $unsigned(((&reg1494) ?
                          reg1181[(3'h6):(3'h5)] : reg1421)));
                    end
                  for (forvar1507 = (1'h0); (forvar1507 < (2'h2)); forvar1507 = (forvar1507 + (1'h1)))
                    begin
                      reg1508 <= reg1176[(4'ha):(3'h5)];
                      reg1509 <= (((!(8'ha9)) <<< wire1155[(1'h0):(1'h0)]) < (~&{$signed(reg1375)}));
                      reg1510 <= $signed({(-$unsigned(reg1253))});
                      reg1511 <= reg1339[(4'hb):(3'h6)];
                    end
                  for (forvar1512 = (1'h0); (forvar1512 < (1'h1)); forvar1512 = (forvar1512 + (1'h1)))
                    begin
                      reg1513 <= ((&$signed($unsigned(forvar1507))) ^~ $signed($signed((^reg1264))));
                      reg1514 <= ((((reg1311 >= reg1206) | $unsigned(reg1397)) >= (~&(reg1423 ?
                          (8'ha2) : (8'hb1)))) == reg1492);
                      reg1515 <= (~reg1166[(3'h4):(2'h3)]);
                      reg1516 <= $unsigned((~&reg1166[(3'h4):(1'h1)]));
                    end
                  for (forvar1517 = (1'h0); (forvar1517 < (1'h0)); forvar1517 = (forvar1517 + (1'h1)))
                    begin
                      reg1518 <= (($signed($unsigned(reg1301)) || $signed(reg1434[(4'ha):(4'h8)])) ?
                          $signed({{reg1451}}) : reg1354);
                      reg1519 <= ((($unsigned(reg1195) ?
                                  {reg1303} : reg1485[(4'hc):(4'ha)]) ?
                              reg1334 : (reg1381 ?
                                  reg1214[(4'h8):(3'h6)] : (~^(8'h9e)))) ?
                          reg1295 : (reg1373[(3'h7):(3'h7)] < (~(reg1397 | (8'hb7)))));
                      reg1520 <= $signed((-$unsigned((+(8'ha6)))));
                    end
                end
              for (forvar1521 = (1'h0); (forvar1521 < (2'h2)); forvar1521 = (forvar1521 + (1'h1)))
                begin
                  for (forvar1522 = (1'h0); (forvar1522 < (2'h2)); forvar1522 = (forvar1522 + (1'h1)))
                    begin
                      reg1523 <= (8'h9d);
                    end
                  if ((~|$unsigned(reg1264[(3'h5):(1'h0)])))
                    begin
                      reg1524 <= ((reg1172[(2'h2):(1'h0)] >> (~|(reg1469 << reg1167))) + reg1421);
                      reg1525 <= (|reg1398);
                      reg1526 <= $signed(reg1224);
                      reg1527 <= reg1358[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg1524 <= (&reg1461[(3'h6):(3'h5)]);
                      reg1525 <= $signed((^(~^$unsigned(reg1483))));
                    end
                end
            end
          else
            begin
              if ((reg1379[(2'h3):(1'h0)] >> $signed(wire1254[(1'h1):(1'h0)])))
                begin
                  if (((reg1276[(1'h0):(1'h0)] ?
                      ($unsigned(reg1451) ?
                          (reg1334 & wire1157) : $signed(reg1214)) : $signed(reg1422)) > $unsigned(reg1422)))
                    begin
                      reg1503 <= reg1391;
                      reg1504 <= reg1208;
                    end
                  else
                    begin
                      reg1503 <= $signed((((reg1380 ?
                              reg1520 : reg1428) ^~ (&forvar1490)) ?
                          (((8'ha3) ? reg1466 : reg1325) ?
                              (reg1223 & reg1243) : (reg1324 ?
                                  reg1527 : reg1502)) : reg1279[(2'h2):(1'h0)]));
                      reg1504 <= reg1367;
                    end
                  for (forvar1505 = (1'h0); (forvar1505 < (1'h0)); forvar1505 = (forvar1505 + (1'h1)))
                    begin
                      reg1506 <= ($unsigned(((wire1154 | reg1293) <<< $unsigned((8'hac)))) < $unsigned(reg1390));
                    end
                  if ((8'hb9))
                    begin
                      reg1507 <= {reg1274[(2'h2):(1'h1)]};
                      reg1508 <= (({forvar1514} ?
                          (^(^reg1389)) : ((reg1181 >= reg1200) ?
                              $unsigned(wire1149) : $unsigned((8'ha3)))) <<< (reg1241[(1'h0):(1'h0)] < $signed((reg1312 & forvar1517))));
                      reg1509 <= $signed((^~$signed(((8'ha2) <<< reg1406))));
                      reg1510 <= reg1370[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg1507 <= $signed({((reg1305 ?
                              reg1409 : reg1288) * $unsigned(forvar1512))});
                      reg1508 <= reg1236;
                    end
                  for (forvar1511 = (1'h0); (forvar1511 < (2'h2)); forvar1511 = (forvar1511 + (1'h1)))
                    begin
                      reg1512 <= {(-$unsigned(forvar1466))};
                      reg1513 <= (reg1415[(1'h1):(1'h0)] ?
                          ((((8'ha0) ? reg1485 : (8'hb1)) ?
                                  (!forvar1475) : (reg1169 && (8'hb9))) ?
                              (!(!reg1199)) : reg1403) : $signed((-(^~reg1340))));
                      reg1514 <= (reg1512[(4'hc):(4'h9)] ?
                          reg1451[(3'h4):(3'h4)] : $signed(((reg1419 || reg1236) + reg1351)));
                      reg1515 <= reg1448;
                    end
                end
              else
                begin
                  if (reg1383[(2'h2):(2'h2)])
                    begin
                      reg1503 <= ($unsigned({reg1228}) ?
                          reg1495 : ($unsigned((reg1441 << reg1346)) ?
                              (^~(forvar1521 <<< (8'ha2))) : $unsigned(reg1314[(1'h0):(1'h0)])));
                      reg1504 <= (reg1339 ? reg1269 : $signed(forvar1484));
                      reg1505 <= wire1255;
                      reg1506 <= reg1242[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1503 <= $unsigned({forvar1507});
                      reg1504 <= ((+reg1385) ?
                          $signed((reg1361 ?
                              reg1245 : reg1421[(4'h8):(3'h6)])) : $signed((|reg1305)));
                      reg1505 <= reg1264[(3'h7):(3'h5)];
                    end
                end
            end
        end
      if ($signed(reg1401))
        begin
          for (forvar1528 = (1'h0); (forvar1528 < (1'h0)); forvar1528 = (forvar1528 + (1'h1)))
            begin
              reg1529 <= reg1364;
              for (forvar1530 = (1'h0); (forvar1530 < (2'h2)); forvar1530 = (forvar1530 + (1'h1)))
                begin
                  if ($signed($signed((|(reg1359 ? reg1162 : reg1513)))))
                    begin
                      reg1531 <= {$unsigned(reg1182[(1'h1):(1'h0)])};
                      reg1532 <= {reg1391};
                      reg1533 <= {reg1246};
                      reg1534 <= (($signed(reg1424[(1'h1):(1'h0)]) ?
                              (~^((8'ha5) ? (8'hb0) : reg1228)) : (reg1459 ?
                                  reg1377[(2'h3):(2'h3)] : (~^reg1179))) ?
                          {(reg1221 ?
                                  $unsigned(reg1289) : (reg1206 ^~ reg1332))} : $signed((reg1327[(3'h7):(3'h6)] < $signed(reg1208))));
                    end
                  else
                    begin
                      reg1531 <= $signed($signed(reg1172[(2'h2):(2'h2)]));
                    end
                  if ($unsigned((reg1198 < (|reg1337))))
                    begin
                      reg1535 <= (reg1279[(3'h6):(2'h2)] ?
                          reg1333 : (^~({reg1295} ?
                              reg1480[(2'h3):(1'h0)] : (reg1166 < reg1313))));
                      reg1536 <= forvar1471;
                      reg1537 <= ((~&($signed((8'ha1)) ?
                              {reg1337} : (~|reg1224))) ?
                          (+{{reg1192}}) : reg1222[(1'h0):(1'h0)]);
                      reg1538 <= ($signed({reg1227[(3'h6):(2'h3)]}) ?
                          {forvar1514[(2'h3):(1'h1)]} : ($unsigned(reg1425[(3'h5):(3'h4)]) * (^$signed(wire1464))));
                    end
                  else
                    begin
                      reg1535 <= ($unsigned(({(8'hb5)} ?
                              ((8'hba) ? reg1527 : (8'hb4)) : (8'ha3))) ?
                          reg1407[(2'h3):(2'h2)] : $signed({$signed(reg1273)}));
                      reg1536 <= ((($signed(reg1267) ?
                              $signed((8'ha4)) : (reg1201 ?
                                  reg1174 : reg1444)) ?
                          (~reg1169[(4'h8):(4'h8)]) : {$unsigned(reg1496)}) + (^$unsigned($unsigned(forvar1507))));
                      reg1537 <= ((~|((forvar1475 ? (8'had) : reg1441) ?
                          $signed(reg1356) : reg1198)) && reg1164);
                      reg1538 <= {(~($signed(reg1422) * (reg1305 ?
                              reg1198 : reg1206)))};
                    end
                  for (forvar1539 = (1'h0); (forvar1539 < (1'h0)); forvar1539 = (forvar1539 + (1'h1)))
                    begin
                      reg1540 <= {(reg1456[(2'h2):(2'h2)] & {(^wire1158)})};
                      reg1541 <= (8'ha5);
                    end
                  for (forvar1542 = (1'h0); (forvar1542 < (1'h1)); forvar1542 = (forvar1542 + (1'h1)))
                    begin
                      reg1543 <= $unsigned((!(-(&reg1311))));
                      reg1544 <= reg1240[(1'h1):(1'h0)];
                    end
                end
              for (forvar1545 = (1'h0); (forvar1545 < (2'h3)); forvar1545 = (forvar1545 + (1'h1)))
                begin
                  for (forvar1546 = (1'h0); (forvar1546 < (2'h3)); forvar1546 = (forvar1546 + (1'h1)))
                    begin
                      reg1547 <= reg1221[(2'h3):(1'h0)];
                      reg1548 <= (&{$signed((&reg1519))});
                    end
                  for (forvar1549 = (1'h0); (forvar1549 < (2'h2)); forvar1549 = (forvar1549 + (1'h1)))
                    begin
                      reg1550 <= reg1202;
                      reg1551 <= $signed(($unsigned($signed(reg1541)) >> ($signed(reg1265) ?
                          $signed(reg1307) : $signed(reg1242))));
                    end
                  if (reg1446)
                    begin
                      reg1552 <= $unsigned($unsigned(reg1317));
                      reg1553 <= reg1411[(1'h1):(1'h0)];
                      reg1554 <= reg1359[(1'h0):(1'h0)];
                      reg1555 <= ($signed(((reg1180 + (8'ha9)) ~^ (reg1354 ?
                              reg1526 : reg1456))) ?
                          $unsigned(wire1159[(3'h5):(1'h0)]) : reg1202[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1552 <= reg1425;
                      reg1553 <= $unsigned((&($signed(reg1184) - reg1387)));
                    end
                  if ($unsigned((-(~(reg1221 ? reg1364 : reg1527)))))
                    begin
                      reg1556 <= $signed((reg1389[(4'he):(3'h4)] ?
                          ((reg1488 > reg1430) ?
                              reg1336 : $signed(reg1487)) : (reg1456[(2'h2):(1'h1)] ?
                              $unsigned(reg1513) : reg1327[(1'h0):(1'h0)])));
                      reg1557 <= (reg1184[(4'h8):(4'h8)] * {reg1344});
                    end
                  else
                    begin
                      reg1556 <= ($unsigned({(reg1346 ?
                              reg1300 : reg1535)}) | {$signed(((8'ha9) ?
                              reg1384 : reg1473))});
                    end
                end
            end
          for (forvar1558 = (1'h0); (forvar1558 < (1'h0)); forvar1558 = (forvar1558 + (1'h1)))
            begin
              for (forvar1559 = (1'h0); (forvar1559 < (2'h2)); forvar1559 = (forvar1559 + (1'h1)))
                begin
                  if ((reg1480[(4'h9):(3'h6)] ?
                      $unsigned(reg1353[(1'h0):(1'h0)]) : reg1264))
                    begin
                      reg1560 <= $unsigned(((~|(reg1191 ? reg1160 : reg1312)) ?
                          $signed({(8'hb1)}) : {((8'ha3) || reg1378)}));
                      reg1561 <= reg1474[(4'he):(4'h8)];
                      reg1562 <= $unsigned((($signed(reg1525) & $unsigned(reg1272)) ?
                          $unsigned((|reg1214)) : $unsigned((reg1422 & reg1373))));
                      reg1563 <= reg1451[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1560 <= ((!{$unsigned(reg1327)}) << $unsigned(((reg1248 ?
                              (8'ha3) : (8'hb7)) ?
                          $unsigned(reg1278) : (~reg1179))));
                      reg1561 <= reg1444[(3'h4):(2'h3)];
                      reg1562 <= (reg1293 ?
                          (reg1220 ?
                              $signed($signed(reg1412)) : $unsigned((-reg1291))) : {({reg1262} ?
                                  reg1178 : ((8'h9d) ^~ reg1362))});
                    end
                end
              for (forvar1564 = (1'h0); (forvar1564 < (2'h3)); forvar1564 = (forvar1564 + (1'h1)))
                begin
                  for (forvar1565 = (1'h0); (forvar1565 < (1'h0)); forvar1565 = (forvar1565 + (1'h1)))
                    begin
                      reg1566 <= $unsigned(reg1482);
                    end
                  if ((~|$signed(reg1328[(3'h6):(1'h1)])))
                    begin
                      reg1567 <= reg1284;
                    end
                  else
                    begin
                      reg1567 <= ($unsigned(reg1173) ?
                          ((reg1260 ? (reg1399 | (8'ha2)) : wire1151) ?
                              ((reg1481 ?
                                  reg1531 : reg1383) + reg1511) : (8'hb2)) : $signed((8'had)));
                      reg1568 <= (-$signed(($signed(reg1405) >> {(8'had)})));
                      reg1569 <= ($signed(((&reg1525) ?
                          (~^wire1464) : (reg1442 ?
                              forvar1497 : reg1195))) <= ((+wire1159[(2'h2):(1'h1)]) ^ $unsigned(reg1196)));
                      reg1570 <= {{{$signed((8'hb1))}}};
                    end
                  for (forvar1571 = (1'h0); (forvar1571 < (1'h1)); forvar1571 = (forvar1571 + (1'h1)))
                    begin
                      reg1572 <= $unsigned(reg1550);
                      reg1573 <= ((!(~reg1389)) ?
                          ({$signed(forvar1546)} || (!reg1184[(1'h0):(1'h0)])) : $signed(($unsigned(reg1529) | ((8'ha2) ?
                              reg1548 : reg1347))));
                    end
                end
              for (forvar1574 = (1'h0); (forvar1574 < (2'h3)); forvar1574 = (forvar1574 + (1'h1)))
                begin
                  for (forvar1575 = (1'h0); (forvar1575 < (1'h1)); forvar1575 = (forvar1575 + (1'h1)))
                    begin
                      reg1576 <= $signed((((reg1371 ?
                              reg1473 : reg1411) || (reg1323 ^ reg1348)) ?
                          reg1523 : ((reg1440 ? reg1291 : (8'ha9)) ?
                              ((8'hba) ?
                                  wire1149 : reg1551) : reg1423[(3'h6):(3'h5)])));
                      reg1577 <= {reg1401};
                      reg1578 <= $signed(reg1316);
                      reg1579 <= $unsigned(reg1173[(3'h4):(2'h3)]);
                    end
                  for (forvar1580 = (1'h0); (forvar1580 < (1'h0)); forvar1580 = (forvar1580 + (1'h1)))
                    begin
                      reg1581 <= ((8'h9c) - reg1317[(3'h5):(3'h5)]);
                      reg1582 <= $signed($signed($signed((&reg1246))));
                    end
                  if ((|(reg1563 ?
                      $signed($unsigned(wire1150)) : {$unsigned(reg1221)})))
                    begin
                      reg1583 <= (((^(reg1222 <= reg1490)) - $unsigned((8'ha3))) << (|$signed(forvar1475[(3'h6):(2'h2)])));
                      reg1584 <= $signed(reg1483[(4'h9):(2'h2)]);
                      reg1585 <= (reg1428[(3'h5):(1'h0)] ?
                          reg1513[(2'h3):(2'h3)] : reg1518);
                    end
                  else
                    begin
                      reg1583 <= (8'ha1);
                      reg1584 <= (reg1359 * $signed((8'hb4)));
                      reg1585 <= reg1494;
                      reg1586 <= (((!$unsigned(forvar1549)) ?
                          reg1174 : reg1569) == reg1240);
                    end
                end
              for (forvar1587 = (1'h0); (forvar1587 < (2'h3)); forvar1587 = (forvar1587 + (1'h1)))
                begin
                  if ($signed($signed(({(8'h9c)} ?
                      reg1441[(3'h6):(3'h5)] : (reg1379 ? (8'ha3) : reg1191)))))
                    begin
                      reg1588 <= (~(reg1184[(4'h8):(2'h2)] ?
                          {(+reg1243)} : $signed(reg1197)));
                      reg1589 <= (&reg1332[(2'h2):(1'h0)]);
                      reg1590 <= (-({(reg1303 ^ reg1311)} < $signed((reg1328 ?
                          forvar1507 : (8'ha4)))));
                    end
                  else
                    begin
                      reg1588 <= $unsigned($unsigned($unsigned(reg1540)));
                      reg1589 <= (~|(+forvar1559[(3'h4):(3'h4)]));
                    end
                  for (forvar1591 = (1'h0); (forvar1591 < (2'h2)); forvar1591 = (forvar1591 + (1'h1)))
                    begin
                      reg1592 <= (^$signed($unsigned({reg1408})));
                      reg1593 <= $signed((($unsigned(reg1573) ~^ $unsigned(reg1472)) ?
                          $unsigned(reg1276[(2'h2):(1'h1)]) : reg1168[(1'h0):(1'h0)]));
                      reg1594 <= reg1570[(1'h1):(1'h1)];
                      reg1595 <= ($signed($unsigned((!(8'ha8)))) ?
                          (~&$signed(reg1405)) : reg1174);
                    end
                  for (forvar1596 = (1'h0); (forvar1596 < (2'h2)); forvar1596 = (forvar1596 + (1'h1)))
                    begin
                      reg1597 <= reg1338;
                      reg1598 <= ((reg1236[(2'h3):(1'h0)] ?
                          ((!reg1240) >>> forvar1580) : (-reg1252)) << reg1182[(3'h5):(3'h4)]);
                      reg1599 <= $unsigned((^(reg1293[(4'h9):(4'h8)] ?
                          $unsigned(reg1434) : (~&(8'ha4)))));
                      reg1600 <= (reg1599[(3'h6):(2'h3)] ?
                          $signed(((reg1592 >> (8'hb6)) ?
                              $unsigned(reg1383) : (reg1172 ~^ reg1233))) : reg1588[(1'h1):(1'h1)]);
                    end
                end
            end
          if ((8'hb2))
            begin
              for (forvar1601 = (1'h0); (forvar1601 < (1'h1)); forvar1601 = (forvar1601 + (1'h1)))
                begin
                  for (forvar1602 = (1'h0); (forvar1602 < (2'h3)); forvar1602 = (forvar1602 + (1'h1)))
                    begin
                      reg1603 <= {$unsigned((!reg1190[(3'h6):(2'h3)]))};
                      reg1604 <= $signed(((~^(reg1161 ^~ reg1527)) ?
                          ((reg1491 ?
                              forvar1549 : reg1512) <= reg1311) : (reg1284 ?
                              (reg1261 ? reg1340 : (8'haf)) : {reg1590})));
                    end
                end
            end
          else
            begin
              if ($unsigned((^~(-$unsigned(reg1313)))))
                begin
                  reg1601 <= reg1333;
                end
              else
                begin
                  for (forvar1601 = (1'h0); (forvar1601 < (1'h0)); forvar1601 = (forvar1601 + (1'h1)))
                    begin
                      reg1602 <= $unsigned((^($unsigned(reg1281) ?
                          (|(8'hb8)) : $signed(forvar1507))));
                    end
                  for (forvar1603 = (1'h0); (forvar1603 < (1'h1)); forvar1603 = (forvar1603 + (1'h1)))
                    begin
                      reg1604 <= $unsigned(((|$unsigned((8'h9c))) >> reg1431[(2'h2):(2'h2)]));
                      reg1605 <= reg1489[(3'h5):(1'h0)];
                      reg1606 <= ($signed((reg1262 ?
                              $signed(reg1547) : forvar1514[(3'h4):(3'h4)])) ?
                          ((reg1266[(1'h1):(1'h1)] ^~ $signed(reg1586)) << (reg1560[(1'h1):(1'h1)] ?
                              reg1261[(2'h2):(2'h2)] : reg1328[(1'h1):(1'h0)])) : $unsigned({{reg1206}}));
                      reg1607 <= ($signed($unsigned((reg1481 ?
                          reg1189 : (8'h9e)))) >= (~|$unsigned($signed(reg1225))));
                    end
                  if ((((~&$signed(reg1466)) >> reg1555) ?
                      {(reg1422 >> $unsigned(reg1508))} : wire1255[(1'h0):(1'h0)]))
                    begin
                      reg1608 <= ($signed({$unsigned(reg1266)}) ?
                          $unsigned($signed((^(8'h9c)))) : (reg1239[(1'h1):(1'h1)] ?
                              reg1188[(3'h4):(1'h1)] : reg1236[(4'ha):(4'h8)]));
                      reg1609 <= ((!reg1429) ?
                          $unsigned((reg1362[(4'hb):(1'h0)] ?
                              (&(8'ha5)) : reg1383)) : $signed({reg1224[(1'h1):(1'h1)]}));
                      reg1610 <= {(^~(((8'ha7) ? reg1251 : reg1607) ?
                              reg1417[(3'h6):(2'h3)] : reg1218))};
                      reg1611 <= $unsigned((!((wire1150 && reg1266) ?
                          ((8'hb1) ?
                              forvar1549 : reg1516) : reg1408[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg1608 <= $unsigned(($unsigned(reg1385) ?
                          forvar1465[(2'h3):(2'h3)] : (((8'ha0) < reg1185) ?
                              reg1229[(1'h1):(1'h0)] : (reg1518 ?
                                  reg1228 : reg1446))));
                      reg1609 <= $signed({$unsigned({reg1186})});
                      reg1610 <= reg1278[(3'h6):(1'h1)];
                    end
                  for (forvar1612 = (1'h0); (forvar1612 < (2'h3)); forvar1612 = (forvar1612 + (1'h1)))
                    begin
                      reg1613 <= reg1413[(1'h0):(1'h0)];
                      reg1614 <= {(-({forvar1558} + {reg1442}))};
                      reg1615 <= (reg1588[(1'h0):(1'h0)] <= forvar1575);
                      reg1616 <= $signed((reg1457 ?
                          {(&reg1253)} : $signed(reg1176)));
                    end
                end
              for (forvar1617 = (1'h0); (forvar1617 < (2'h3)); forvar1617 = (forvar1617 + (1'h1)))
                begin
                  reg1618 <= $unsigned(($unsigned(reg1537) & $unsigned(reg1606[(1'h0):(1'h0)])));
                  reg1619 <= wire1159;
                end
            end
        end
      else
        begin
          for (forvar1528 = (1'h0); (forvar1528 < (2'h3)); forvar1528 = (forvar1528 + (1'h1)))
            begin
              if ((~|$unsigned(reg1292)))
                begin
                  for (forvar1529 = (1'h0); (forvar1529 < (2'h3)); forvar1529 = (forvar1529 + (1'h1)))
                    begin
                      reg1530 <= $signed(((~^reg1288) ?
                          forvar1512[(3'h4):(1'h1)] : {reg1476}));
                      reg1531 <= reg1411;
                      reg1532 <= forvar1514[(3'h4):(1'h1)];
                      reg1533 <= $unsigned((~&(8'ha2)));
                    end
                  for (forvar1534 = (1'h0); (forvar1534 < (1'h0)); forvar1534 = (forvar1534 + (1'h1)))
                    begin
                      reg1535 <= $signed(($signed($unsigned(reg1166)) <= (((8'hab) <<< reg1382) ?
                          $unsigned((8'ha0)) : (~|(8'hab)))));
                      reg1536 <= ($unsigned({$unsigned(reg1432)}) * (reg1532 ?
                          {$unsigned(reg1323)} : reg1588));
                      reg1537 <= reg1619[(2'h2):(2'h2)];
                    end
                  for (forvar1538 = (1'h0); (forvar1538 < (1'h1)); forvar1538 = (forvar1538 + (1'h1)))
                    begin
                      reg1539 <= reg1193;
                      reg1540 <= {$signed(($unsigned(reg1326) ?
                              (~^reg1214) : reg1220[(4'hc):(4'hc)]))};
                    end
                  for (forvar1541 = (1'h0); (forvar1541 < (2'h3)); forvar1541 = (forvar1541 + (1'h1)))
                    begin
                      reg1542 <= reg1540;
                      reg1543 <= ($signed(($signed(reg1283) == $unsigned(reg1317))) ?
                          {(-reg1199[(2'h2):(1'h0)])} : $signed(({reg1476} ?
                              (reg1313 ? reg1265 : reg1371) : (reg1618 ?
                                  (8'ha7) : (8'haa)))));
                      reg1544 <= (~&(!((~&(8'hb6)) ?
                          reg1429[(1'h0):(1'h0)] : $signed(reg1164))));
                      reg1545 <= (|reg1273[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar1529 = (1'h0); (forvar1529 < (2'h3)); forvar1529 = (forvar1529 + (1'h1)))
                    begin
                      reg1530 <= (reg1189[(4'h9):(3'h4)] ?
                          ((-reg1171) ?
                              wire1150[(3'h5):(1'h1)] : $signed((reg1293 >> reg1311))) : ({$signed((8'hb9))} ?
                              reg1469[(3'h6):(3'h5)] : {(reg1252 >>> reg1430)}));
                      reg1531 <= reg1371;
                    end
                  if (((($signed(reg1523) >> reg1243) ?
                      reg1421[(3'h6):(3'h4)] : ($unsigned(forvar1564) <<< wire1151)) ^~ forvar1539))
                    begin
                      reg1532 <= $unsigned($signed($signed((^reg1183))));
                      reg1533 <= ((reg1478 ?
                          (|{reg1451}) : (!forvar1546)) ~^ reg1519[(3'h7):(3'h6)]);
                      reg1534 <= {reg1422[(3'h4):(2'h2)]};
                      reg1535 <= reg1578[(4'h8):(2'h3)];
                    end
                  else
                    begin
                      reg1532 <= ((({reg1332} ?
                              ((8'hb3) > reg1509) : (forvar1602 + reg1234)) * {(reg1260 >> reg1204)}) ?
                          (^(reg1570 ?
                              (reg1168 << reg1171) : $signed(reg1347))) : $signed(($unsigned(reg1606) > (reg1355 ?
                              reg1394 : reg1234))));
                      reg1533 <= $unsigned(reg1421);
                      reg1534 <= reg1274;
                      reg1535 <= (8'ha2);
                    end
                  for (forvar1536 = (1'h0); (forvar1536 < (1'h0)); forvar1536 = (forvar1536 + (1'h1)))
                    begin
                      reg1537 <= forvar1484;
                      reg1538 <= (~&$unsigned((~&(forvar1564 ?
                          forvar1612 : reg1517))));
                    end
                  reg1539 <= forvar1465[(1'h0):(1'h0)];
                end
              for (forvar1546 = (1'h0); (forvar1546 < (1'h1)); forvar1546 = (forvar1546 + (1'h1)))
                begin
                  for (forvar1547 = (1'h0); (forvar1547 < (2'h3)); forvar1547 = (forvar1547 + (1'h1)))
                    begin
                      reg1548 <= reg1601;
                      reg1549 <= $unsigned((((~(8'ha1)) ?
                          $unsigned(reg1445) : $signed(reg1371)) >> {{reg1507}}));
                    end
                end
            end
          if (reg1553[(1'h0):(1'h0)])
            begin
              for (forvar1550 = (1'h0); (forvar1550 < (1'h0)); forvar1550 = (forvar1550 + (1'h1)))
                begin
                  if (reg1300[(2'h2):(1'h0)])
                    begin
                      reg1551 <= $unsigned($unsigned(((reg1602 ^~ (8'h9c)) || reg1168)));
                    end
                  else
                    begin
                      reg1551 <= $signed((+forvar1564[(4'h8):(3'h4)]));
                      reg1552 <= $signed(($signed($signed((8'hb6))) != ((+reg1589) ?
                          reg1614 : ((8'hb8) <<< forvar1475))));
                      reg1553 <= reg1491[(3'h5):(3'h5)];
                    end
                end
              reg1554 <= ((8'hb3) ?
                  reg1291[(3'h5):(3'h4)] : (((reg1459 * reg1491) << (~&reg1225)) ?
                      {$unsigned(reg1171)} : {{reg1181}}));
              reg1555 <= reg1326;
            end
          else
            begin
              for (forvar1550 = (1'h0); (forvar1550 < (2'h2)); forvar1550 = (forvar1550 + (1'h1)))
                begin
                  reg1551 <= ({(!reg1488[(2'h2):(1'h1)])} | (reg1265 ?
                      reg1267[(1'h1):(1'h0)] : (~|(reg1524 ?
                          reg1288 : reg1184))));
                  for (forvar1552 = (1'h0); (forvar1552 < (2'h2)); forvar1552 = (forvar1552 + (1'h1)))
                    begin
                      reg1553 <= (($unsigned($signed(reg1277)) ?
                              ($signed(reg1553) ?
                                  forvar1549 : $unsigned(forvar1542)) : ($unsigned(reg1246) > $unsigned((8'hba)))) ?
                          (~&reg1477) : $unsigned($signed((reg1487 ?
                              reg1312 : reg1555))));
                      reg1554 <= (reg1614 >> reg1447);
                      reg1555 <= reg1444;
                      reg1556 <= (($unsigned($signed(reg1338)) ?
                          reg1308[(1'h1):(1'h1)] : reg1446[(2'h2):(1'h0)]) || $signed($unsigned((+(8'h9d)))));
                    end
                  for (forvar1557 = (1'h0); (forvar1557 < (2'h2)); forvar1557 = (forvar1557 + (1'h1)))
                    begin
                      reg1558 <= (($signed(reg1597) >= $signed(reg1264)) ?
                          (~^($signed(reg1189) || $unsigned(reg1177))) : ($unsigned((!reg1585)) ?
                              (reg1517 & forvar1534) : ($unsigned(reg1347) ?
                                  forvar1484 : reg1576[(1'h0):(1'h0)])));
                      reg1559 <= ({reg1404[(2'h3):(2'h2)]} && (~^((^reg1160) >= (reg1322 >>> reg1178))));
                      reg1560 <= $unsigned((^((!reg1214) ?
                          (reg1422 ? reg1339 : reg1429) : $unsigned(reg1160))));
                      reg1561 <= $signed(($unsigned(reg1529[(2'h2):(2'h2)]) ?
                          reg1284[(1'h0):(1'h0)] : $unsigned(reg1251)));
                    end
                end
              for (forvar1562 = (1'h0); (forvar1562 < (1'h1)); forvar1562 = (forvar1562 + (1'h1)))
                begin
                  for (forvar1563 = (1'h0); (forvar1563 < (2'h3)); forvar1563 = (forvar1563 + (1'h1)))
                    begin
                      reg1564 <= $signed(forvar1591);
                      reg1565 <= $signed((|(~^reg1609[(4'hf):(3'h5)])));
                      reg1566 <= ($unsigned($unsigned(reg1262)) != ($signed((^(8'hb0))) && $unsigned(((8'hb7) != reg1270))));
                    end
                end
            end
        end
      if ((-(^~$signed($unsigned(reg1453)))))
        begin
          for (forvar1620 = (1'h0); (forvar1620 < (2'h2)); forvar1620 = (forvar1620 + (1'h1)))
            begin
              for (forvar1621 = (1'h0); (forvar1621 < (1'h1)); forvar1621 = (forvar1621 + (1'h1)))
                begin
                  if ($unsigned((((reg1323 ^~ reg1396) << reg1442) ?
                      $unsigned((8'ha8)) : ($signed(forvar1574) & forvar1591[(3'h5):(1'h0)]))))
                    begin
                      reg1622 <= ($unsigned($unsigned(reg1213)) * reg1428[(3'h6):(1'h0)]);
                      reg1623 <= $signed(reg1413[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg1622 <= wire1157;
                      reg1623 <= ((^((~^reg1541) ?
                          reg1180[(4'ha):(4'ha)] : forvar1542)) >>> $unsigned(reg1538[(3'h7):(2'h3)]));
                    end
                end
            end
          reg1624 <= ($unsigned((wire1155[(4'hb):(4'hb)] ?
                  reg1606[(4'ha):(1'h1)] : (reg1456 ? reg1462 : reg1474))) ?
              reg1181[(3'h6):(2'h3)] : ($signed($signed(reg1178)) ?
                  (8'had) : forvar1484[(3'h4):(3'h4)]));
          for (forvar1625 = (1'h0); (forvar1625 < (2'h3)); forvar1625 = (forvar1625 + (1'h1)))
            begin
              for (forvar1626 = (1'h0); (forvar1626 < (1'h0)); forvar1626 = (forvar1626 + (1'h1)))
                begin
                  reg1627 <= $unsigned((8'hb2));
                  if ($signed((reg1281[(1'h1):(1'h1)] == $unsigned($unsigned(reg1327)))))
                    begin
                      reg1628 <= {reg1539[(4'hf):(3'h7)]};
                    end
                  else
                    begin
                      reg1628 <= reg1180[(2'h2):(2'h2)];
                      reg1629 <= $unsigned(reg1322);
                      reg1630 <= (($unsigned($signed(reg1508)) << ((reg1373 << reg1328) ?
                              reg1572[(1'h0):(1'h0)] : $signed(reg1229))) ?
                          reg1428[(4'h9):(1'h1)] : $unsigned($signed((reg1523 >>> reg1380))));
                    end
                  if ((~^((forvar1550 ? $unsigned(reg1267) : $signed(reg1627)) ?
                      {$signed(reg1399)} : (reg1177[(5'h10):(1'h1)] ?
                          reg1188[(2'h3):(2'h2)] : reg1517[(4'h9):(3'h5)]))))
                    begin
                      reg1631 <= $unsigned($unsigned(reg1529));
                      reg1632 <= $signed((((+reg1215) <<< (^reg1523)) << $signed(reg1489[(2'h2):(1'h1)])));
                    end
                  else
                    begin
                      reg1631 <= (-forvar1558);
                    end
                end
              if ((~^reg1477[(1'h1):(1'h0)]))
                begin
                  for (forvar1633 = (1'h0); (forvar1633 < (2'h3)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= (^~reg1417[(4'h8):(1'h1)]);
                    end
                  for (forvar1635 = (1'h0); (forvar1635 < (1'h0)); forvar1635 = (forvar1635 + (1'h1)))
                    begin
                      reg1636 <= (&((|reg1212[(3'h5):(2'h3)]) ?
                          wire1151[(1'h0):(1'h0)] : (reg1180[(4'hc):(1'h1)] || $unsigned(reg1344))));
                    end
                  for (forvar1637 = (1'h0); (forvar1637 < (2'h2)); forvar1637 = (forvar1637 + (1'h1)))
                    begin
                      reg1638 <= (^$signed(($signed(reg1486) ?
                          (reg1239 ?
                              reg1247 : reg1461) : (reg1379 ^~ reg1200))));
                      reg1639 <= (~($signed((^~(8'hb5))) << reg1477[(1'h0):(1'h0)]));
                      reg1640 <= $signed($unsigned($unsigned((reg1599 > reg1458))));
                    end
                end
              else
                begin
                  for (forvar1633 = (1'h0); (forvar1633 < (2'h2)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= reg1527;
                      reg1635 <= $signed(reg1453);
                      reg1636 <= ((reg1503 ?
                          (reg1339 ?
                              reg1375 : reg1219[(1'h0):(1'h0)]) : {$signed(reg1461)}) + $unsigned({reg1377[(3'h4):(3'h4)]}));
                    end
                  reg1637 <= {($signed(((8'h9d) ?
                          forvar1626 : (8'hb4))) + reg1479[(2'h2):(1'h1)])};
                  for (forvar1638 = (1'h0); (forvar1638 < (1'h1)); forvar1638 = (forvar1638 + (1'h1)))
                    begin
                      reg1639 <= ($unsigned($signed((reg1226 * reg1537))) ?
                          (reg1160[(1'h1):(1'h0)] * $unsigned((reg1410 ?
                              reg1536 : reg1351))) : reg1323);
                    end
                  for (forvar1640 = (1'h0); (forvar1640 < (1'h0)); forvar1640 = (forvar1640 + (1'h1)))
                    begin
                      reg1641 <= (|$signed($unsigned(reg1189)));
                      reg1642 <= $unsigned((~&(reg1389[(3'h6):(3'h6)] <<< {(8'h9f)})));
                      reg1643 <= ((reg1167 < $signed((~^forvar1503))) ?
                          $signed(reg1463) : {{((8'had) ? reg1453 : (8'hb3))}});
                    end
                end
              for (forvar1644 = (1'h0); (forvar1644 < (2'h3)); forvar1644 = (forvar1644 + (1'h1)))
                begin
                  reg1645 <= ($signed($signed($unsigned(forvar1545))) || (8'hba));
                  if (((($unsigned(reg1481) <= ((8'h9d) >= reg1360)) ^ (8'ha7)) ^ forvar1633))
                    begin
                      reg1646 <= $signed(({$signed(reg1333)} == reg1223));
                      reg1647 <= ($signed(forvar1575[(1'h1):(1'h1)]) ?
                          ($unsigned({reg1646}) ?
                              reg1358[(3'h4):(3'h4)] : ({(8'ha3)} ?
                                  {forvar1563} : (~^(8'hac)))) : $unsigned({(forvar1541 ?
                                  reg1289 : reg1536)}));
                    end
                  else
                    begin
                      reg1646 <= reg1373[(4'hf):(4'he)];
                      reg1647 <= reg1599;
                      reg1648 <= reg1518;
                      reg1649 <= (8'ha5);
                    end
                  if ($signed(reg1331))
                    begin
                      reg1650 <= (8'ha9);
                      reg1651 <= {((^~$unsigned(reg1266)) ?
                              reg1635 : ((reg1409 ^ reg1415) ?
                                  {reg1301} : (forvar1565 || (8'hb2))))};
                    end
                  else
                    begin
                      reg1650 <= reg1321[(1'h0):(1'h0)];
                      reg1651 <= (8'hb5);
                      reg1652 <= (~&{$unsigned($signed(reg1496))});
                    end
                  for (forvar1653 = (1'h0); (forvar1653 < (2'h2)); forvar1653 = (forvar1653 + (1'h1)))
                    begin
                      reg1654 <= (~^(8'h9c));
                    end
                end
            end
        end
      else
        begin
          for (forvar1620 = (1'h0); (forvar1620 < (2'h3)); forvar1620 = (forvar1620 + (1'h1)))
            begin
              for (forvar1621 = (1'h0); (forvar1621 < (1'h0)); forvar1621 = (forvar1621 + (1'h1)))
                begin
                  if ($unsigned(((reg1532[(2'h3):(2'h2)] * reg1611) ^ ($unsigned(reg1170) < reg1245[(3'h7):(1'h0)]))))
                    begin
                      reg1622 <= $signed((~$signed((~&reg1576))));
                      reg1623 <= (reg1227[(1'h0):(1'h0)] >> {reg1245[(4'ha):(2'h3)]});
                    end
                  else
                    begin
                      reg1622 <= reg1654[(4'h9):(2'h2)];
                    end
                  reg1624 <= ((8'ha3) ?
                      $unsigned(({reg1457} ?
                          $signed(reg1509) : (reg1639 * reg1160))) : (~$signed(reg1544)));
                  reg1625 <= reg1169;
                end
              if ($unsigned(reg1406[(1'h0):(1'h0)]))
                begin
                  if ($signed((-$unsigned($signed(reg1474)))))
                    begin
                      reg1626 <= (+reg1250);
                      reg1627 <= ((reg1213[(1'h0):(1'h0)] ?
                          (!$unsigned(reg1278)) : (|forvar1565[(2'h2):(1'h0)])) && (!(^reg1334[(4'he):(3'h5)])));
                      reg1628 <= reg1589[(4'he):(4'he)];
                    end
                  else
                    begin
                      reg1626 <= ($unsigned({reg1175[(3'h4):(2'h2)]}) >>> reg1605);
                    end
                  if (($signed($signed((reg1457 > forvar1621))) ?
                      reg1411[(1'h0):(1'h0)] : ($signed($unsigned(reg1166)) && reg1348[(3'h7):(1'h0)])))
                    begin
                      reg1629 <= forvar1475[(1'h0):(1'h0)];
                      reg1630 <= {$unsigned(((reg1190 ^~ reg1300) ?
                              $signed(reg1542) : reg1429))};
                      reg1631 <= (&reg1611[(4'hb):(3'h4)]);
                      reg1632 <= reg1188[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1629 <= $signed(reg1594[(1'h1):(1'h1)]);
                      reg1630 <= $signed((^reg1515));
                    end
                  if ($unsigned((reg1179[(3'h5):(1'h0)] ?
                      (~$unsigned(wire1464)) : ($signed(reg1409) && (~^reg1626)))))
                    begin
                      reg1633 <= ($unsigned(reg1611[(3'h4):(2'h2)]) & ((reg1431[(2'h3):(2'h3)] != (reg1543 ?
                          reg1473 : reg1504)) && reg1334[(4'h8):(3'h7)]));
                      reg1634 <= reg1508;
                      reg1635 <= $unsigned(reg1642);
                    end
                  else
                    begin
                      reg1633 <= $signed((&$unsigned($signed(reg1273))));
                      reg1634 <= {($unsigned((~|reg1400)) <= $signed(reg1640))};
                    end
                end
              else
                begin
                  reg1626 <= $signed(($signed(reg1223) ?
                      $unsigned($signed(reg1632)) : wire1151[(2'h2):(1'h1)]));
                  for (forvar1627 = (1'h0); (forvar1627 < (2'h2)); forvar1627 = (forvar1627 + (1'h1)))
                    begin
                      reg1628 <= forvar1471;
                      reg1629 <= ($unsigned(reg1181) || (!($unsigned((8'haa)) * $signed(reg1573))));
                    end
                end
              for (forvar1636 = (1'h0); (forvar1636 < (2'h2)); forvar1636 = (forvar1636 + (1'h1)))
                begin
                  for (forvar1637 = (1'h0); (forvar1637 < (1'h1)); forvar1637 = (forvar1637 + (1'h1)))
                    begin
                      reg1638 <= ({((~&reg1576) >= reg1473[(2'h2):(1'h0)])} ?
                          ($unsigned({(8'hb1)}) <<< $unsigned($signed(forvar1617))) : (~|$unsigned((+reg1466))));
                      reg1639 <= ($unsigned(reg1379) - $signed(($unsigned((8'hb3)) || reg1565[(1'h1):(1'h0)])));
                    end
                end
              reg1640 <= ((reg1412[(3'h6):(1'h0)] & forvar1546[(2'h2):(1'h0)]) ~^ forvar1617);
            end
        end
    end
  assign wire1655 = ((~|((reg1339 ? reg1289 : reg1225) ?
                        (~|reg1595) : reg1623)) >>> $unsigned(reg1347[(2'h3):(1'h0)]));
  assign wire1656 = {(reg1418[(1'h0):(1'h0)] != $signed(reg1601[(1'h1):(1'h0)]))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3045  (y, clk, wire3049, wire3048, wire3047, wire3046);
  output wire [(32'h14a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire3049;
  input wire [(4'ha):(1'h0)] wire3048;
  input wire signed [(4'h8):(1'h0)] wire3047;
  input wire signed [(3'h5):(1'h0)] wire3046;
  wire signed [(3'h4):(1'h0)] wire3416;
  wire signed [(2'h3):(1'h0)] wire3385;
  wire [(3'h7):(1'h0)] wire3055;
  wire signed [(4'hc):(1'h0)] wire3054;
  wire [(4'hc):(1'h0)] wire3053;
  wire [(4'he):(1'h0)] wire3052;
  wire [(3'h6):(1'h0)] wire3051;
  wire [(3'h4):(1'h0)] wire3050;
  reg [(2'h3):(1'h0)] reg3415 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3414 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3413 = (1'h0);
  reg [(4'h8):(1'h0)] reg3410 = (1'h0);
  reg [(5'h10):(1'h0)] reg3391 = (1'h0);
  reg [(3'h7):(1'h0)] reg3408 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3407 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3406 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3405 = (1'h0);
  reg [(2'h2):(1'h0)] reg3404 = (1'h0);
  reg [(4'hd):(1'h0)] reg3403 = (1'h0);
  reg [(4'hd):(1'h0)] reg3401 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3400 = (1'h0);
  reg [(2'h3):(1'h0)] reg3398 = (1'h0);
  reg [(4'he):(1'h0)] reg3396 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3395 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3394 = (1'h0);
  reg [(3'h4):(1'h0)] reg3393 = (1'h0);
  reg [(5'h10):(1'h0)] reg3392 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3389 = (1'h0);
  reg [(3'h7):(1'h0)] reg3388 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3412 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3411 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3409 = (1'h0);
  reg [(4'he):(1'h0)] forvar3402 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3399 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3397 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3391 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3390 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3387 = (1'h0);
  assign y = {wire3416,
                 wire3385,
                 wire3055,
                 wire3054,
                 wire3053,
                 wire3052,
                 wire3051,
                 wire3050,
                 reg3415,
                 reg3414,
                 reg3413,
                 reg3410,
                 reg3391,
                 reg3408,
                 reg3407,
                 reg3406,
                 reg3405,
                 reg3404,
                 reg3403,
                 reg3401,
                 reg3400,
                 reg3398,
                 reg3396,
                 reg3395,
                 reg3394,
                 reg3393,
                 reg3392,
                 reg3389,
                 reg3388,
                 forvar3412,
                 forvar3411,
                 forvar3409,
                 forvar3402,
                 forvar3399,
                 forvar3397,
                 forvar3391,
                 forvar3390,
                 forvar3387,
                 (1'h0)};
  assign wire3050 = wire3048;
  assign wire3051 = $signed((~(^wire3048[(3'h7):(1'h1)])));
  assign wire3052 = (wire3048 < wire3050);
  assign wire3053 = (!$unsigned((!(!wire3051))));
  assign wire3054 = (~|wire3048[(3'h4):(1'h1)]);
  assign wire3055 = $signed($signed(wire3051));
  module3056 #() modinst3386 (wire3385, clk, wire3052, wire3053, wire3054, wire3055);
  always
    @(posedge clk) begin
      for (forvar3387 = (1'h0); (forvar3387 < (1'h0)); forvar3387 = (forvar3387 + (1'h1)))
        begin
          reg3388 <= {({wire3047} ?
                  $signed(wire3052[(4'hc):(3'h7)]) : (|(~&wire3046)))};
          reg3389 <= $signed(wire3049[(4'h8):(3'h5)]);
          if (({$signed(wire3054)} ?
              wire3053 : (~$signed((wire3053 ? wire3052 : wire3047)))))
            begin
              for (forvar3390 = (1'h0); (forvar3390 < (1'h0)); forvar3390 = (forvar3390 + (1'h1)))
                begin
                  for (forvar3391 = (1'h0); (forvar3391 < (2'h2)); forvar3391 = (forvar3391 + (1'h1)))
                    begin
                      reg3392 <= wire3046[(2'h3):(2'h3)];
                      reg3393 <= wire3055;
                      reg3394 <= (({(forvar3387 ~^ (8'ha4))} ?
                              (~|$unsigned((8'ha3))) : {((8'haa) ?
                                      wire3052 : forvar3390)}) ?
                          {$signed(reg3392)} : ({wire3055} ?
                              {((8'hb8) && reg3388)} : wire3050[(2'h2):(1'h0)]));
                    end
                  if ($unsigned(((8'h9d) ?
                      $signed((~wire3054)) : (!$signed((8'hb1))))))
                    begin
                      reg3395 <= ($signed($unsigned($unsigned(reg3388))) ?
                          $signed(reg3393[(1'h0):(1'h0)]) : wire3052);
                    end
                  else
                    begin
                      reg3395 <= {$signed(wire3053[(2'h2):(2'h2)])};
                      reg3396 <= (~&(^(wire3385[(2'h3):(1'h0)] <= $signed(forvar3391))));
                    end
                end
              if ($signed($signed((&reg3389))))
                begin
                  for (forvar3397 = (1'h0); (forvar3397 < (1'h0)); forvar3397 = (forvar3397 + (1'h1)))
                    begin
                      reg3398 <= ($unsigned($signed((reg3388 + (8'hae)))) <<< $unsigned($unsigned(reg3394)));
                    end
                end
              else
                begin
                  for (forvar3397 = (1'h0); (forvar3397 < (1'h1)); forvar3397 = (forvar3397 + (1'h1)))
                    begin
                      reg3398 <= reg3388[(1'h0):(1'h0)];
                    end
                  for (forvar3399 = (1'h0); (forvar3399 < (1'h1)); forvar3399 = (forvar3399 + (1'h1)))
                    begin
                      reg3400 <= reg3392[(4'he):(4'h9)];
                      reg3401 <= (($signed($signed(wire3048)) <<< (((8'h9d) ?
                              reg3398 : reg3392) < (wire3047 << forvar3397))) ?
                          reg3393 : (^~{((8'hb7) <= (8'h9e))}));
                    end
                  for (forvar3402 = (1'h0); (forvar3402 < (1'h1)); forvar3402 = (forvar3402 + (1'h1)))
                    begin
                      reg3403 <= $signed(($signed(reg3396) ?
                          (~^$signed(forvar3402)) : $unsigned((~&reg3393))));
                      reg3404 <= reg3400;
                    end
                  if ({{$signed(wire3052[(3'h6):(2'h2)])}})
                    begin
                      reg3405 <= ({$signed(forvar3397[(1'h1):(1'h0)])} ?
                          (reg3396[(1'h0):(1'h0)] ?
                              reg3400 : wire3055[(1'h0):(1'h0)]) : reg3394);
                      reg3406 <= (8'haf);
                      reg3407 <= (-$signed(((wire3046 < forvar3402) ?
                          wire3051 : $unsigned(reg3405))));
                      reg3408 <= $unsigned(wire3051);
                    end
                  else
                    begin
                      reg3405 <= ((-((~reg3408) ?
                              $signed(wire3050) : reg3405)) ?
                          (~&((reg3406 ? reg3400 : (8'hb2)) ?
                              $unsigned(reg3405) : reg3406[(3'h4):(1'h1)])) : reg3395[(4'h8):(3'h5)]);
                      reg3406 <= $signed($unsigned(forvar3391));
                      reg3407 <= wire3048;
                    end
                end
            end
          else
            begin
              for (forvar3390 = (1'h0); (forvar3390 < (2'h2)); forvar3390 = (forvar3390 + (1'h1)))
                begin
                  if ((~|forvar3399))
                    begin
                      reg3391 <= $signed(($signed($signed(forvar3399)) ^~ ($unsigned(forvar3391) ^ (forvar3399 <= forvar3391))));
                    end
                  else
                    begin
                      reg3391 <= (8'hb3);
                      reg3392 <= {reg3400[(2'h3):(1'h0)]};
                      reg3393 <= ($unsigned($unsigned($signed(forvar3387))) | ({$signed(reg3403)} <<< ({reg3392} ?
                          reg3398[(1'h1):(1'h0)] : (reg3394 ?
                              reg3408 : wire3050))));
                      reg3394 <= reg3401;
                    end
                end
              reg3395 <= {($unsigned((forvar3402 ? wire3047 : wire3048)) ?
                      (wire3053[(3'h6):(3'h6)] ?
                          $unsigned((8'h9f)) : (wire3050 ?
                              forvar3390 : reg3393)) : $unsigned($signed(forvar3390)))};
            end
          for (forvar3409 = (1'h0); (forvar3409 < (2'h3)); forvar3409 = (forvar3409 + (1'h1)))
            begin
              reg3410 <= $signed(((|$signed(reg3396)) ?
                  forvar3409 : reg3403[(4'hd):(4'hc)]));
              for (forvar3411 = (1'h0); (forvar3411 < (1'h1)); forvar3411 = (forvar3411 + (1'h1)))
                begin
                  for (forvar3412 = (1'h0); (forvar3412 < (2'h3)); forvar3412 = (forvar3412 + (1'h1)))
                    begin
                      reg3413 <= (~{(8'ha7)});
                      reg3414 <= (~&$unsigned($unsigned((reg3396 ?
                          forvar3411 : reg3388))));
                    end
                end
            end
        end
      reg3415 <= $unsigned((!((forvar3412 ? reg3393 : reg3414) >= wire3050)));
    end
  assign wire3416 = $unsigned($unsigned(((reg3406 ? reg3405 : reg3403) ?
                        reg3394 : reg3401)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2039
#(parameter param3041 = {(((~|(8'hb2)) ? ((8'hae) ? (8'ha3) : (8'had)) : ((8'hb6) ? (8'hb1) : (8'hb1))) ? (~&(8'hb4)) : (((8'hb1) <<< (8'hb4)) != ((8'h9e) ? (8'ha2) : (8'hb8))))})
(y, clk, wire2044, wire2043, wire2042, wire2041, wire2040);
  output wire [(32'h1113):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire2044;
  input wire [(5'h10):(1'h0)] wire2043;
  input wire [(3'h4):(1'h0)] wire2042;
  input wire signed [(3'h7):(1'h0)] wire2041;
  input wire signed [(5'h10):(1'h0)] wire2040;
  wire signed [(4'hf):(1'h0)] wire3039;
  wire [(4'ha):(1'h0)] wire2578;
  wire signed [(4'ha):(1'h0)] wire2504;
  wire [(3'h6):(1'h0)] wire2502;
  wire signed [(3'h4):(1'h0)] wire2235;
  wire [(4'h8):(1'h0)] wire2234;
  reg signed [(5'h10):(1'h0)] reg2577 = (1'h0);
  reg [(3'h6):(1'h0)] reg2576 = (1'h0);
  reg [(5'h10):(1'h0)] reg2575 = (1'h0);
  reg [(4'hc):(1'h0)] reg2574 = (1'h0);
  reg [(2'h3):(1'h0)] reg2572 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2571 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2570 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2569 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2567 = (1'h0);
  reg [(3'h4):(1'h0)] reg2564 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2563 = (1'h0);
  reg [(4'hb):(1'h0)] reg2562 = (1'h0);
  reg [(4'ha):(1'h0)] reg2560 = (1'h0);
  reg [(2'h2):(1'h0)] reg2559 = (1'h0);
  reg [(3'h6):(1'h0)] reg2558 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2557 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2554 = (1'h0);
  reg [(4'ha):(1'h0)] reg2552 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2551 = (1'h0);
  reg [(4'h9):(1'h0)] reg2550 = (1'h0);
  reg [(4'hb):(1'h0)] reg2542 = (1'h0);
  reg [(3'h4):(1'h0)] reg2549 = (1'h0);
  reg [(3'h7):(1'h0)] reg2548 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2547 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2546 = (1'h0);
  reg [(2'h3):(1'h0)] reg2545 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2544 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2543 = (1'h0);
  reg [(2'h2):(1'h0)] reg2541 = (1'h0);
  reg [(4'hf):(1'h0)] reg2540 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2539 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2538 = (1'h0);
  reg [(2'h3):(1'h0)] reg2537 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2536 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2535 = (1'h0);
  reg [(2'h3):(1'h0)] reg2534 = (1'h0);
  reg [(4'h8):(1'h0)] reg2533 = (1'h0);
  reg [(3'h4):(1'h0)] reg2531 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2527 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2532 = (1'h0);
  reg [(5'h10):(1'h0)] reg2530 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2529 = (1'h0);
  reg [(2'h2):(1'h0)] reg2528 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2521 = (1'h0);
  reg [(3'h5):(1'h0)] reg2525 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2524 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2523 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2522 = (1'h0);
  reg [(4'h8):(1'h0)] reg2520 = (1'h0);
  reg [(3'h7):(1'h0)] reg2519 = (1'h0);
  reg [(2'h2):(1'h0)] reg2515 = (1'h0);
  reg [(4'he):(1'h0)] reg2518 = (1'h0);
  reg [(4'hb):(1'h0)] reg2517 = (1'h0);
  reg [(3'h5):(1'h0)] reg2514 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2513 = (1'h0);
  reg [(3'h7):(1'h0)] reg2512 = (1'h0);
  reg [(4'ha):(1'h0)] reg2510 = (1'h0);
  reg [(4'ha):(1'h0)] reg2509 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2508 = (1'h0);
  reg [(2'h3):(1'h0)] reg2507 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2048 = (1'h0);
  reg [(3'h4):(1'h0)] reg2050 = (1'h0);
  reg [(4'h9):(1'h0)] reg2051 = (1'h0);
  reg [(4'h9):(1'h0)] reg2052 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2046 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2047 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2049 = (1'h0);
  reg [(3'h5):(1'h0)] reg2053 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2054 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2055 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2056 = (1'h0);
  reg [(4'hc):(1'h0)] reg2057 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2059 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2060 = (1'h0);
  reg [(4'h9):(1'h0)] reg2061 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2064 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2065 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2066 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2067 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2069 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2071 = (1'h0);
  reg [(4'he):(1'h0)] reg2072 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2073 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2074 = (1'h0);
  reg [(2'h2):(1'h0)] reg2076 = (1'h0);
  reg [(4'hf):(1'h0)] reg2077 = (1'h0);
  reg [(4'hf):(1'h0)] reg2078 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2079 = (1'h0);
  reg [(3'h6):(1'h0)] reg2080 = (1'h0);
  reg [(4'hd):(1'h0)] reg2081 = (1'h0);
  reg [(2'h3):(1'h0)] reg2082 = (1'h0);
  reg [(4'hb):(1'h0)] reg2083 = (1'h0);
  reg [(4'ha):(1'h0)] reg2084 = (1'h0);
  reg [(2'h2):(1'h0)] reg2085 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2088 = (1'h0);
  reg [(4'h9):(1'h0)] reg2091 = (1'h0);
  reg [(3'h4):(1'h0)] reg2092 = (1'h0);
  reg [(4'he):(1'h0)] reg2093 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2094 = (1'h0);
  reg [(2'h2):(1'h0)] reg2096 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2098 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2099 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2100 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2101 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2102 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2103 = (1'h0);
  reg [(4'h9):(1'h0)] reg2104 = (1'h0);
  reg [(4'hf):(1'h0)] reg2106 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2107 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2108 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2109 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2095 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2097 = (1'h0);
  reg [(3'h5):(1'h0)] reg2110 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2114 = (1'h0);
  reg [(4'he):(1'h0)] reg2115 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2116 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2117 = (1'h0);
  reg [(3'h7):(1'h0)] reg2118 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2120 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2121 = (1'h0);
  reg [(3'h4):(1'h0)] reg2122 = (1'h0);
  reg [(4'hd):(1'h0)] reg2123 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2124 = (1'h0);
  reg [(3'h5):(1'h0)] reg2125 = (1'h0);
  reg [(3'h6):(1'h0)] reg2126 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2127 = (1'h0);
  reg [(4'hc):(1'h0)] reg2128 = (1'h0);
  reg [(4'hd):(1'h0)] reg2130 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2131 = (1'h0);
  reg [(4'he):(1'h0)] reg2132 = (1'h0);
  reg [(4'hf):(1'h0)] reg2129 = (1'h0);
  reg [(4'he):(1'h0)] reg2133 = (1'h0);
  reg [(4'he):(1'h0)] reg2134 = (1'h0);
  reg [(4'h9):(1'h0)] reg2112 = (1'h0);
  reg [(4'ha):(1'h0)] reg2113 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2119 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2137 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2140 = (1'h0);
  reg [(4'hc):(1'h0)] reg2141 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2142 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2143 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2144 = (1'h0);
  reg [(3'h5):(1'h0)] reg2145 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2146 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2148 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2149 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2150 = (1'h0);
  reg [(3'h4):(1'h0)] reg2152 = (1'h0);
  reg [(4'h9):(1'h0)] reg2153 = (1'h0);
  reg [(4'hb):(1'h0)] reg2154 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2155 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2156 = (1'h0);
  reg [(3'h5):(1'h0)] reg2147 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2151 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2159 = (1'h0);
  reg [(4'hd):(1'h0)] reg2160 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2161 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2162 = (1'h0);
  reg [(4'he):(1'h0)] reg2166 = (1'h0);
  reg [(4'ha):(1'h0)] reg2167 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2169 = (1'h0);
  reg [(4'hc):(1'h0)] reg2170 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2172 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2173 = (1'h0);
  reg [(4'hd):(1'h0)] reg2174 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2175 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2177 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2178 = (1'h0);
  reg [(4'hf):(1'h0)] reg2179 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2180 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2182 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2183 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2185 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2186 = (1'h0);
  reg [(4'he):(1'h0)] reg2187 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2188 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2189 = (1'h0);
  reg [(4'hf):(1'h0)] reg2190 = (1'h0);
  reg [(2'h2):(1'h0)] reg2191 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2193 = (1'h0);
  reg [(4'hc):(1'h0)] reg2194 = (1'h0);
  reg [(4'hc):(1'h0)] reg2195 = (1'h0);
  reg [(2'h2):(1'h0)] reg2197 = (1'h0);
  reg [(4'hd):(1'h0)] reg2198 = (1'h0);
  reg [(4'he):(1'h0)] reg2199 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2201 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2202 = (1'h0);
  reg [(4'hc):(1'h0)] reg2203 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2204 = (1'h0);
  reg [(4'h8):(1'h0)] reg2205 = (1'h0);
  reg [(3'h5):(1'h0)] reg2206 = (1'h0);
  reg [(4'he):(1'h0)] reg2210 = (1'h0);
  reg [(4'hf):(1'h0)] reg2211 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2212 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2213 = (1'h0);
  reg [(3'h6):(1'h0)] reg2214 = (1'h0);
  reg [(4'hd):(1'h0)] reg2215 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2216 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2217 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2218 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2209 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2222 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2223 = (1'h0);
  reg [(4'hb):(1'h0)] reg2224 = (1'h0);
  reg [(2'h3):(1'h0)] reg2226 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2227 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2228 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2229 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2230 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2231 = (1'h0);
  reg [(5'h10):(1'h0)] reg2232 = (1'h0);
  reg [(4'hc):(1'h0)] reg2233 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2238 = (1'h0);
  reg [(2'h2):(1'h0)] reg2239 = (1'h0);
  reg [(4'hc):(1'h0)] reg2240 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2241 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2242 = (1'h0);
  reg [(2'h3):(1'h0)] reg2243 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2244 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2246 = (1'h0);
  reg [(3'h5):(1'h0)] reg2247 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2248 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2249 = (1'h0);
  reg [(4'h8):(1'h0)] reg2250 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2251 = (1'h0);
  reg [(4'ha):(1'h0)] reg2253 = (1'h0);
  reg [(4'hf):(1'h0)] reg2252 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2255 = (1'h0);
  reg [(3'h5):(1'h0)] reg2257 = (1'h0);
  reg [(4'hf):(1'h0)] reg2258 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2259 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2260 = (1'h0);
  reg [(3'h6):(1'h0)] reg2261 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2263 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2264 = (1'h0);
  reg [(3'h5):(1'h0)] reg2266 = (1'h0);
  reg [(4'hb):(1'h0)] reg2267 = (1'h0);
  reg [(4'h8):(1'h0)] reg2262 = (1'h0);
  reg [(2'h2):(1'h0)] reg2265 = (1'h0);
  reg [(4'ha):(1'h0)] reg2268 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2269 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2271 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2272 = (1'h0);
  reg [(4'hf):(1'h0)] reg2273 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2275 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2276 = (1'h0);
  reg [(3'h6):(1'h0)] reg2277 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2278 = (1'h0);
  reg [(2'h3):(1'h0)] reg2279 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2280 = (1'h0);
  reg [(2'h2):(1'h0)] reg2281 = (1'h0);
  reg [(3'h4):(1'h0)] reg2282 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2270 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2274 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2284 = (1'h0);
  reg [(3'h6):(1'h0)] reg2285 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2286 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2287 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2289 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2290 = (1'h0);
  reg [(4'hd):(1'h0)] reg2293 = (1'h0);
  reg [(4'h9):(1'h0)] reg2294 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2295 = (1'h0);
  reg [(4'h9):(1'h0)] reg2296 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2299 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2300 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2301 = (1'h0);
  reg [(3'h7):(1'h0)] reg2303 = (1'h0);
  reg [(3'h6):(1'h0)] reg2304 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2305 = (1'h0);
  reg [(2'h2):(1'h0)] reg2306 = (1'h0);
  reg [(3'h6):(1'h0)] reg2307 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2302 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2288 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2291 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2297 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2298 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2309 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2310 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2311 = (1'h0);
  reg [(3'h6):(1'h0)] reg2313 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2314 = (1'h0);
  reg [(4'hf):(1'h0)] reg2315 = (1'h0);
  reg [(4'h9):(1'h0)] reg2316 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2245 = (1'h0);
  reg [(3'h7):(1'h0)] reg2254 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2256 = (1'h0);
  reg [(4'hb):(1'h0)] reg2237 = (1'h0);
  reg [(4'hb):(1'h0)] reg2283 = (1'h0);
  reg [(4'h8):(1'h0)] reg2292 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2312 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2308 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2319 = (1'h0);
  reg [(4'hf):(1'h0)] reg2320 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2322 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2323 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2324 = (1'h0);
  reg [(4'h9):(1'h0)] reg2327 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2328 = (1'h0);
  reg [(2'h3):(1'h0)] reg2329 = (1'h0);
  reg [(3'h6):(1'h0)] reg2331 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2333 = (1'h0);
  reg [(4'ha):(1'h0)] reg2334 = (1'h0);
  reg [(4'h8):(1'h0)] reg2335 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2336 = (1'h0);
  reg [(3'h5):(1'h0)] reg2337 = (1'h0);
  reg [(3'h6):(1'h0)] reg2339 = (1'h0);
  reg [(4'h8):(1'h0)] reg2340 = (1'h0);
  reg [(4'ha):(1'h0)] reg2343 = (1'h0);
  reg [(3'h7):(1'h0)] reg2345 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2346 = (1'h0);
  reg [(5'h10):(1'h0)] reg2347 = (1'h0);
  reg [(2'h2):(1'h0)] reg2348 = (1'h0);
  reg [(4'hd):(1'h0)] reg2349 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2350 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2351 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2352 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2354 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2355 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2356 = (1'h0);
  reg [(2'h3):(1'h0)] reg2357 = (1'h0);
  reg [(3'h7):(1'h0)] reg2358 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2359 = (1'h0);
  reg [(4'hc):(1'h0)] reg2360 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2361 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2362 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2365 = (1'h0);
  reg [(4'he):(1'h0)] reg2367 = (1'h0);
  reg [(2'h2):(1'h0)] reg2368 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2369 = (1'h0);
  reg [(2'h3):(1'h0)] reg2370 = (1'h0);
  reg [(4'hf):(1'h0)] reg2372 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2373 = (1'h0);
  reg [(4'he):(1'h0)] reg2374 = (1'h0);
  reg [(3'h5):(1'h0)] reg2375 = (1'h0);
  reg [(4'ha):(1'h0)] reg2376 = (1'h0);
  reg [(3'h7):(1'h0)] reg2377 = (1'h0);
  reg [(4'hb):(1'h0)] reg2378 = (1'h0);
  reg [(4'h9):(1'h0)] reg2379 = (1'h0);
  reg [(3'h5):(1'h0)] reg2381 = (1'h0);
  reg [(3'h4):(1'h0)] reg2382 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2383 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2384 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2385 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2386 = (1'h0);
  reg [(4'h9):(1'h0)] reg2387 = (1'h0);
  reg [(3'h7):(1'h0)] reg2388 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2389 = (1'h0);
  reg [(4'ha):(1'h0)] reg2391 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2392 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2573 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2568 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2566 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2565 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2561 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2556 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2555 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2553 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2549 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2547 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2539 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2528 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2542 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2531 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2527 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2526 = (1'h0);
  reg [(4'he):(1'h0)] forvar2521 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2514 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2512 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2516 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2515 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2511 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2506 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2505 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2390 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2381 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2380 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2371 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2366 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2364 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2363 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2353 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2344 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2342 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2341 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2338 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2332 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2330 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2326 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2325 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2319 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2321 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2318 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2317 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2306 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2304 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2295 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2281 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2280 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2273 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2269 = (1'h0);
  reg [(4'he):(1'h0)] forvar2266 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2241 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2260 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2255 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2248 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2242 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2309 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2312 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2308 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2301 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2290 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2285 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2303 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2302 = (1'h0);
  reg [(4'he):(1'h0)] forvar2298 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2297 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2292 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2291 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2288 = (1'h0);
  reg [(4'he):(1'h0)] forvar2283 = (1'h0);
  reg [(4'he):(1'h0)] forvar2274 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2270 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2264 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2265 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2262 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2256 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2254 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2249 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2252 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2245 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2237 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2236 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2228 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2225 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2221 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2220 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2219 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2212 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2210 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2209 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2208 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2207 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2200 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2190 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2186 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2196 = (1'h0);
  reg [(4'he):(1'h0)] forvar2192 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2184 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2181 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2176 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2171 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2168 = (1'h0);
  reg [(4'he):(1'h0)] forvar2165 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2164 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2163 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2158 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2157 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2152 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2149 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2151 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2147 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2139 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2138 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2136 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2135 = (1'h0);
  reg [(4'he):(1'h0)] forvar2115 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2131 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2125 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2129 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2119 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2113 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2112 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2111 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2096 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2105 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2097 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2095 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2090 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2089 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2087 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2086 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2075 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2070 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2068 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2063 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2062 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2058 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2051 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2049 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2047 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2046 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2045 = (1'h0);
  assign y = {wire3039,
                 wire2578,
                 wire2504,
                 wire2502,
                 wire2235,
                 wire2234,
                 reg2577,
                 reg2576,
                 reg2575,
                 reg2574,
                 reg2572,
                 reg2571,
                 reg2570,
                 reg2569,
                 reg2567,
                 reg2564,
                 reg2563,
                 reg2562,
                 reg2560,
                 reg2559,
                 reg2558,
                 reg2557,
                 reg2554,
                 reg2552,
                 reg2551,
                 reg2550,
                 reg2542,
                 reg2549,
                 reg2548,
                 reg2547,
                 reg2546,
                 reg2545,
                 reg2544,
                 reg2543,
                 reg2541,
                 reg2540,
                 reg2539,
                 reg2538,
                 reg2537,
                 reg2536,
                 reg2535,
                 reg2534,
                 reg2533,
                 reg2531,
                 reg2527,
                 reg2532,
                 reg2530,
                 reg2529,
                 reg2528,
                 reg2521,
                 reg2525,
                 reg2524,
                 reg2523,
                 reg2522,
                 reg2520,
                 reg2519,
                 reg2515,
                 reg2518,
                 reg2517,
                 reg2514,
                 reg2513,
                 reg2512,
                 reg2510,
                 reg2509,
                 reg2508,
                 reg2507,
                 reg2048,
                 reg2050,
                 reg2051,
                 reg2052,
                 reg2046,
                 reg2047,
                 reg2049,
                 reg2053,
                 reg2054,
                 reg2055,
                 reg2056,
                 reg2057,
                 reg2059,
                 reg2060,
                 reg2061,
                 reg2064,
                 reg2065,
                 reg2066,
                 reg2067,
                 reg2069,
                 reg2071,
                 reg2072,
                 reg2073,
                 reg2074,
                 reg2076,
                 reg2077,
                 reg2078,
                 reg2079,
                 reg2080,
                 reg2081,
                 reg2082,
                 reg2083,
                 reg2084,
                 reg2085,
                 reg2088,
                 reg2091,
                 reg2092,
                 reg2093,
                 reg2094,
                 reg2096,
                 reg2098,
                 reg2099,
                 reg2100,
                 reg2101,
                 reg2102,
                 reg2103,
                 reg2104,
                 reg2106,
                 reg2107,
                 reg2108,
                 reg2109,
                 reg2095,
                 reg2097,
                 reg2110,
                 reg2114,
                 reg2115,
                 reg2116,
                 reg2117,
                 reg2118,
                 reg2120,
                 reg2121,
                 reg2122,
                 reg2123,
                 reg2124,
                 reg2125,
                 reg2126,
                 reg2127,
                 reg2128,
                 reg2130,
                 reg2131,
                 reg2132,
                 reg2129,
                 reg2133,
                 reg2134,
                 reg2112,
                 reg2113,
                 reg2119,
                 reg2137,
                 reg2140,
                 reg2141,
                 reg2142,
                 reg2143,
                 reg2144,
                 reg2145,
                 reg2146,
                 reg2148,
                 reg2149,
                 reg2150,
                 reg2152,
                 reg2153,
                 reg2154,
                 reg2155,
                 reg2156,
                 reg2147,
                 reg2151,
                 reg2159,
                 reg2160,
                 reg2161,
                 reg2162,
                 reg2166,
                 reg2167,
                 reg2169,
                 reg2170,
                 reg2172,
                 reg2173,
                 reg2174,
                 reg2175,
                 reg2177,
                 reg2178,
                 reg2179,
                 reg2180,
                 reg2182,
                 reg2183,
                 reg2185,
                 reg2186,
                 reg2187,
                 reg2188,
                 reg2189,
                 reg2190,
                 reg2191,
                 reg2193,
                 reg2194,
                 reg2195,
                 reg2197,
                 reg2198,
                 reg2199,
                 reg2201,
                 reg2202,
                 reg2203,
                 reg2204,
                 reg2205,
                 reg2206,
                 reg2210,
                 reg2211,
                 reg2212,
                 reg2213,
                 reg2214,
                 reg2215,
                 reg2216,
                 reg2217,
                 reg2218,
                 reg2209,
                 reg2222,
                 reg2223,
                 reg2224,
                 reg2226,
                 reg2227,
                 reg2228,
                 reg2229,
                 reg2230,
                 reg2231,
                 reg2232,
                 reg2233,
                 reg2238,
                 reg2239,
                 reg2240,
                 reg2241,
                 reg2242,
                 reg2243,
                 reg2244,
                 reg2246,
                 reg2247,
                 reg2248,
                 reg2249,
                 reg2250,
                 reg2251,
                 reg2253,
                 reg2252,
                 reg2255,
                 reg2257,
                 reg2258,
                 reg2259,
                 reg2260,
                 reg2261,
                 reg2263,
                 reg2264,
                 reg2266,
                 reg2267,
                 reg2262,
                 reg2265,
                 reg2268,
                 reg2269,
                 reg2271,
                 reg2272,
                 reg2273,
                 reg2275,
                 reg2276,
                 reg2277,
                 reg2278,
                 reg2279,
                 reg2280,
                 reg2281,
                 reg2282,
                 reg2270,
                 reg2274,
                 reg2284,
                 reg2285,
                 reg2286,
                 reg2287,
                 reg2289,
                 reg2290,
                 reg2293,
                 reg2294,
                 reg2295,
                 reg2296,
                 reg2299,
                 reg2300,
                 reg2301,
                 reg2303,
                 reg2304,
                 reg2305,
                 reg2306,
                 reg2307,
                 reg2302,
                 reg2288,
                 reg2291,
                 reg2297,
                 reg2298,
                 reg2309,
                 reg2310,
                 reg2311,
                 reg2313,
                 reg2314,
                 reg2315,
                 reg2316,
                 reg2245,
                 reg2254,
                 reg2256,
                 reg2237,
                 reg2283,
                 reg2292,
                 reg2312,
                 reg2308,
                 reg2319,
                 reg2320,
                 reg2322,
                 reg2323,
                 reg2324,
                 reg2327,
                 reg2328,
                 reg2329,
                 reg2331,
                 reg2333,
                 reg2334,
                 reg2335,
                 reg2336,
                 reg2337,
                 reg2339,
                 reg2340,
                 reg2343,
                 reg2345,
                 reg2346,
                 reg2347,
                 reg2348,
                 reg2349,
                 reg2350,
                 reg2351,
                 reg2352,
                 reg2354,
                 reg2355,
                 reg2356,
                 reg2357,
                 reg2358,
                 reg2359,
                 reg2360,
                 reg2361,
                 reg2362,
                 reg2365,
                 reg2367,
                 reg2368,
                 reg2369,
                 reg2370,
                 reg2372,
                 reg2373,
                 reg2374,
                 reg2375,
                 reg2376,
                 reg2377,
                 reg2378,
                 reg2379,
                 reg2381,
                 reg2382,
                 reg2383,
                 reg2384,
                 reg2385,
                 reg2386,
                 reg2387,
                 reg2388,
                 reg2389,
                 reg2391,
                 reg2392,
                 forvar2573,
                 forvar2568,
                 forvar2566,
                 forvar2565,
                 forvar2561,
                 forvar2556,
                 forvar2555,
                 forvar2553,
                 forvar2549,
                 forvar2547,
                 forvar2539,
                 forvar2528,
                 forvar2542,
                 forvar2531,
                 forvar2527,
                 forvar2526,
                 forvar2521,
                 forvar2514,
                 forvar2512,
                 forvar2516,
                 forvar2515,
                 forvar2511,
                 forvar2506,
                 forvar2505,
                 forvar2390,
                 forvar2381,
                 forvar2380,
                 forvar2371,
                 forvar2366,
                 forvar2364,
                 forvar2363,
                 forvar2353,
                 forvar2344,
                 forvar2342,
                 forvar2341,
                 forvar2338,
                 forvar2332,
                 forvar2330,
                 forvar2326,
                 forvar2325,
                 forvar2319,
                 forvar2321,
                 forvar2318,
                 forvar2317,
                 forvar2306,
                 forvar2304,
                 forvar2295,
                 forvar2281,
                 forvar2280,
                 forvar2273,
                 forvar2269,
                 forvar2266,
                 forvar2241,
                 forvar2260,
                 forvar2255,
                 forvar2248,
                 forvar2242,
                 forvar2309,
                 forvar2312,
                 forvar2308,
                 forvar2301,
                 forvar2290,
                 forvar2285,
                 forvar2303,
                 forvar2302,
                 forvar2298,
                 forvar2297,
                 forvar2292,
                 forvar2291,
                 forvar2288,
                 forvar2283,
                 forvar2274,
                 forvar2270,
                 forvar2264,
                 forvar2265,
                 forvar2262,
                 forvar2256,
                 forvar2254,
                 forvar2249,
                 forvar2252,
                 forvar2245,
                 forvar2237,
                 forvar2236,
                 forvar2228,
                 forvar2225,
                 forvar2221,
                 forvar2220,
                 forvar2219,
                 forvar2212,
                 forvar2210,
                 forvar2209,
                 forvar2208,
                 forvar2207,
                 forvar2200,
                 forvar2190,
                 forvar2186,
                 forvar2196,
                 forvar2192,
                 forvar2184,
                 forvar2181,
                 forvar2176,
                 forvar2171,
                 forvar2168,
                 forvar2165,
                 forvar2164,
                 forvar2163,
                 forvar2158,
                 forvar2157,
                 forvar2152,
                 forvar2149,
                 forvar2151,
                 forvar2147,
                 forvar2139,
                 forvar2138,
                 forvar2136,
                 forvar2135,
                 forvar2115,
                 forvar2131,
                 forvar2125,
                 forvar2129,
                 forvar2119,
                 forvar2113,
                 forvar2112,
                 forvar2111,
                 forvar2096,
                 forvar2105,
                 forvar2097,
                 forvar2095,
                 forvar2090,
                 forvar2089,
                 forvar2087,
                 forvar2086,
                 forvar2075,
                 forvar2070,
                 forvar2068,
                 forvar2063,
                 forvar2062,
                 forvar2058,
                 forvar2051,
                 forvar2049,
                 forvar2047,
                 forvar2046,
                 forvar2045,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ({wire2042[(1'h1):(1'h0)]})
        begin
          for (forvar2045 = (1'h0); (forvar2045 < (2'h3)); forvar2045 = (forvar2045 + (1'h1)))
            begin
              for (forvar2046 = (1'h0); (forvar2046 < (2'h3)); forvar2046 = (forvar2046 + (1'h1)))
                begin
                  for (forvar2047 = (1'h0); (forvar2047 < (2'h2)); forvar2047 = (forvar2047 + (1'h1)))
                    begin
                      reg2048 <= ((^~wire2040[(3'h7):(2'h3)]) >= wire2041);
                    end
                  for (forvar2049 = (1'h0); (forvar2049 < (2'h2)); forvar2049 = (forvar2049 + (1'h1)))
                    begin
                      reg2050 <= wire2040;
                      reg2051 <= (wire2040[(2'h2):(2'h2)] ?
                          $signed(wire2044[(2'h3):(1'h1)]) : (reg2048[(3'h5):(1'h1)] != (8'hb7)));
                      reg2052 <= (((8'h9d) ?
                              forvar2047[(3'h5):(1'h1)] : $unsigned(reg2051[(2'h3):(1'h0)])) ?
                          ({{(8'ha7)}} ?
                              ({forvar2049} >= $unsigned(forvar2045)) : ($signed(forvar2045) ?
                                  (-wire2040) : $unsigned((8'hb3)))) : ($unsigned($unsigned(forvar2049)) <<< forvar2049));
                    end
                end
            end
        end
      else
        begin
          for (forvar2045 = (1'h0); (forvar2045 < (2'h3)); forvar2045 = (forvar2045 + (1'h1)))
            begin
              reg2046 <= (~($unsigned($unsigned(wire2044)) ?
                  (~|(forvar2046 ^~ wire2043)) : forvar2045[(3'h5):(2'h3)]));
              if (($unsigned($unsigned($signed(forvar2049))) ^ $signed(reg2048[(4'h8):(3'h6)])))
                begin
                  if (reg2046[(1'h0):(1'h0)])
                    begin
                      reg2047 <= wire2040[(4'hb):(4'hb)];
                      reg2048 <= {$unsigned(forvar2045)};
                      reg2049 <= $unsigned((~forvar2045));
                    end
                  else
                    begin
                      reg2047 <= {($signed(reg2048[(2'h2):(2'h2)]) ?
                              wire2044[(2'h2):(1'h0)] : wire2043)};
                      reg2048 <= $signed(wire2041[(3'h5):(1'h1)]);
                      reg2049 <= forvar2045[(3'h4):(3'h4)];
                    end
                end
              else
                begin
                  for (forvar2047 = (1'h0); (forvar2047 < (1'h1)); forvar2047 = (forvar2047 + (1'h1)))
                    begin
                      reg2048 <= ($unsigned((!(forvar2047 ?
                          wire2041 : reg2050))) <<< ((-(~reg2052)) > ($unsigned(forvar2045) < (reg2052 && forvar2045))));
                      reg2049 <= forvar2047[(2'h2):(1'h1)];
                      reg2050 <= (wire2043[(2'h2):(1'h0)] ?
                          (forvar2049[(2'h2):(2'h2)] ?
                              $unsigned(wire2043[(4'hf):(1'h0)]) : ((reg2048 >>> forvar2046) >= (~^forvar2045))) : $signed(wire2044[(1'h0):(1'h0)]));
                    end
                  for (forvar2051 = (1'h0); (forvar2051 < (1'h1)); forvar2051 = (forvar2051 + (1'h1)))
                    begin
                      reg2052 <= reg2048;
                      reg2053 <= (+reg2051[(3'h6):(3'h6)]);
                    end
                  if ((((!$signed(wire2044)) >>> wire2043[(4'h9):(4'h9)]) >> (((reg2052 && wire2043) << $signed(forvar2049)) << $unsigned(reg2050[(1'h0):(1'h0)]))))
                    begin
                      reg2054 <= wire2044;
                      reg2055 <= {{forvar2046[(3'h4):(3'h4)]}};
                      reg2056 <= $signed(forvar2046);
                    end
                  else
                    begin
                      reg2054 <= (!$unsigned($signed(reg2052)));
                      reg2055 <= (reg2052[(3'h4):(2'h2)] >>> reg2056[(4'hd):(1'h0)]);
                      reg2056 <= $signed((($unsigned(reg2054) ?
                              reg2049 : $signed(reg2046)) ?
                          reg2049 : (~&$signed((8'ha0)))));
                      reg2057 <= wire2044;
                    end
                end
              for (forvar2058 = (1'h0); (forvar2058 < (1'h1)); forvar2058 = (forvar2058 + (1'h1)))
                begin
                  reg2059 <= (~reg2049[(2'h2):(2'h2)]);
                  if (((^~((+reg2053) * $unsigned(reg2053))) << wire2043))
                    begin
                      reg2060 <= wire2044;
                      reg2061 <= $unsigned(($signed(reg2060) >> $signed((reg2055 ?
                          reg2047 : reg2059))));
                    end
                  else
                    begin
                      reg2060 <= reg2054[(4'hc):(4'hc)];
                    end
                end
            end
          for (forvar2062 = (1'h0); (forvar2062 < (2'h2)); forvar2062 = (forvar2062 + (1'h1)))
            begin
              for (forvar2063 = (1'h0); (forvar2063 < (2'h3)); forvar2063 = (forvar2063 + (1'h1)))
                begin
                  if ((forvar2049 ?
                      $unsigned(((8'ha2) >> {reg2053})) : (reg2046 >>> ((-reg2048) > (reg2056 && (8'ha0))))))
                    begin
                      reg2064 <= $signed(((!(^~reg2059)) >> ({forvar2046} ?
                          reg2050[(1'h1):(1'h1)] : (reg2047 ?
                              forvar2058 : (8'hb8)))));
                      reg2065 <= ((~^(reg2047 <= reg2056[(3'h6):(2'h2)])) <<< $unsigned(($unsigned(reg2047) ?
                          (reg2061 ? wire2042 : reg2049) : (^reg2048))));
                      reg2066 <= (|(^~((forvar2046 ? wire2040 : reg2059) ?
                          $signed(forvar2051) : $unsigned(reg2052))));
                      reg2067 <= (forvar2063 ?
                          reg2052[(1'h1):(1'h1)] : reg2050);
                    end
                  else
                    begin
                      reg2064 <= ((reg2060 ?
                          {(reg2057 ^ reg2059)} : ((forvar2062 * reg2046) >> (~reg2049))) - $signed($unsigned({forvar2063})));
                    end
                end
            end
          for (forvar2068 = (1'h0); (forvar2068 < (1'h0)); forvar2068 = (forvar2068 + (1'h1)))
            begin
              reg2069 <= ($signed((+$unsigned(reg2060))) ?
                  reg2047[(4'hb):(3'h5)] : forvar2068[(2'h2):(2'h2)]);
              for (forvar2070 = (1'h0); (forvar2070 < (2'h2)); forvar2070 = (forvar2070 + (1'h1)))
                begin
                  if ({((&(reg2067 * forvar2062)) ?
                          forvar2047 : (^forvar2049))})
                    begin
                      reg2071 <= forvar2062;
                      reg2072 <= $unsigned(({$signed(reg2059)} == reg2056[(4'h8):(1'h1)]));
                      reg2073 <= $signed($signed($signed((forvar2062 >>> reg2065))));
                      reg2074 <= (~|$unsigned((reg2059 <= reg2065)));
                    end
                  else
                    begin
                      reg2071 <= ($unsigned(forvar2062[(1'h0):(1'h0)]) - $unsigned(forvar2046[(2'h2):(1'h0)]));
                      reg2072 <= (reg2048 && ((~reg2061) < $unsigned((forvar2047 ?
                          forvar2046 : reg2071))));
                    end
                end
              for (forvar2075 = (1'h0); (forvar2075 < (1'h0)); forvar2075 = (forvar2075 + (1'h1)))
                begin
                  if ($signed((~^$unsigned($unsigned((8'hba))))))
                    begin
                      reg2076 <= forvar2068;
                      reg2077 <= reg2076;
                      reg2078 <= reg2049[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2076 <= (wire2040[(4'hc):(4'hc)] ?
                          ((+$signed(forvar2045)) - ({reg2047} ?
                              (~|reg2052) : {reg2067})) : $signed(($signed(reg2059) ?
                              (wire2040 >= reg2076) : $signed(forvar2062))));
                      reg2077 <= $signed(reg2077[(2'h3):(2'h2)]);
                    end
                  if ((reg2052[(3'h7):(2'h2)] ?
                      (forvar2068 ?
                          ((forvar2047 > forvar2063) ?
                              $signed(reg2049) : (reg2059 ?
                                  reg2053 : forvar2058)) : $unsigned(((8'haa) <<< wire2042))) : $unsigned((~|wire2041[(3'h6):(3'h5)]))))
                    begin
                      reg2079 <= {(~&reg2051)};
                      reg2080 <= (-$signed({reg2048}));
                      reg2081 <= $unsigned($unsigned((forvar2051 >> (reg2055 >> forvar2063))));
                    end
                  else
                    begin
                      reg2079 <= reg2053;
                      reg2080 <= (^((reg2061 ?
                              $unsigned(forvar2051) : $signed(reg2065)) ?
                          reg2055[(4'h9):(1'h0)] : $unsigned($unsigned(reg2049))));
                      reg2081 <= (!reg2081[(4'h9):(2'h3)]);
                    end
                  if ($signed((~&forvar2058[(4'hd):(2'h3)])))
                    begin
                      reg2082 <= ({(reg2057 ?
                              forvar2063 : $unsigned(reg2049))} <<< $signed($unsigned((reg2073 && forvar2058))));
                    end
                  else
                    begin
                      reg2082 <= reg2074;
                      reg2083 <= reg2056;
                      reg2084 <= ($signed(reg2055[(5'h10):(4'ha)]) ?
                          wire2043 : {($unsigned(reg2078) ?
                                  (8'ha7) : $signed(reg2060))});
                    end
                end
              reg2085 <= wire2044[(2'h3):(1'h0)];
            end
          for (forvar2086 = (1'h0); (forvar2086 < (2'h2)); forvar2086 = (forvar2086 + (1'h1)))
            begin
              for (forvar2087 = (1'h0); (forvar2087 < (2'h2)); forvar2087 = (forvar2087 + (1'h1)))
                begin
                  reg2088 <= ($signed(forvar2049) && $unsigned((&(|(8'h9f)))));
                end
              for (forvar2089 = (1'h0); (forvar2089 < (2'h3)); forvar2089 = (forvar2089 + (1'h1)))
                begin
                  for (forvar2090 = (1'h0); (forvar2090 < (2'h3)); forvar2090 = (forvar2090 + (1'h1)))
                    begin
                      reg2091 <= $unsigned(reg2047[(4'hf):(4'ha)]);
                      reg2092 <= (forvar2063 ?
                          wire2042 : $signed(((wire2043 ~^ (8'hb5)) ?
                              (~&reg2079) : (reg2064 > reg2071))));
                      reg2093 <= reg2049;
                      reg2094 <= ($unsigned(reg2083) ?
                          {($unsigned(reg2074) ?
                                  (reg2050 <<< forvar2062) : $signed(reg2054))} : (reg2093[(4'hb):(2'h3)] ?
                              (~(reg2083 ^ reg2046)) : $signed($unsigned(reg2081))));
                    end
                end
              if ((forvar2047 - $unsigned(wire2043)))
                begin
                  for (forvar2095 = (1'h0); (forvar2095 < (2'h3)); forvar2095 = (forvar2095 + (1'h1)))
                    begin
                      reg2096 <= ((-({(8'ha8)} >>> $unsigned(reg2080))) ?
                          (^~$signed(reg2082)) : reg2057[(1'h0):(1'h0)]);
                    end
                  for (forvar2097 = (1'h0); (forvar2097 < (1'h1)); forvar2097 = (forvar2097 + (1'h1)))
                    begin
                      reg2098 <= $unsigned({$signed(reg2074[(1'h1):(1'h0)])});
                      reg2099 <= $signed($unsigned($unsigned(reg2091[(1'h1):(1'h0)])));
                      reg2100 <= $unsigned(forvar2062);
                    end
                  if (reg2064)
                    begin
                      reg2101 <= (-wire2040);
                      reg2102 <= ($unsigned($unsigned($signed(reg2047))) >> reg2084);
                      reg2103 <= ((reg2096[(2'h2):(1'h0)] ?
                          $unsigned(reg2073) : forvar2068) + $unsigned($signed($signed(forvar2058))));
                      reg2104 <= (^~(~reg2051[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg2101 <= (+(forvar2070 ?
                          $signed((!wire2040)) : $unsigned($unsigned((8'ha3)))));
                      reg2102 <= $unsigned(reg2049[(2'h3):(1'h1)]);
                      reg2103 <= $unsigned((+(-reg2061)));
                      reg2104 <= (8'ha3);
                    end
                  for (forvar2105 = (1'h0); (forvar2105 < (2'h2)); forvar2105 = (forvar2105 + (1'h1)))
                    begin
                      reg2106 <= ((wire2044 ~^ $unsigned((reg2069 ?
                              reg2050 : (8'ha1)))) ?
                          (~^wire2043) : (&forvar2086));
                      reg2107 <= reg2053[(1'h1):(1'h0)];
                      reg2108 <= (~&$signed({$unsigned(wire2044)}));
                      reg2109 <= reg2080[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  reg2095 <= $signed(reg2107);
                  for (forvar2096 = (1'h0); (forvar2096 < (2'h3)); forvar2096 = (forvar2096 + (1'h1)))
                    begin
                      reg2097 <= reg2048[(3'h4):(2'h3)];
                      reg2098 <= $unsigned(($unsigned((+(8'hb8))) ?
                          ((forvar2095 ?
                              (8'hab) : reg2071) - $unsigned(forvar2087)) : reg2082));
                      reg2099 <= (reg2101 > $signed((reg2088 | wire2042)));
                      reg2100 <= $unsigned($unsigned(($signed((8'h9c)) ?
                          (~(8'hab)) : reg2064[(4'he):(1'h1)])));
                    end
                  reg2101 <= reg2103;
                end
              reg2110 <= reg2091[(3'h7):(1'h1)];
            end
        end
      for (forvar2111 = (1'h0); (forvar2111 < (1'h1)); forvar2111 = (forvar2111 + (1'h1)))
        begin
          if (($unsigned(((reg2104 ? reg2066 : reg2057) ?
              (reg2066 * wire2043) : $unsigned(reg2080))) <<< $unsigned({(reg2048 ?
                  forvar2051 : reg2101)})))
            begin
              for (forvar2112 = (1'h0); (forvar2112 < (1'h0)); forvar2112 = (forvar2112 + (1'h1)))
                begin
                  for (forvar2113 = (1'h0); (forvar2113 < (2'h2)); forvar2113 = (forvar2113 + (1'h1)))
                    begin
                      reg2114 <= {{(^(wire2041 ? (8'hac) : reg2096))}};
                      reg2115 <= $signed($signed(reg2056));
                      reg2116 <= $unsigned(forvar2113[(4'h8):(3'h7)]);
                      reg2117 <= (reg2074 ^~ ($signed($unsigned(forvar2062)) ?
                          $signed(reg2066[(2'h3):(2'h2)]) : reg2054));
                    end
                  reg2118 <= $unsigned((&forvar2090));
                  for (forvar2119 = (1'h0); (forvar2119 < (2'h3)); forvar2119 = (forvar2119 + (1'h1)))
                    begin
                      reg2120 <= (reg2109 ?
                          ((reg2060 - reg2046) ?
                              {(^(8'hb0))} : $unsigned({reg2097})) : ($unsigned(forvar2049) ?
                              reg2057 : reg2066));
                    end
                  if (($unsigned(reg2088) ?
                      {reg2050[(1'h0):(1'h0)]} : (forvar2049 ?
                          wire2040 : ((~&reg2101) ?
                              forvar2049[(4'h9):(2'h3)] : ((8'h9d) ?
                                  reg2110 : reg2109)))))
                    begin
                      reg2121 <= ($signed(wire2041) ?
                          $unsigned($signed((reg2054 ?
                              (8'hac) : (8'hb6)))) : ({reg2095} ?
                              $signed((forvar2058 ?
                                  forvar2113 : reg2120)) : ((&(8'hb7)) ?
                                  $signed(wire2041) : (reg2060 ?
                                      reg2076 : wire2043))));
                      reg2122 <= (($unsigned(forvar2070[(1'h1):(1'h0)]) ?
                              wire2043[(4'ha):(1'h1)] : (((8'ha6) << reg2115) == (+reg2072))) ?
                          (($unsigned(reg2065) ^~ (reg2050 * forvar2063)) ?
                              (|wire2044) : {reg2065[(3'h4):(3'h4)]}) : (8'haa));
                      reg2123 <= $signed((reg2096[(1'h1):(1'h0)] << (wire2044 + (forvar2049 | reg2065))));
                      reg2124 <= (^~reg2052);
                    end
                  else
                    begin
                      reg2121 <= forvar2062;
                    end
                end
              if ((reg2071 ?
                  (((+reg2122) * (~reg2051)) ?
                      $signed(reg2061[(4'h9):(2'h3)]) : (~^(-forvar2086))) : $unsigned({reg2055[(3'h4):(1'h0)]})))
                begin
                  if ((^$unsigned($unsigned(reg2121[(2'h2):(1'h0)]))))
                    begin
                      reg2125 <= ((&reg2102) >> $unsigned(reg2110));
                      reg2126 <= {({((8'hac) * forvar2097)} >> (|{(8'hb8)}))};
                      reg2127 <= $unsigned(((~&reg2047) ?
                          reg2103[(4'hb):(4'hb)] : reg2079));
                      reg2128 <= $unsigned($signed($signed($unsigned(reg2127))));
                    end
                  else
                    begin
                      reg2125 <= ((&(+reg2121)) ?
                          (forvar2090[(3'h5):(1'h1)] || (reg2118 ?
                              (reg2064 ?
                                  forvar2111 : (8'haf)) : $unsigned(reg2097))) : $signed(((8'hb3) || $signed(reg2078))));
                      reg2126 <= (($unsigned($unsigned(forvar2097)) == {$signed(forvar2068)}) && $unsigned(((-reg2064) >= $signed(reg2093))));
                    end
                  for (forvar2129 = (1'h0); (forvar2129 < (2'h3)); forvar2129 = (forvar2129 + (1'h1)))
                    begin
                      reg2130 <= forvar2113;
                      reg2131 <= {(reg2104 - wire2043)};
                      reg2132 <= reg2073[(2'h2):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar2125 = (1'h0); (forvar2125 < (1'h1)); forvar2125 = (forvar2125 + (1'h1)))
                    begin
                      reg2126 <= reg2115;
                      reg2127 <= (+(reg2117[(1'h0):(1'h0)] != reg2057[(3'h4):(3'h4)]));
                      reg2128 <= $signed((forvar2096[(3'h4):(3'h4)] ?
                          $signed($unsigned(reg2110)) : ((reg2096 <<< (8'hb4)) ?
                              (!reg2095) : $unsigned(reg2046))));
                      reg2129 <= (~|$unsigned(((reg2107 << reg2060) ?
                          (reg2072 ? reg2048 : reg2131) : forvar2058)));
                    end
                  reg2130 <= (wire2044 ?
                      {(~$signed(reg2059))} : forvar2051[(1'h0):(1'h0)]);
                  for (forvar2131 = (1'h0); (forvar2131 < (2'h2)); forvar2131 = (forvar2131 + (1'h1)))
                    begin
                      reg2132 <= {reg2085};
                      reg2133 <= (reg2057[(3'h6):(3'h4)] ?
                          (^~reg2127) : ($unsigned((~^(8'hba))) <<< ((reg2079 + reg2094) == (reg2103 ?
                              forvar2068 : reg2067))));
                    end
                  reg2134 <= reg2048;
                end
            end
          else
            begin
              if (((8'hac) ?
                  (^($signed(reg2101) ?
                      (reg2102 >>> (8'ha2)) : (forvar2068 ^ reg2081))) : ({(reg2091 >>> wire2044)} & wire2040)))
                begin
                  if (reg2082)
                    begin
                      reg2112 <= forvar2097;
                      reg2113 <= reg2084;
                      reg2114 <= $signed((((reg2117 ?
                              forvar2131 : reg2132) < $signed(reg2106)) ?
                          reg2056 : $signed((reg2127 ? (8'had) : (8'hb2)))));
                    end
                  else
                    begin
                      reg2112 <= $unsigned($signed({$unsigned(reg2106)}));
                    end
                  for (forvar2115 = (1'h0); (forvar2115 < (2'h3)); forvar2115 = (forvar2115 + (1'h1)))
                    begin
                      reg2116 <= (8'h9f);
                      reg2117 <= (^({(~reg2047)} > $signed((reg2061 ?
                          forvar2105 : reg2092))));
                      reg2118 <= ((($signed(forvar2047) > $signed(reg2061)) ?
                              (+{reg2132}) : reg2061[(1'h1):(1'h0)]) ?
                          ($unsigned(reg2123) | reg2121[(1'h0):(1'h0)]) : ({reg2095[(2'h3):(1'h1)]} ?
                              (+(reg2117 ?
                                  reg2133 : reg2129)) : (~|{reg2096})));
                      reg2119 <= reg2094[(1'h1):(1'h0)];
                    end
                  if ($signed($signed(forvar2113[(2'h2):(1'h1)])))
                    begin
                      reg2120 <= (((forvar2119 ?
                              $unsigned(reg2080) : (~reg2077)) ^ reg2082) ?
                          {$signed(reg2115[(4'hc):(2'h3)])} : reg2132[(3'h4):(2'h2)]);
                      reg2121 <= ((reg2110[(1'h0):(1'h0)] >> $signed((forvar2075 << reg2132))) ~^ {reg2130[(3'h6):(3'h6)]});
                    end
                  else
                    begin
                      reg2120 <= ((-forvar2096) > $signed(((reg2125 ?
                          forvar2089 : reg2054) >= $unsigned(reg2092))));
                      reg2121 <= reg2047;
                      reg2122 <= $signed($signed($signed($signed(forvar2063))));
                    end
                end
              else
                begin
                  if (reg2060)
                    begin
                      reg2112 <= $unsigned(reg2072);
                      reg2113 <= forvar2131[(3'h6):(2'h3)];
                    end
                  else
                    begin
                      reg2112 <= $signed($signed($signed(reg2107[(2'h3):(2'h2)])));
                      reg2113 <= (~|reg2099[(4'h9):(2'h3)]);
                      reg2114 <= ({{$unsigned((8'had))}} ^~ {$signed((forvar2115 >> reg2083))});
                    end
                  if ((8'h9c))
                    begin
                      reg2115 <= (~|(($signed(reg2117) ? (-reg2094) : reg2096) ?
                          reg2115[(2'h3):(2'h3)] : {(-(8'h9c))}));
                    end
                  else
                    begin
                      reg2115 <= ($signed($unsigned(reg2059)) ?
                          ((reg2128[(3'h6):(2'h3)] ? reg2128 : {reg2055}) ?
                              $unsigned($signed(forvar2131)) : ((~reg2114) ~^ (-(8'ha0)))) : reg2108);
                      reg2116 <= (~^((^(forvar2105 ? (8'hb9) : reg2096)) ?
                          reg2095[(4'ha):(4'ha)] : ((reg2093 ^~ (8'hb7)) - (8'hb3))));
                    end
                end
            end
        end
      for (forvar2135 = (1'h0); (forvar2135 < (2'h3)); forvar2135 = (forvar2135 + (1'h1)))
        begin
          for (forvar2136 = (1'h0); (forvar2136 < (1'h0)); forvar2136 = (forvar2136 + (1'h1)))
            begin
              reg2137 <= (^~(({reg2123} ?
                  reg2091[(3'h5):(1'h0)] : forvar2070[(2'h3):(2'h3)]) >> $unsigned(forvar2049[(3'h4):(1'h1)])));
              for (forvar2138 = (1'h0); (forvar2138 < (2'h3)); forvar2138 = (forvar2138 + (1'h1)))
                begin
                  for (forvar2139 = (1'h0); (forvar2139 < (1'h0)); forvar2139 = (forvar2139 + (1'h1)))
                    begin
                      reg2140 <= {(reg2080[(2'h2):(2'h2)] >> ({reg2122} << (~|forvar2113)))};
                      reg2141 <= reg2110;
                      reg2142 <= $signed($signed(forvar2135));
                    end
                  if ($unsigned({reg2132}))
                    begin
                      reg2143 <= reg2055;
                      reg2144 <= {reg2059[(4'hb):(4'h9)]};
                      reg2145 <= reg2095[(3'h5):(3'h5)];
                      reg2146 <= (-$signed(forvar2046));
                    end
                  else
                    begin
                      reg2143 <= forvar2139[(3'h7):(3'h7)];
                      reg2144 <= ($signed(forvar2045[(3'h5):(1'h1)]) ?
                          reg2076 : ((-(reg2146 >> wire2041)) >= ($unsigned(reg2092) ?
                              reg2074 : ((8'ha4) ? reg2098 : reg2125))));
                      reg2145 <= $unsigned((~|$unsigned((8'ha7))));
                    end
                end
            end
          if ((~&$signed((!forvar2095[(3'h7):(2'h2)]))))
            begin
              if (({(!(reg2088 ? reg2140 : reg2064))} ?
                  reg2142[(4'hc):(4'ha)] : $unsigned(reg2120[(1'h0):(1'h0)])))
                begin
                  for (forvar2147 = (1'h0); (forvar2147 < (2'h3)); forvar2147 = (forvar2147 + (1'h1)))
                    begin
                      reg2148 <= forvar2129;
                      reg2149 <= wire2044[(2'h3):(2'h2)];
                      reg2150 <= ($signed($signed(reg2146)) ?
                          $signed(reg2129[(4'h9):(3'h5)]) : $signed(($unsigned(reg2127) ?
                              (8'hb3) : $unsigned(reg2076))));
                    end
                  for (forvar2151 = (1'h0); (forvar2151 < (1'h1)); forvar2151 = (forvar2151 + (1'h1)))
                    begin
                      reg2152 <= reg2076;
                      reg2153 <= $unsigned($unsigned(reg2106));
                    end
                  if (($unsigned(reg2096) || (-reg2144[(3'h5):(3'h4)])))
                    begin
                      reg2154 <= ($unsigned($unsigned(reg2121[(1'h1):(1'h0)])) <<< reg2099[(3'h7):(2'h3)]);
                      reg2155 <= reg2148[(1'h1):(1'h1)];
                      reg2156 <= (forvar2136[(3'h5):(3'h5)] ?
                          $signed(reg2078) : forvar2147);
                    end
                  else
                    begin
                      reg2154 <= (({(^forvar2049)} ?
                          ((!reg2148) & (reg2108 ?
                              reg2064 : forvar2139)) : (+$unsigned((8'hb8)))) && reg2145);
                      reg2155 <= reg2093;
                      reg2156 <= forvar2105;
                    end
                end
              else
                begin
                  reg2147 <= $signed($unsigned((~&reg2102[(3'h4):(2'h3)])));
                  reg2148 <= reg2059;
                  for (forvar2149 = (1'h0); (forvar2149 < (2'h2)); forvar2149 = (forvar2149 + (1'h1)))
                    begin
                      reg2150 <= {$unsigned(((reg2077 ? reg2110 : reg2078) ?
                              (reg2067 * reg2096) : reg2108[(1'h0):(1'h0)]))};
                      reg2151 <= (~{(&$signed(reg2053))});
                    end
                  for (forvar2152 = (1'h0); (forvar2152 < (2'h2)); forvar2152 = (forvar2152 + (1'h1)))
                    begin
                      reg2153 <= {forvar2086[(3'h7):(3'h5)]};
                      reg2154 <= (reg2093 > ($unsigned(reg2149) != ((~^reg2155) ?
                          {reg2123} : (forvar2111 ? reg2130 : (8'h9f)))));
                      reg2155 <= (~^$signed({(reg2116 >= forvar2062)}));
                      reg2156 <= (($unsigned(wire2044) ?
                              ((!reg2073) ^ (|reg2098)) : ({reg2142} ?
                                  $unsigned(reg2102) : $signed(reg2141))) ?
                          {$unsigned((reg2080 > reg2123))} : {$signed(reg2143)});
                    end
                end
              for (forvar2157 = (1'h0); (forvar2157 < (2'h2)); forvar2157 = (forvar2157 + (1'h1)))
                begin
                  for (forvar2158 = (1'h0); (forvar2158 < (1'h0)); forvar2158 = (forvar2158 + (1'h1)))
                    begin
                      reg2159 <= $unsigned((((!reg2131) ?
                          forvar2151 : forvar2136) | {reg2100[(4'h8):(1'h1)]}));
                      reg2160 <= reg2047[(4'h8):(4'h8)];
                      reg2161 <= (((forvar2119[(3'h6):(2'h3)] ^~ $signed(forvar2086)) ?
                              reg2093[(1'h0):(1'h0)] : ({reg2076} ~^ forvar2149)) ?
                          {$signed({(8'h9f)})} : ($signed($signed(reg2054)) >= reg2125[(2'h2):(2'h2)]));
                    end
                end
            end
          else
            begin
              reg2147 <= reg2079[(3'h7):(1'h0)];
            end
          reg2162 <= forvar2151;
          for (forvar2163 = (1'h0); (forvar2163 < (2'h3)); forvar2163 = (forvar2163 + (1'h1)))
            begin
              for (forvar2164 = (1'h0); (forvar2164 < (1'h0)); forvar2164 = (forvar2164 + (1'h1)))
                begin
                  for (forvar2165 = (1'h0); (forvar2165 < (2'h2)); forvar2165 = (forvar2165 + (1'h1)))
                    begin
                      reg2166 <= $unsigned(forvar2063);
                    end
                  reg2167 <= {$signed(((8'ha7) > forvar2138[(1'h1):(1'h0)]))};
                  for (forvar2168 = (1'h0); (forvar2168 < (2'h3)); forvar2168 = (forvar2168 + (1'h1)))
                    begin
                      reg2169 <= ((reg2053 ?
                          (forvar2149 ?
                              {reg2127} : $signed(forvar2068)) : ((forvar2164 <= reg2153) | (reg2128 >> reg2066))) << (reg2103[(3'h6):(1'h0)] >> $signed(reg2069[(3'h7):(2'h2)])));
                      reg2170 <= $signed((^reg2108[(2'h2):(1'h0)]));
                    end
                  for (forvar2171 = (1'h0); (forvar2171 < (2'h3)); forvar2171 = (forvar2171 + (1'h1)))
                    begin
                      reg2172 <= $unsigned((-((reg2094 ? reg2052 : forvar2047) ?
                          {reg2048} : (~|forvar2139))));
                      reg2173 <= (~&(reg2142 <<< ($signed((8'ha7)) ^~ {reg2102})));
                      reg2174 <= (&(^(reg2137 >> forvar2089[(1'h1):(1'h1)])));
                      reg2175 <= forvar2136;
                    end
                end
              if ($unsigned({(-(~&(8'hba)))}))
                begin
                  for (forvar2176 = (1'h0); (forvar2176 < (2'h3)); forvar2176 = (forvar2176 + (1'h1)))
                    begin
                      reg2177 <= {{$signed(forvar2138[(1'h1):(1'h0)])}};
                      reg2178 <= (!(($unsigned(reg2095) ?
                          (forvar2158 ?
                              forvar2129 : forvar2147) : {wire2041}) >>> reg2177));
                    end
                end
              else
                begin
                  for (forvar2176 = (1'h0); (forvar2176 < (1'h1)); forvar2176 = (forvar2176 + (1'h1)))
                    begin
                      reg2177 <= reg2112[(1'h1):(1'h1)];
                      reg2178 <= ($signed(reg2133) ?
                          reg2092 : (~&$unsigned((reg2149 ^~ reg2145))));
                      reg2179 <= ($signed(($unsigned(forvar2090) || (&forvar2063))) ?
                          $signed(forvar2070[(2'h2):(1'h1)]) : (($signed(reg2066) ?
                              $unsigned(reg2159) : (forvar2151 << forvar2135)) >= {$signed((8'ha3))}));
                      reg2180 <= (|$unsigned($unsigned({reg2162})));
                    end
                  for (forvar2181 = (1'h0); (forvar2181 < (2'h2)); forvar2181 = (forvar2181 + (1'h1)))
                    begin
                      reg2182 <= reg2120;
                      reg2183 <= (reg2052[(3'h4):(1'h0)] ?
                          $signed(((8'hab) ?
                              reg2095 : reg2149)) : ($signed($signed(reg2052)) ?
                              (reg2172 ?
                                  $signed(reg2117) : (!reg2124)) : ((reg2091 ?
                                  reg2103 : (8'ha2)) * forvar2051[(1'h1):(1'h0)])));
                    end
                end
              if (reg2126)
                begin
                  for (forvar2184 = (1'h0); (forvar2184 < (2'h3)); forvar2184 = (forvar2184 + (1'h1)))
                    begin
                      reg2185 <= ($signed(($unsigned(reg2060) ?
                          (reg2064 >= reg2082) : $unsigned(forvar2125))) * $signed($signed(reg2117)));
                      reg2186 <= reg2100[(4'hd):(1'h0)];
                      reg2187 <= {reg2151[(2'h2):(2'h2)]};
                      reg2188 <= $signed(reg2085[(2'h2):(1'h1)]);
                    end
                  if ($unsigned(reg2073[(3'h7):(3'h6)]))
                    begin
                      reg2189 <= ($signed((reg2118 | (~^reg2178))) ?
                          $unsigned(forvar2063[(1'h1):(1'h0)]) : $signed(((reg2125 != reg2049) ?
                              (forvar2111 ?
                                  reg2056 : reg2079) : $unsigned(reg2182))));
                      reg2190 <= $signed($signed(reg2134));
                    end
                  else
                    begin
                      reg2189 <= ($unsigned(forvar2089) >= reg2190);
                      reg2190 <= $unsigned((reg2190[(1'h0):(1'h0)] && reg2148));
                      reg2191 <= (forvar2089[(3'h5):(3'h4)] ?
                          (8'hb5) : forvar2058);
                    end
                  for (forvar2192 = (1'h0); (forvar2192 < (1'h1)); forvar2192 = (forvar2192 + (1'h1)))
                    begin
                      reg2193 <= reg2071;
                      reg2194 <= (forvar2096[(1'h0):(1'h0)] <= reg2066);
                      reg2195 <= (~reg2140[(2'h2):(2'h2)]);
                    end
                  for (forvar2196 = (1'h0); (forvar2196 < (2'h2)); forvar2196 = (forvar2196 + (1'h1)))
                    begin
                      reg2197 <= ($signed((~$unsigned(reg2057))) ^~ (reg2101 ?
                          $signed((^reg2122)) : (forvar2135[(4'h9):(3'h7)] ?
                              $unsigned((8'hba)) : (~reg2167))));
                      reg2198 <= (reg2194[(1'h1):(1'h0)] ?
                          $unsigned($unsigned($signed((8'hb1)))) : (&({reg2078} + {reg2069})));
                      reg2199 <= (|$signed(forvar2051));
                    end
                end
              else
                begin
                  for (forvar2184 = (1'h0); (forvar2184 < (2'h2)); forvar2184 = (forvar2184 + (1'h1)))
                    begin
                      reg2185 <= ($unsigned(forvar2138[(3'h4):(1'h0)]) ?
                          $signed(($unsigned(forvar2136) || $signed(reg2048))) : forvar2095[(1'h1):(1'h0)]);
                    end
                  for (forvar2186 = (1'h0); (forvar2186 < (2'h3)); forvar2186 = (forvar2186 + (1'h1)))
                    begin
                      reg2187 <= $signed((+$unsigned($signed(reg2092))));
                      reg2188 <= ({$signed({forvar2068})} & (8'ha2));
                      reg2189 <= (!((~^(forvar2164 >= reg2114)) ?
                          ($unsigned((8'ha5)) > (forvar2058 ^ (8'ha1))) : reg2060));
                    end
                  for (forvar2190 = (1'h0); (forvar2190 < (1'h1)); forvar2190 = (forvar2190 + (1'h1)))
                    begin
                      reg2191 <= $unsigned(reg2188[(3'h5):(2'h2)]);
                    end
                end
              for (forvar2200 = (1'h0); (forvar2200 < (1'h1)); forvar2200 = (forvar2200 + (1'h1)))
                begin
                  if (((($unsigned(reg2142) ~^ (~&forvar2135)) ?
                      reg2185 : ((^(8'hb7)) ? reg2107 : reg2085)) & (8'hb6)))
                    begin
                      reg2201 <= forvar2200[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2201 <= $signed(forvar2090);
                      reg2202 <= forvar2105;
                    end
                  if (($unsigned((+(!reg2117))) <<< $unsigned($unsigned($signed((8'ha6))))))
                    begin
                      reg2203 <= reg2121;
                      reg2204 <= (($signed($signed(forvar2090)) ?
                              {$unsigned(reg2056)} : reg2170[(3'h5):(1'h1)]) ?
                          (8'hb4) : (8'ha6));
                      reg2205 <= reg2154;
                      reg2206 <= $unsigned(forvar2086);
                    end
                  else
                    begin
                      reg2203 <= $unsigned(((~|$signed(forvar2151)) && $signed(wire2042)));
                      reg2204 <= reg2197[(1'h0):(1'h0)];
                      reg2205 <= reg2114[(4'h9):(3'h5)];
                    end
                end
            end
        end
      for (forvar2207 = (1'h0); (forvar2207 < (2'h3)); forvar2207 = (forvar2207 + (1'h1)))
        begin
          for (forvar2208 = (1'h0); (forvar2208 < (2'h3)); forvar2208 = (forvar2208 + (1'h1)))
            begin
              if (($signed(reg2110[(3'h4):(2'h3)]) << (-$unsigned(((8'hb7) ?
                  reg2143 : (8'ha1))))))
                begin
                  for (forvar2209 = (1'h0); (forvar2209 < (1'h1)); forvar2209 = (forvar2209 + (1'h1)))
                    begin
                      reg2210 <= $unsigned((reg2162 ?
                          $signed({reg2132}) : $signed($unsigned(forvar2190))));
                      reg2211 <= (8'h9c);
                    end
                  if (((|($signed(reg2193) ? reg2074 : reg2076)) ?
                      reg2107 : (~(8'ha2))))
                    begin
                      reg2212 <= (~(reg2054 > $unsigned($signed((8'ha8)))));
                      reg2213 <= forvar2138;
                    end
                  else
                    begin
                      reg2212 <= $unsigned(($signed($unsigned(reg2059)) < ((&reg2177) ?
                          {(8'hb8)} : $unsigned(forvar2086))));
                      reg2213 <= reg2166;
                      reg2214 <= (~reg2121[(1'h1):(1'h0)]);
                      reg2215 <= (8'ha0);
                    end
                  if ((^~($signed($signed(forvar2068)) ?
                      (^~(forvar2115 ^ reg2102)) : {((8'hab) ?
                              reg2115 : (8'hb7))})))
                    begin
                      reg2216 <= $unsigned($unsigned((^~reg2130[(1'h1):(1'h1)])));
                      reg2217 <= ($unsigned($unsigned($unsigned(reg2098))) >= ({reg2188} - reg2199[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg2216 <= $signed((8'ha6));
                      reg2217 <= (&((~|(reg2124 ? reg2099 : (8'hb5))) ?
                          $signed((forvar2151 ?
                              reg2166 : forvar2135)) : (reg2130[(4'hb):(4'ha)] ^ (reg2191 ?
                              (8'haa) : (8'ha3)))));
                      reg2218 <= $unsigned($unsigned(({(8'hb5)} << {reg2201})));
                    end
                end
              else
                begin
                  reg2209 <= reg2113[(3'h6):(1'h1)];
                  for (forvar2210 = (1'h0); (forvar2210 < (2'h3)); forvar2210 = (forvar2210 + (1'h1)))
                    begin
                      reg2211 <= $signed((reg2170[(2'h2):(1'h1)] ?
                          (8'hb8) : ((reg2214 ? reg2194 : (8'haf)) ?
                              reg2073[(5'h10):(5'h10)] : wire2042)));
                    end
                  for (forvar2212 = (1'h0); (forvar2212 < (2'h3)); forvar2212 = (forvar2212 + (1'h1)))
                    begin
                      reg2213 <= (($unsigned(forvar2135) ?
                              (reg2049 ?
                                  ((8'ha8) ?
                                      reg2084 : reg2182) : (~^(8'ha1))) : reg2191) ?
                          $unsigned($signed($signed(forvar2113))) : $signed(reg2149));
                      reg2214 <= ($signed($signed((^~reg2194))) && (reg2067 ?
                          ((reg2053 || reg2102) << (forvar2184 || reg2091)) : (!(reg2069 ?
                              reg2141 : (8'hb5)))));
                      reg2215 <= reg2127;
                    end
                end
            end
          for (forvar2219 = (1'h0); (forvar2219 < (1'h0)); forvar2219 = (forvar2219 + (1'h1)))
            begin
              for (forvar2220 = (1'h0); (forvar2220 < (2'h3)); forvar2220 = (forvar2220 + (1'h1)))
                begin
                  for (forvar2221 = (1'h0); (forvar2221 < (1'h0)); forvar2221 = (forvar2221 + (1'h1)))
                    begin
                      reg2222 <= reg2079;
                      reg2223 <= $signed(($unsigned((|reg2151)) ?
                          reg2098[(2'h2):(1'h0)] : (reg2128 <= (forvar2046 ^~ forvar2210))));
                      reg2224 <= $signed($unsigned(($signed(reg2113) >> $signed(forvar2090))));
                    end
                end
              for (forvar2225 = (1'h0); (forvar2225 < (2'h3)); forvar2225 = (forvar2225 + (1'h1)))
                begin
                  if (($unsigned(((8'ha1) != {(8'ha8)})) ~^ reg2101))
                    begin
                      reg2226 <= (($signed((|forvar2151)) ?
                              $signed($signed(reg2083)) : {(^~reg2191)}) ?
                          reg2091 : {$signed((reg2125 ? (8'h9f) : reg2121))});
                    end
                  else
                    begin
                      reg2226 <= wire2042[(1'h0):(1'h0)];
                    end
                end
              if ((({forvar2192} <= $signed((reg2104 ? reg2123 : reg2141))) ?
                  ($signed(((8'h9e) != reg2060)) && (|(~&(8'hac)))) : (-forvar2115)))
                begin
                  if ((^forvar2147))
                    begin
                      reg2227 <= reg2154;
                      reg2228 <= (-(8'h9e));
                      reg2229 <= (+($unsigned((reg2118 ^ reg2130)) ?
                          $signed($signed(forvar2208)) : (forvar2138[(3'h4):(1'h1)] ?
                              reg2147 : (forvar2221 << (8'ha0)))));
                    end
                  else
                    begin
                      reg2227 <= reg2064;
                    end
                  if ($unsigned($unsigned({{reg2091}})))
                    begin
                      reg2230 <= $signed($unsigned(reg2193));
                    end
                  else
                    begin
                      reg2230 <= forvar2181;
                      reg2231 <= ($unsigned($unsigned({reg2110})) - $signed((~reg2229)));
                      reg2232 <= reg2120[(1'h0):(1'h0)];
                      reg2233 <= $unsigned(reg2074);
                    end
                end
              else
                begin
                  reg2227 <= ($unsigned((8'hba)) ^~ ($unsigned(reg2229) == {reg2185[(3'h5):(1'h1)]}));
                  for (forvar2228 = (1'h0); (forvar2228 < (2'h2)); forvar2228 = (forvar2228 + (1'h1)))
                    begin
                      reg2229 <= $signed(forvar2070);
                    end
                  if ($signed(($signed({reg2144}) ?
                      forvar2111[(1'h1):(1'h1)] : (forvar2049[(4'h8):(2'h2)] ?
                          $signed(reg2188) : (|reg2182)))))
                    begin
                      reg2230 <= reg2215[(4'ha):(4'ha)];
                      reg2231 <= ({{(^reg2214)}} >= ((forvar2075 ?
                          reg2233[(4'h9):(2'h3)] : (forvar2151 ?
                              reg2179 : reg2065)) * reg2188[(2'h2):(1'h1)]));
                      reg2232 <= $unsigned(((&reg2131) ?
                          reg2073[(3'h5):(2'h2)] : reg2115));
                      reg2233 <= forvar2058[(4'h9):(4'h9)];
                    end
                  else
                    begin
                      reg2230 <= ($unsigned((8'ha7)) == (&(&forvar2171[(4'ha):(2'h2)])));
                      reg2231 <= (reg2088[(3'h4):(1'h0)] ?
                          reg2160[(4'h8):(4'h8)] : (~&(reg2112 ?
                              (8'ha1) : forvar2096)));
                    end
                end
            end
        end
    end
  assign wire2234 = reg2140;
  assign wire2235 = $unsigned($signed(reg2127[(1'h1):(1'h1)]));
  always
    @(posedge clk) begin
      if ($signed($unsigned((!((8'hba) ? reg2096 : reg2078)))))
        begin
          for (forvar2236 = (1'h0); (forvar2236 < (1'h0)); forvar2236 = (forvar2236 + (1'h1)))
            begin
              if ({reg2197[(2'h2):(2'h2)]})
                begin
                  for (forvar2237 = (1'h0); (forvar2237 < (1'h1)); forvar2237 = (forvar2237 + (1'h1)))
                    begin
                      reg2238 <= $unsigned((reg2233[(4'ha):(3'h7)] >>> $unsigned((~reg2159))));
                      reg2239 <= {(reg2180[(1'h0):(1'h0)] ?
                              (~|(reg2102 <<< reg2211)) : $unsigned(reg2162))};
                      reg2240 <= ((^(8'ha4)) ?
                          (!$unsigned((reg2205 > reg2117))) : (|reg2054));
                    end
                  if ((^((&(&reg2142)) ~^ reg2060[(1'h1):(1'h1)])))
                    begin
                      reg2241 <= $signed((({wire2235} & reg2209) ?
                          reg2169 : (reg2211[(4'ha):(4'h8)] ?
                              (reg2186 ? reg2218 : reg2130) : (~reg2120))));
                    end
                  else
                    begin
                      reg2241 <= $signed(reg2175);
                      reg2242 <= (({(~^reg2211)} | {$signed(reg2054)}) ?
                          {reg2226} : reg2215[(2'h2):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar2237 = (1'h0); (forvar2237 < (1'h0)); forvar2237 = (forvar2237 + (1'h1)))
                    begin
                      reg2238 <= reg2115[(2'h3):(1'h1)];
                      reg2239 <= ($unsigned((~^(reg2050 ?
                          reg2186 : reg2222))) && reg2046);
                      reg2240 <= $unsigned($signed(reg2114));
                      reg2241 <= reg2156;
                    end
                  if ($unsigned(reg2173))
                    begin
                      reg2242 <= $unsigned((reg2178 ?
                          {$signed(reg2189)} : (~reg2129)));
                    end
                  else
                    begin
                      reg2242 <= (({(reg2230 * reg2239)} ?
                              (~&(reg2209 >= reg2129)) : reg2125) ?
                          $signed($unsigned((reg2142 + (8'hac)))) : (+$signed(reg2093[(4'hb):(3'h7)])));
                      reg2243 <= reg2048[(2'h2):(1'h0)];
                    end
                end
            end
          if (({((reg2124 ?
                  reg2210 : reg2097) * $signed(reg2084))} != $signed((|(reg2095 == reg2194)))))
            begin
              reg2244 <= $signed(reg2177);
              for (forvar2245 = (1'h0); (forvar2245 < (2'h3)); forvar2245 = (forvar2245 + (1'h1)))
                begin
                  reg2246 <= $unsigned(wire2042[(3'h4):(1'h0)]);
                  reg2247 <= $signed(($signed((reg2240 ?
                      reg2226 : reg2092)) ^~ ((&(8'hb5)) ?
                      reg2092[(1'h1):(1'h0)] : (reg2198 - reg2178))));
                  if (((($unsigned((8'haa)) ?
                      (reg2046 ? reg2121 : reg2133) : (reg2113 ?
                          reg2066 : reg2149)) >> (~|{(8'ha4)})) < $signed(reg2241)))
                    begin
                      reg2248 <= reg2201[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2248 <= $unsigned(reg2093[(4'hd):(3'h7)]);
                      reg2249 <= reg2170[(3'h6):(3'h4)];
                      reg2250 <= $unsigned($signed((&$signed(reg2206))));
                      reg2251 <= reg2118[(1'h0):(1'h0)];
                    end
                  for (forvar2252 = (1'h0); (forvar2252 < (2'h3)); forvar2252 = (forvar2252 + (1'h1)))
                    begin
                      reg2253 <= $unsigned(reg2082[(2'h3):(2'h3)]);
                    end
                end
            end
          else
            begin
              reg2244 <= ((~reg2082[(2'h2):(2'h2)]) || {$unsigned(reg2095[(1'h1):(1'h0)])});
              if (reg2153[(4'h8):(3'h7)])
                begin
                  for (forvar2245 = (1'h0); (forvar2245 < (1'h0)); forvar2245 = (forvar2245 + (1'h1)))
                    begin
                      reg2246 <= (8'hb9);
                      reg2247 <= (~((reg2148[(1'h0):(1'h0)] - {reg2215}) ?
                          (~&(reg2061 ?
                              reg2232 : reg2206)) : ({reg2150} & $signed(reg2131))));
                      reg2248 <= $unsigned($signed($unsigned(((8'haf) ?
                          reg2047 : reg2211))));
                    end
                  for (forvar2249 = (1'h0); (forvar2249 < (1'h1)); forvar2249 = (forvar2249 + (1'h1)))
                    begin
                      reg2250 <= reg2187[(4'h8):(1'h1)];
                      reg2251 <= $unsigned($signed($unsigned((~(8'hae)))));
                      reg2252 <= ((((~reg2108) != reg2238) << {$unsigned(wire2043)}) > reg2118);
                      reg2253 <= $unsigned((^~($unsigned(reg2194) ?
                          $unsigned(reg2098) : (^reg2191))));
                    end
                  for (forvar2254 = (1'h0); (forvar2254 < (2'h2)); forvar2254 = (forvar2254 + (1'h1)))
                    begin
                      reg2255 <= $signed($unsigned(reg2051[(1'h0):(1'h0)]));
                    end
                  for (forvar2256 = (1'h0); (forvar2256 < (2'h3)); forvar2256 = (forvar2256 + (1'h1)))
                    begin
                      reg2257 <= ($unsigned($signed($signed((8'hba)))) > ($signed((8'ha6)) ?
                          $unsigned((8'h9f)) : (reg2095 * (+reg2065))));
                      reg2258 <= reg2180;
                    end
                end
              else
                begin
                  for (forvar2245 = (1'h0); (forvar2245 < (2'h3)); forvar2245 = (forvar2245 + (1'h1)))
                    begin
                      reg2246 <= $signed($signed(reg2145));
                    end
                end
              if (reg2116[(2'h2):(1'h1)])
                begin
                  if ({(~reg2048)})
                    begin
                      reg2259 <= reg2204[(3'h6):(1'h0)];
                    end
                  else
                    begin
                      reg2259 <= wire2235;
                      reg2260 <= (reg2185 > reg2239);
                      reg2261 <= (((~&$unsigned(reg2201)) ^ ((reg2170 == reg2162) ?
                              $unsigned(reg2054) : (+reg2064))) ?
                          ({(reg2119 ?
                                  (8'hba) : reg2123)} << $unsigned($signed(reg2110))) : reg2074[(2'h2):(2'h2)]);
                    end
                  for (forvar2262 = (1'h0); (forvar2262 < (1'h1)); forvar2262 = (forvar2262 + (1'h1)))
                    begin
                      reg2263 <= (~^$signed((8'hac)));
                      reg2264 <= reg2222;
                    end
                  for (forvar2265 = (1'h0); (forvar2265 < (1'h1)); forvar2265 = (forvar2265 + (1'h1)))
                    begin
                      reg2266 <= $signed(($unsigned($signed((8'ha2))) && (wire2044 ?
                          (reg2162 ?
                              reg2217 : reg2226) : reg2241[(3'h4):(1'h1)])));
                      reg2267 <= (^~(((forvar2254 <<< reg2078) ?
                              (!forvar2265) : $signed(reg2227)) ?
                          reg2229[(2'h2):(2'h2)] : ((reg2227 ?
                              reg2076 : reg2218) * (reg2112 || reg2153))));
                    end
                end
              else
                begin
                  if ((^(~&forvar2245)))
                    begin
                      reg2259 <= $signed($signed($signed(reg2244)));
                    end
                  else
                    begin
                      reg2259 <= $unsigned($unsigned(reg2100[(4'hf):(4'hc)]));
                      reg2260 <= $signed(reg2244);
                      reg2261 <= ($unsigned(reg2126[(3'h4):(2'h3)]) > $signed(reg2127[(4'ha):(3'h5)]));
                      reg2262 <= $signed((($signed(reg2144) ?
                              reg2251 : $unsigned(reg2239)) ?
                          (reg2091 ?
                              reg2246[(3'h4):(2'h2)] : $unsigned(reg2098)) : ({forvar2252} < (^reg2067))));
                    end
                  reg2263 <= (reg2137 ?
                      reg2069 : ($unsigned({reg2054}) ^ reg2213));
                  for (forvar2264 = (1'h0); (forvar2264 < (1'h0)); forvar2264 = (forvar2264 + (1'h1)))
                    begin
                      reg2265 <= reg2057;
                      reg2266 <= (|$unsigned((8'hb1)));
                      reg2267 <= $unsigned($signed({$unsigned(reg2053)}));
                      reg2268 <= ($unsigned((~|(reg2223 ? (8'haf) : reg2100))) ?
                          $signed($unsigned((wire2040 | reg2150))) : ((!$signed(reg2206)) ^ (8'ha1)));
                    end
                  reg2269 <= (({(reg2243 ? reg2223 : reg2201)} ?
                          forvar2262[(1'h0):(1'h0)] : {$signed(reg2175)}) ?
                      $unsigned(((reg2052 ? reg2187 : (8'ha7)) ?
                          (~&reg2227) : $unsigned((8'hb6)))) : reg2178);
                end
              if ($unsigned($unsigned($signed($signed(reg2085)))))
                begin
                  for (forvar2270 = (1'h0); (forvar2270 < (2'h3)); forvar2270 = (forvar2270 + (1'h1)))
                    begin
                      reg2271 <= reg2046[(1'h0):(1'h0)];
                      reg2272 <= $unsigned($unsigned(((+(8'hb5)) << (reg2257 ?
                          reg2202 : reg2162))));
                      reg2273 <= $unsigned($signed(reg2091[(2'h2):(2'h2)]));
                    end
                  for (forvar2274 = (1'h0); (forvar2274 < (2'h3)); forvar2274 = (forvar2274 + (1'h1)))
                    begin
                      reg2275 <= reg2217[(1'h1):(1'h1)];
                      reg2276 <= $unsigned(reg2224[(3'h4):(1'h1)]);
                      reg2277 <= $unsigned((&reg2130[(3'h6):(2'h3)]));
                      reg2278 <= reg2112;
                    end
                  if ($signed({reg2114[(3'h6):(1'h0)]}))
                    begin
                      reg2279 <= $signed(($signed((reg2076 ~^ reg2094)) ?
                          $signed((reg2262 ~^ reg2187)) : reg2095));
                      reg2280 <= (((&$signed(reg2151)) ?
                              ($signed(reg2249) >= $unsigned((8'haf))) : reg2114[(3'h7):(3'h6)]) ?
                          $unsigned((~^reg2206)) : ($unsigned($unsigned(reg2119)) ?
                              (reg2085[(1'h0):(1'h0)] ?
                                  $signed(reg2050) : $signed(reg2078)) : ((~^reg2053) ?
                                  (reg2047 * reg2224) : reg2241)));
                    end
                  else
                    begin
                      reg2279 <= reg2097;
                      reg2280 <= ($unsigned(reg2054[(1'h1):(1'h1)]) ?
                          reg2148[(1'h0):(1'h0)] : ($unsigned(reg2276) ?
                              ($signed(reg2149) << $unsigned(reg2130)) : (((8'hb4) + reg2280) >> (reg2248 ?
                                  reg2230 : reg2132))));
                      reg2281 <= $signed(reg2124);
                      reg2282 <= (^~reg2215[(3'h6):(1'h0)]);
                    end
                end
              else
                begin
                  reg2270 <= {(~|$unsigned(reg2246))};
                  if ($signed($signed(reg2261[(1'h0):(1'h0)])))
                    begin
                      reg2271 <= (reg2134[(4'hc):(4'h8)] >>> (8'ha4));
                      reg2272 <= (!reg2229[(3'h4):(1'h0)]);
                      reg2273 <= reg2150;
                    end
                  else
                    begin
                      reg2271 <= {reg2079[(3'h5):(1'h1)]};
                    end
                  reg2274 <= reg2146;
                  if (reg2206[(2'h3):(2'h3)])
                    begin
                      reg2275 <= {reg2173[(1'h1):(1'h1)]};
                    end
                  else
                    begin
                      reg2275 <= reg2167[(4'ha):(3'h5)];
                      reg2276 <= reg2175[(4'ha):(4'h8)];
                      reg2277 <= (reg2178[(1'h1):(1'h0)] >>> $signed((~&reg2161)));
                      reg2278 <= ((&((reg2202 >> reg2186) ^ (reg2246 | reg2055))) << (~^reg2255[(2'h2):(2'h2)]));
                    end
                end
            end
          if (($signed((8'hb3)) ? reg2094 : ((~&reg2271) <<< reg2088)))
            begin
              for (forvar2283 = (1'h0); (forvar2283 < (1'h1)); forvar2283 = (forvar2283 + (1'h1)))
                begin
                  if ((~&reg2083))
                    begin
                      reg2284 <= (forvar2249[(1'h0):(1'h0)] && ($signed(((8'hae) ?
                          forvar2256 : reg2106)) << reg2274));
                      reg2285 <= {$unsigned($unsigned(reg2133))};
                    end
                  else
                    begin
                      reg2284 <= (($signed({(8'hba)}) <<< ($unsigned(reg2263) ?
                          (reg2274 ?
                              reg2226 : reg2104) : (8'ha0))) || $signed($unsigned((reg2211 ?
                          reg2148 : reg2246))));
                      reg2285 <= (&$signed(reg2141[(2'h2):(1'h0)]));
                      reg2286 <= $signed({{{reg2253}}});
                    end
                  reg2287 <= (reg2172[(1'h0):(1'h0)] + $signed((reg2209[(3'h7):(3'h6)] <<< $unsigned(reg2179))));
                  for (forvar2288 = (1'h0); (forvar2288 < (2'h3)); forvar2288 = (forvar2288 + (1'h1)))
                    begin
                      reg2289 <= (~&reg2183[(1'h1):(1'h1)]);
                    end
                  if (($signed($unsigned((reg2109 ?
                      (8'hb5) : reg2194))) >>> (^~$signed((reg2120 ?
                      reg2233 : reg2183)))))
                    begin
                      reg2290 <= $unsigned(reg2054[(3'h7):(1'h1)]);
                    end
                  else
                    begin
                      reg2290 <= $unsigned($unsigned(($signed((8'hb3)) ^~ (^~(8'ha8)))));
                    end
                end
              for (forvar2291 = (1'h0); (forvar2291 < (1'h0)); forvar2291 = (forvar2291 + (1'h1)))
                begin
                  for (forvar2292 = (1'h0); (forvar2292 < (1'h1)); forvar2292 = (forvar2292 + (1'h1)))
                    begin
                      reg2293 <= ((~^$unsigned(reg2203)) <= (8'ha8));
                      reg2294 <= $signed(($signed($signed(reg2050)) | ((reg2154 ~^ reg2161) ?
                          reg2065 : (forvar2264 ? forvar2274 : reg2285))));
                      reg2295 <= forvar2236;
                      reg2296 <= reg2106;
                    end
                end
              for (forvar2297 = (1'h0); (forvar2297 < (2'h2)); forvar2297 = (forvar2297 + (1'h1)))
                begin
                  for (forvar2298 = (1'h0); (forvar2298 < (1'h1)); forvar2298 = (forvar2298 + (1'h1)))
                    begin
                      reg2299 <= reg2188;
                      reg2300 <= ((|$signed({reg2116})) && $unsigned($signed(reg2251[(1'h0):(1'h0)])));
                      reg2301 <= {$signed(reg2167)};
                    end
                end
              if (reg2141[(3'h5):(1'h0)])
                begin
                  for (forvar2302 = (1'h0); (forvar2302 < (2'h3)); forvar2302 = (forvar2302 + (1'h1)))
                    begin
                      reg2303 <= (((+reg2094[(3'h4):(1'h0)]) ?
                          ((reg2127 ^ (8'ha9)) >>> reg2264) : ($signed((8'ha2)) >>> (forvar2256 << (8'ha5)))) & (8'hb2));
                    end
                  if ((^~{reg2078}))
                    begin
                      reg2304 <= {$signed(reg2115[(2'h3):(2'h2)])};
                    end
                  else
                    begin
                      reg2304 <= $signed((($unsigned(reg2239) >= $unsigned(reg2173)) > (~&reg2290[(3'h4):(2'h3)])));
                      reg2305 <= $signed(($unsigned({reg2232}) ?
                          $signed((reg2050 - reg2277)) : (reg2243[(1'h0):(1'h0)] ?
                              reg2238[(2'h2):(2'h2)] : $unsigned(reg2125))));
                      reg2306 <= ($unsigned(((~^reg2211) ?
                          $unsigned(reg2055) : (^~(8'ha7)))) >= $unsigned(reg2161));
                      reg2307 <= reg2306[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  reg2302 <= reg2250[(3'h7):(2'h3)];
                  for (forvar2303 = (1'h0); (forvar2303 < (2'h2)); forvar2303 = (forvar2303 + (1'h1)))
                    begin
                      reg2304 <= (~^(((reg2241 - reg2161) ?
                              {reg2098} : reg2140) ?
                          reg2212 : $unsigned((|reg2102))));
                    end
                  reg2305 <= $signed(reg2287);
                end
            end
          else
            begin
              for (forvar2283 = (1'h0); (forvar2283 < (2'h2)); forvar2283 = (forvar2283 + (1'h1)))
                begin
                  reg2284 <= $signed({(~(~reg2277))});
                end
              for (forvar2285 = (1'h0); (forvar2285 < (2'h3)); forvar2285 = (forvar2285 + (1'h1)))
                begin
                  if ((reg2187 >>> {$signed(reg2055)}))
                    begin
                      reg2286 <= $signed($unsigned($unsigned((reg2223 + reg2278))));
                    end
                  else
                    begin
                      reg2286 <= reg2120;
                      reg2287 <= (reg2250 ?
                          {(((8'h9e) ?
                                  (8'ha8) : reg2227) ^ (~&reg2173))} : $signed((8'hb1)));
                      reg2288 <= $unsigned((^(reg2214 - (reg2054 ?
                          reg2067 : reg2048))));
                      reg2289 <= $signed((~(|(reg2061 ? reg2186 : reg2275))));
                    end
                  for (forvar2290 = (1'h0); (forvar2290 < (2'h3)); forvar2290 = (forvar2290 + (1'h1)))
                    begin
                      reg2291 <= {$unsigned(((reg2259 ^~ reg2178) ?
                              reg2052 : reg2122))};
                    end
                  for (forvar2292 = (1'h0); (forvar2292 < (2'h3)); forvar2292 = (forvar2292 + (1'h1)))
                    begin
                      reg2293 <= reg2189[(3'h6):(1'h0)];
                      reg2294 <= (~$signed(reg2173));
                      reg2295 <= (reg2188 ?
                          $signed(reg2092) : {($signed(reg2084) <= {reg2294})});
                      reg2296 <= reg2253[(3'h7):(1'h1)];
                    end
                  if ($unsigned($unsigned((forvar2262[(2'h2):(1'h0)] + reg2177[(3'h4):(2'h2)]))))
                    begin
                      reg2297 <= $unsigned(reg2057);
                      reg2298 <= {$signed(reg2134)};
                      reg2299 <= $signed($signed(((&reg2066) ?
                          reg2046[(2'h2):(2'h2)] : (reg2250 ^ forvar2245))));
                    end
                  else
                    begin
                      reg2297 <= (-($signed(forvar2236) && $unsigned((reg2186 ?
                          reg2066 : reg2287))));
                      reg2298 <= reg2193;
                      reg2299 <= (|reg2275);
                      reg2300 <= (|reg2253);
                    end
                end
              for (forvar2301 = (1'h0); (forvar2301 < (2'h2)); forvar2301 = (forvar2301 + (1'h1)))
                begin
                  for (forvar2302 = (1'h0); (forvar2302 < (2'h3)); forvar2302 = (forvar2302 + (1'h1)))
                    begin
                      reg2303 <= $signed($unsigned(reg2051));
                    end
                end
              reg2304 <= (((reg2264 ? {(8'hba)} : $signed(reg2188)) ?
                  (~^{reg2305}) : reg2201) + reg2115);
            end
          for (forvar2308 = (1'h0); (forvar2308 < (1'h1)); forvar2308 = (forvar2308 + (1'h1)))
            begin
              if ($unsigned((-(reg2065[(3'h4):(1'h1)] & $unsigned((8'hb8))))))
                begin
                  if (reg2147)
                    begin
                      reg2309 <= reg2159[(4'ha):(3'h4)];
                      reg2310 <= reg2179[(3'h5):(1'h1)];
                      reg2311 <= $signed($signed(reg2210[(3'h7):(2'h3)]));
                    end
                  else
                    begin
                      reg2309 <= {$signed($signed((reg2300 || reg2053)))};
                    end
                  for (forvar2312 = (1'h0); (forvar2312 < (1'h0)); forvar2312 = (forvar2312 + (1'h1)))
                    begin
                      reg2313 <= reg2183;
                      reg2314 <= (($signed((reg2108 > (8'hb0))) ?
                              ((&reg2079) == reg2186[(1'h0):(1'h0)]) : (8'hb6)) ?
                          $signed(((reg2161 ? reg2116 : reg2242) ?
                              $unsigned((8'h9e)) : (reg2281 > reg2125))) : $unsigned((reg2116 ?
                              (reg2080 ? (8'ha0) : reg2097) : reg2259)));
                      reg2315 <= $unsigned($signed({$unsigned((8'ha0))}));
                      reg2316 <= reg2246[(4'h9):(3'h4)];
                    end
                end
              else
                begin
                  for (forvar2309 = (1'h0); (forvar2309 < (2'h2)); forvar2309 = (forvar2309 + (1'h1)))
                    begin
                      reg2310 <= ($signed((!forvar2252)) * ({(reg2115 ?
                                  (8'hba) : (8'hb9))} ?
                          ((reg2060 + reg2241) ?
                              reg2231[(3'h5):(3'h5)] : reg2162[(3'h5):(1'h1)]) : reg2304[(2'h2):(1'h1)]));
                    end
                  reg2311 <= $signed((-(~|reg2301[(3'h4):(2'h3)])));
                  for (forvar2312 = (1'h0); (forvar2312 < (1'h0)); forvar2312 = (forvar2312 + (1'h1)))
                    begin
                      reg2313 <= {$unsigned($signed((reg2107 <<< reg2222)))};
                    end
                end
            end
        end
      else
        begin
          if ((~&reg2284))
            begin
              for (forvar2236 = (1'h0); (forvar2236 < (2'h3)); forvar2236 = (forvar2236 + (1'h1)))
                begin
                  for (forvar2237 = (1'h0); (forvar2237 < (2'h2)); forvar2237 = (forvar2237 + (1'h1)))
                    begin
                      reg2238 <= reg2271;
                      reg2239 <= reg2284;
                      reg2240 <= $signed(reg2281);
                      reg2241 <= reg2195;
                    end
                  for (forvar2242 = (1'h0); (forvar2242 < (1'h1)); forvar2242 = (forvar2242 + (1'h1)))
                    begin
                      reg2243 <= {(forvar2308[(2'h2):(1'h1)] ?
                              reg2056 : $signed(((8'hae) ?
                                  reg2279 : reg2264)))};
                      reg2244 <= ((~&{reg2239}) ?
                          reg2175 : $unsigned((~(reg2144 ?
                              (8'hb2) : reg2162))));
                      reg2245 <= $signed({$signed($unsigned(reg2098))});
                    end
                  reg2246 <= (reg2084 >> reg2281[(1'h0):(1'h0)]);
                  reg2247 <= $unsigned(reg2224[(3'h7):(3'h6)]);
                end
              for (forvar2248 = (1'h0); (forvar2248 < (1'h0)); forvar2248 = (forvar2248 + (1'h1)))
                begin
                  if (reg2130[(2'h3):(2'h3)])
                    begin
                      reg2249 <= $signed($unsigned($unsigned((reg2173 ?
                          reg2279 : reg2223))));
                      reg2250 <= (~&$signed(reg2175[(4'he):(4'h8)]));
                      reg2251 <= $unsigned((({(8'ha3)} ?
                          reg2149[(2'h2):(1'h1)] : $unsigned(reg2110)) >> (~|(reg2169 ?
                          reg2241 : reg2209))));
                      reg2252 <= (8'ha2);
                    end
                  else
                    begin
                      reg2249 <= $unsigned((reg2274[(2'h3):(1'h0)] != $unsigned((reg2095 ?
                          reg2215 : reg2091))));
                      reg2250 <= (reg2153 ?
                          reg2189[(3'h6):(3'h6)] : $unsigned(reg2084[(3'h5):(2'h2)]));
                    end
                  if ($signed(((|$signed(reg2275)) ?
                      (8'ha3) : reg2262[(1'h1):(1'h1)])))
                    begin
                      reg2253 <= $signed((~(reg2270[(2'h3):(1'h1)] > (reg2266 ?
                          reg2276 : reg2271))));
                      reg2254 <= ($signed($signed((^~forvar2312))) ?
                          (&(~reg2296)) : (~^$signed((reg2204 ?
                              forvar2301 : reg2170))));
                    end
                  else
                    begin
                      reg2253 <= $signed((reg2085 ?
                          $unsigned($unsigned(reg2261)) : forvar2254[(3'h7):(3'h7)]));
                      reg2254 <= (reg2218[(2'h2):(2'h2)] ?
                          $signed((reg2264 & (reg2154 ?
                              (8'hb8) : reg2080))) : (reg2107[(1'h1):(1'h1)] >> (reg2250[(3'h4):(1'h0)] ?
                              ((8'haa) ? forvar2301 : reg2107) : reg2048)));
                    end
                  for (forvar2255 = (1'h0); (forvar2255 < (2'h2)); forvar2255 = (forvar2255 + (1'h1)))
                    begin
                      reg2256 <= $unsigned(reg2078[(4'ha):(1'h1)]);
                      reg2257 <= ($unsigned($signed($signed(reg2084))) ?
                          reg2272 : ($unsigned($unsigned(reg2303)) ?
                              $unsigned($signed(reg2251)) : $unsigned((8'haf))));
                    end
                  if (reg2253[(1'h1):(1'h0)])
                    begin
                      reg2258 <= reg2084[(4'ha):(4'h9)];
                      reg2259 <= forvar2265;
                    end
                  else
                    begin
                      reg2258 <= reg2282;
                    end
                end
              if ((^{reg2084}))
                begin
                  for (forvar2260 = (1'h0); (forvar2260 < (1'h1)); forvar2260 = (forvar2260 + (1'h1)))
                    begin
                      reg2261 <= {reg2255[(4'h9):(1'h0)]};
                    end
                  for (forvar2262 = (1'h0); (forvar2262 < (1'h1)); forvar2262 = (forvar2262 + (1'h1)))
                    begin
                      reg2263 <= (reg2116 != ((^~(reg2103 ?
                          forvar2308 : reg2108)) || (^~forvar2262)));
                      reg2264 <= $unsigned(({(~&reg2109)} ?
                          (-reg2082) : reg2302[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  if ((reg2300[(3'h4):(1'h1)] ?
                      ($signed((-(8'hae))) ^ (forvar2245[(1'h0):(1'h0)] ^ $signed(forvar2308))) : ({reg2223} ?
                          reg2169 : (~(reg2215 ? forvar2308 : reg2048)))))
                    begin
                      reg2260 <= reg2278;
                    end
                  else
                    begin
                      reg2260 <= $unsigned(forvar2312);
                    end
                  if (reg2197)
                    begin
                      reg2261 <= ({((reg2095 - (8'hb5)) * ((8'ha8) ?
                                  reg2137 : wire2041))} ?
                          ($unsigned((+reg2175)) ?
                              (^(&reg2049)) : reg2159[(3'h5):(1'h1)]) : ($unsigned($unsigned(forvar2274)) & ((reg2210 <<< reg2303) || reg2119)));
                      reg2262 <= reg2099;
                      reg2263 <= $signed(forvar2274);
                      reg2264 <= wire2235[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2261 <= $signed(reg2215[(3'h4):(2'h2)]);
                      reg2262 <= $signed((8'ha3));
                      reg2263 <= reg2189;
                    end
                end
            end
          else
            begin
              if (reg2282)
                begin
                  for (forvar2236 = (1'h0); (forvar2236 < (2'h2)); forvar2236 = (forvar2236 + (1'h1)))
                    begin
                      reg2237 <= forvar2288;
                      reg2238 <= (($signed($signed(reg2153)) < $unsigned($signed(reg2153))) ?
                          ((8'hb6) ^ $signed(reg2112)) : reg2142[(3'h7):(3'h5)]);
                      reg2239 <= ($signed(reg2053[(1'h0):(1'h0)]) ~^ $unsigned($signed((+forvar2302))));
                      reg2240 <= ({$signed((reg2187 ? reg2106 : reg2091))} ?
                          $unsigned($unsigned((reg2262 ?
                              forvar2237 : reg2167))) : (!(|$unsigned(reg2202))));
                    end
                  for (forvar2241 = (1'h0); (forvar2241 < (1'h0)); forvar2241 = (forvar2241 + (1'h1)))
                    begin
                      reg2242 <= $unsigned($unsigned(forvar2274[(3'h7):(3'h4)]));
                      reg2243 <= {{($unsigned(reg2189) || (8'hb7))}};
                    end
                  reg2244 <= (8'hb9);
                end
              else
                begin
                  for (forvar2236 = (1'h0); (forvar2236 < (2'h2)); forvar2236 = (forvar2236 + (1'h1)))
                    begin
                      reg2237 <= (forvar2264 == (($unsigned(reg2243) ?
                          reg2264 : reg2205) >> $unsigned((^reg2098))));
                      reg2238 <= $signed({$unsigned($unsigned(forvar2260))});
                      reg2239 <= ({$signed((reg2267 + wire2041))} >>> (^(~reg2301)));
                      reg2240 <= wire2041;
                    end
                  reg2241 <= reg2110;
                  if (($signed(((~|reg2074) ?
                      reg2249[(3'h5):(1'h0)] : reg2132[(4'h8):(2'h3)])) < ((((8'h9f) ?
                      reg2123 : reg2266) >= (~reg2313)) - $signed($signed((8'ha2))))))
                    begin
                      reg2242 <= ($unsigned($signed((~&reg2115))) ?
                          reg2316[(2'h2):(1'h0)] : reg2114[(4'h9):(4'h9)]);
                    end
                  else
                    begin
                      reg2242 <= {reg2217[(3'h5):(2'h2)]};
                      reg2243 <= $unsigned(((reg2179[(1'h1):(1'h0)] ?
                              reg2300 : $signed(reg2185)) ?
                          (-(reg2310 ?
                              reg2260 : reg2242)) : $unsigned({(8'haf)})));
                      reg2244 <= ($signed((reg2191 ?
                              reg2223[(1'h1):(1'h0)] : (reg2134 + reg2270))) ?
                          (~|(~&reg2095)) : $unsigned(reg2307));
                    end
                  if (($signed($signed(reg2175)) || $signed($signed(reg2137))))
                    begin
                      reg2245 <= $signed((8'hb2));
                    end
                  else
                    begin
                      reg2245 <= $signed($signed(reg2115));
                      reg2246 <= reg2137;
                      reg2247 <= (reg2277 && (8'h9c));
                    end
                end
            end
          for (forvar2265 = (1'h0); (forvar2265 < (2'h3)); forvar2265 = (forvar2265 + (1'h1)))
            begin
              if ($signed({$unsigned($signed(reg2066))}))
                begin
                  for (forvar2266 = (1'h0); (forvar2266 < (2'h2)); forvar2266 = (forvar2266 + (1'h1)))
                    begin
                      reg2267 <= reg2098;
                      reg2268 <= (~&((reg2240[(2'h3):(1'h0)] ?
                              reg2188 : $unsigned(reg2080)) ?
                          (&reg2146[(4'hb):(1'h1)]) : (reg2194[(1'h0):(1'h0)] ?
                              reg2309 : (reg2293 ^~ reg2118))));
                    end
                  reg2269 <= ($signed((!(~reg2097))) == (~reg2060));
                  for (forvar2270 = (1'h0); (forvar2270 < (2'h2)); forvar2270 = (forvar2270 + (1'h1)))
                    begin
                      reg2271 <= $signed(reg2188);
                    end
                  if ({{reg2294}})
                    begin
                      reg2272 <= (($signed(reg2110) ?
                              (^(reg2140 || reg2256)) : $signed($signed(reg2107))) ?
                          (~(~&reg2140[(1'h1):(1'h1)])) : reg2109[(1'h1):(1'h1)]);
                      reg2273 <= (((reg2046[(2'h2):(1'h0)] > $signed((8'hb0))) ?
                              ($signed(forvar2252) ?
                                  {reg2233} : $unsigned(reg2166)) : ($unsigned(reg2291) ?
                                  {(8'ha6)} : $unsigned(reg2273))) ?
                          (~&($unsigned((8'hb6)) >>> $signed(reg2205))) : $unsigned(reg2237[(2'h3):(1'h0)]));
                      reg2274 <= reg2307;
                    end
                  else
                    begin
                      reg2272 <= reg2187[(1'h1):(1'h0)];
                      reg2273 <= (!reg2172);
                      reg2274 <= reg2239[(2'h2):(1'h1)];
                    end
                end
              else
                begin
                  if ((|(reg2122[(1'h1):(1'h1)] ^~ {(^~reg2216)})))
                    begin
                      reg2266 <= ({(reg2257 ? $signed((8'hb3)) : (~|reg2223))} ?
                          (({reg2223} && (reg2130 >= reg2131)) == (+(&reg2113))) : reg2161[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg2266 <= forvar2248[(2'h2):(2'h2)];
                      reg2267 <= $signed(reg2288);
                      reg2268 <= (reg2285[(1'h0):(1'h0)] & $unsigned((reg2137 ?
                          $unsigned(reg2122) : $unsigned(reg2228))));
                    end
                  for (forvar2269 = (1'h0); (forvar2269 < (2'h3)); forvar2269 = (forvar2269 + (1'h1)))
                    begin
                      reg2270 <= $unsigned($signed((+(~|(8'hb7)))));
                      reg2271 <= {reg2084};
                      reg2272 <= (~($unsigned({(8'ha5)}) >> ($signed((8'ha6)) ?
                          (+(8'hb3)) : reg2202)));
                    end
                  for (forvar2273 = (1'h0); (forvar2273 < (2'h2)); forvar2273 = (forvar2273 + (1'h1)))
                    begin
                      reg2274 <= reg2271;
                      reg2275 <= $unsigned($signed({(reg2080 <<< (8'hb1))}));
                      reg2276 <= reg2228;
                    end
                  if (reg2255[(3'h7):(3'h6)])
                    begin
                      reg2277 <= {$unsigned($unsigned(((8'hb6) + reg2166)))};
                      reg2278 <= (^$unsigned((reg2263 ?
                          $unsigned(forvar2241) : (reg2129 >>> wire2234))));
                      reg2279 <= reg2309;
                    end
                  else
                    begin
                      reg2277 <= reg2119;
                      reg2278 <= (reg2297[(3'h5):(2'h2)] & (~&reg2093));
                    end
                end
              for (forvar2280 = (1'h0); (forvar2280 < (2'h2)); forvar2280 = (forvar2280 + (1'h1)))
                begin
                  for (forvar2281 = (1'h0); (forvar2281 < (1'h0)); forvar2281 = (forvar2281 + (1'h1)))
                    begin
                      reg2282 <= $signed((({reg2286} > $unsigned(reg2160)) >>> reg2174[(4'hd):(3'h4)]));
                      reg2283 <= reg2182;
                      reg2284 <= reg2069;
                    end
                  for (forvar2285 = (1'h0); (forvar2285 < (1'h0)); forvar2285 = (forvar2285 + (1'h1)))
                    begin
                      reg2286 <= $signed({(-reg2079)});
                      reg2287 <= $unsigned($signed({reg2272}));
                      reg2288 <= $signed(reg2248);
                      reg2289 <= ((8'hae) ? reg2272 : reg2305[(1'h1):(1'h0)]);
                    end
                  if ($unsigned($unsigned($unsigned((forvar2303 - reg2267)))))
                    begin
                      reg2290 <= (((~^(~^reg2047)) ?
                          ({reg2160} ?
                              (reg2202 >> reg2161) : reg2250) : reg2222) - ($unsigned($unsigned(reg2306)) ?
                          reg2095[(2'h2):(1'h0)] : ((reg2161 ?
                                  forvar2309 : reg2101) ?
                              $signed(reg2263) : $signed(reg2050))));
                    end
                  else
                    begin
                      reg2290 <= (reg2194 ?
                          ({(reg2210 ? reg2213 : reg2283)} ?
                              $signed(reg2052) : ($unsigned(reg2173) ~^ reg2102[(1'h0):(1'h0)])) : ((((8'ha5) ?
                                      reg2210 : reg2072) ?
                                  $unsigned((8'hb4)) : (reg2260 <<< reg2082)) ?
                              ($signed(reg2148) ?
                                  (~|reg2104) : (reg2109 ?
                                      forvar2237 : (8'hba))) : reg2303));
                      reg2291 <= reg2178[(1'h0):(1'h0)];
                      reg2292 <= $signed((^$unsigned((reg2301 != (8'ha3)))));
                    end
                end
              if ((~(reg2095[(3'h4):(1'h1)] < reg2182)))
                begin
                  if ((^(~|$unsigned($unsigned(reg2304)))))
                    begin
                      reg2293 <= (|reg2057);
                    end
                  else
                    begin
                      reg2293 <= $signed($unsigned({(reg2073 & reg2116)}));
                      reg2294 <= (8'haf);
                    end
                  for (forvar2295 = (1'h0); (forvar2295 < (2'h3)); forvar2295 = (forvar2295 + (1'h1)))
                    begin
                      reg2296 <= (~^(((reg2082 ?
                              reg2122 : reg2266) | (~|reg2134)) ?
                          (reg2272[(3'h5):(2'h2)] + (reg2188 << reg2081)) : (8'ha2)));
                      reg2297 <= reg2282;
                      reg2298 <= $unsigned((reg2123[(2'h3):(1'h1)] != $unsigned({forvar2249})));
                      reg2299 <= ((((reg2293 ? reg2249 : reg2284) ?
                              reg2077 : reg2067) << (forvar2273[(4'h9):(3'h7)] >>> ((8'ha9) + reg2177))) ?
                          (~|{(reg2074 ?
                                  reg2245 : reg2121)}) : (reg2133[(4'hd):(3'h6)] >> {reg2293}));
                    end
                end
              else
                begin
                  reg2293 <= reg2079;
                  reg2294 <= $unsigned({$signed($signed(reg2254))});
                  for (forvar2295 = (1'h0); (forvar2295 < (2'h2)); forvar2295 = (forvar2295 + (1'h1)))
                    begin
                      reg2296 <= reg2298[(1'h0):(1'h0)];
                      reg2297 <= $signed($signed($signed($signed((8'hb1)))));
                      reg2298 <= ({$unsigned((-reg2179))} ~^ (8'hb0));
                      reg2299 <= reg2098[(3'h4):(2'h3)];
                    end
                  if ((reg2103 ? reg2202 : $signed(reg2132)))
                    begin
                      reg2300 <= (~&$signed(forvar2242));
                      reg2301 <= $signed((~(8'hac)));
                    end
                  else
                    begin
                      reg2300 <= reg2132[(3'h5):(3'h5)];
                    end
                end
            end
          reg2302 <= (^$signed((^~$unsigned(reg2276))));
          for (forvar2303 = (1'h0); (forvar2303 < (2'h3)); forvar2303 = (forvar2303 + (1'h1)))
            begin
              if (($unsigned((8'ha5)) && (-$unsigned($unsigned(reg2239)))))
                begin
                  for (forvar2304 = (1'h0); (forvar2304 < (2'h3)); forvar2304 = (forvar2304 + (1'h1)))
                    begin
                      reg2305 <= reg2232;
                      reg2306 <= ($signed(($unsigned(reg2050) ?
                              (wire2043 ?
                                  reg2215 : reg2128) : reg2178[(2'h2):(2'h2)])) ?
                          reg2238[(1'h0):(1'h0)] : $unsigned(reg2288));
                      reg2307 <= {reg2231[(3'h5):(2'h3)]};
                    end
                  for (forvar2308 = (1'h0); (forvar2308 < (1'h0)); forvar2308 = (forvar2308 + (1'h1)))
                    begin
                      reg2309 <= reg2053[(1'h0):(1'h0)];
                      reg2310 <= (-($unsigned($signed((8'haa))) ?
                          reg2288 : $signed(reg2257)));
                      reg2311 <= reg2100[(1'h1):(1'h1)];
                      reg2312 <= {$signed($unsigned($signed(reg2277)))};
                    end
                end
              else
                begin
                  if ((8'ha2))
                    begin
                      reg2304 <= (~&(reg2302 && {(reg2175 ?
                              forvar2264 : reg2197)}));
                      reg2305 <= (($unsigned(((8'hae) ? (8'hb6) : (8'haa))) ?
                          (reg2167[(2'h2):(1'h0)] << (reg2278 ?
                              forvar2254 : reg2054)) : (reg2293 ?
                              $signed(reg2270) : {reg2212})) ^~ reg2067[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg2304 <= {$signed({reg2247[(1'h1):(1'h1)]})};
                    end
                  for (forvar2306 = (1'h0); (forvar2306 < (1'h1)); forvar2306 = (forvar2306 + (1'h1)))
                    begin
                      reg2307 <= reg2215[(3'h7):(2'h2)];
                    end
                  if (reg2185)
                    begin
                      reg2308 <= (reg2287 ?
                          $unsigned((forvar2297 <= (^~reg2212))) : reg2097[(2'h3):(1'h1)]);
                      reg2309 <= ($signed(reg2213) - ($signed((reg2123 ?
                              reg2201 : (8'hac))) ?
                          $signed((reg2205 ?
                              reg2299 : forvar2297)) : $unsigned($signed(reg2100))));
                      reg2310 <= {(|$signed((~|forvar2285)))};
                      reg2311 <= ((((reg2204 || reg2228) >> $signed(reg2190)) << forvar2262) ?
                          reg2307[(2'h3):(1'h0)] : ($signed($signed(reg2211)) ?
                              ($signed((8'ha4)) <<< ((8'ha5) ?
                                  reg2148 : (8'hb3))) : {(reg2186 ?
                                      reg2290 : reg2193)}));
                    end
                  else
                    begin
                      reg2308 <= reg2172[(1'h1):(1'h1)];
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2317 = (1'h0); (forvar2317 < (2'h2)); forvar2317 = (forvar2317 + (1'h1)))
        begin
          for (forvar2318 = (1'h0); (forvar2318 < (2'h2)); forvar2318 = (forvar2318 + (1'h1)))
            begin
              if (reg2305[(2'h2):(2'h2)])
                begin
                  if (reg2093[(3'h4):(1'h1)])
                    begin
                      reg2319 <= ($signed($unsigned(reg2304[(3'h4):(1'h0)])) >= ((8'haa) + reg2307[(3'h5):(3'h5)]));
                    end
                  else
                    begin
                      reg2319 <= $unsigned(reg2187[(4'hb):(2'h2)]);
                    end
                  reg2320 <= reg2056[(4'h8):(3'h5)];
                  for (forvar2321 = (1'h0); (forvar2321 < (1'h1)); forvar2321 = (forvar2321 + (1'h1)))
                    begin
                      reg2322 <= $unsigned($unsigned({reg2113}));
                      reg2323 <= $unsigned((&({(8'ha6)} ^~ (|reg2092))));
                    end
                  reg2324 <= (($unsigned($unsigned(reg2119)) ~^ reg2067[(2'h3):(2'h3)]) ?
                      (reg2144[(3'h4):(2'h2)] ?
                          $unsigned(reg2238[(2'h2):(2'h2)]) : reg2320) : (reg2202 ?
                          reg2094[(4'hb):(1'h1)] : (^~((8'hb8) ?
                              reg2050 : (8'haf)))));
                end
              else
                begin
                  for (forvar2319 = (1'h0); (forvar2319 < (1'h1)); forvar2319 = (forvar2319 + (1'h1)))
                    begin
                      reg2320 <= $signed($unsigned($signed((!reg2217))));
                    end
                end
              for (forvar2325 = (1'h0); (forvar2325 < (1'h0)); forvar2325 = (forvar2325 + (1'h1)))
                begin
                  for (forvar2326 = (1'h0); (forvar2326 < (2'h2)); forvar2326 = (forvar2326 + (1'h1)))
                    begin
                      reg2327 <= (($unsigned(reg2315) ?
                              $unsigned(reg2067) : {$unsigned(reg2263)}) ?
                          (+($signed((8'h9d)) - (8'ha1))) : (8'hb9));
                      reg2328 <= ($unsigned(((|reg2156) & (reg2116 ?
                              (8'hb9) : (8'ha8)))) ?
                          (($unsigned(reg2131) ?
                                  $signed(reg2281) : (reg2245 >= reg2066)) ?
                              (8'ha2) : wire2234[(3'h7):(2'h2)]) : ((~&(reg2049 - reg2194)) ?
                              $unsigned($unsigned(reg2162)) : reg2314[(3'h7):(3'h6)]));
                      reg2329 <= ($signed(reg2169[(2'h3):(1'h1)]) >> reg2214);
                    end
                  for (forvar2330 = (1'h0); (forvar2330 < (1'h0)); forvar2330 = (forvar2330 + (1'h1)))
                    begin
                      reg2331 <= (^(reg2049 ?
                          ({reg2091} ?
                              $unsigned(reg2194) : reg2217) : (~^reg2191)));
                    end
                  for (forvar2332 = (1'h0); (forvar2332 < (1'h0)); forvar2332 = (forvar2332 + (1'h1)))
                    begin
                      reg2333 <= reg2096[(1'h0):(1'h0)];
                      reg2334 <= ((8'haf) | ((~|$signed(reg2069)) ?
                          forvar2319[(2'h2):(2'h2)] : {(!reg2155)}));
                    end
                  if ((reg2323 * reg2256))
                    begin
                      reg2335 <= (reg2193 ?
                          $unsigned({reg2324}) : ($signed($signed(reg2224)) ~^ {(8'hae)}));
                      reg2336 <= $signed($unsigned($unsigned(reg2323)));
                      reg2337 <= (&(&$unsigned((reg2237 <<< wire2040))));
                    end
                  else
                    begin
                      reg2335 <= reg2173[(4'h9):(3'h7)];
                      reg2336 <= $unsigned($signed(wire2235[(2'h2):(1'h0)]));
                    end
                end
              for (forvar2338 = (1'h0); (forvar2338 < (2'h2)); forvar2338 = (forvar2338 + (1'h1)))
                begin
                  reg2339 <= ($signed($signed({reg2198})) != $unsigned(reg2294[(4'h9):(1'h0)]));
                end
            end
          reg2340 <= $signed(reg2294);
          for (forvar2341 = (1'h0); (forvar2341 < (1'h1)); forvar2341 = (forvar2341 + (1'h1)))
            begin
              for (forvar2342 = (1'h0); (forvar2342 < (2'h3)); forvar2342 = (forvar2342 + (1'h1)))
                begin
                  reg2343 <= (reg2302[(2'h2):(1'h0)] ^ {$unsigned((~^reg2108))});
                end
              for (forvar2344 = (1'h0); (forvar2344 < (1'h1)); forvar2344 = (forvar2344 + (1'h1)))
                begin
                  if ((~^{wire2042}))
                    begin
                      reg2345 <= ($unsigned(reg2257[(2'h3):(2'h3)]) <= reg2343);
                      reg2346 <= reg2117;
                    end
                  else
                    begin
                      reg2345 <= reg2191;
                      reg2346 <= $unsigned($unsigned($signed(reg2106[(4'hb):(3'h7)])));
                    end
                  if ((8'ha0))
                    begin
                      reg2347 <= (8'h9c);
                    end
                  else
                    begin
                      reg2347 <= $unsigned(reg2059);
                      reg2348 <= reg2316[(2'h3):(1'h1)];
                    end
                  if (reg2276)
                    begin
                      reg2349 <= $signed((|reg2286));
                    end
                  else
                    begin
                      reg2349 <= ($unsigned(reg2115) ?
                          $signed((~&reg2113[(3'h7):(3'h5)])) : ($unsigned(reg2114) ?
                              reg2057[(3'h7):(3'h5)] : reg2194));
                      reg2350 <= reg2099;
                      reg2351 <= $unsigned(($unsigned($unsigned((8'ha5))) ?
                          ((reg2261 ? reg2335 : (8'hb0)) ?
                              (^(8'ha5)) : reg2265[(1'h0):(1'h0)]) : ((reg2301 ?
                              reg2179 : reg2278) ~^ (reg2267 ?
                              reg2126 : reg2061))));
                      reg2352 <= ($signed((~((8'ha7) << (8'ha9)))) ?
                          reg2237[(2'h3):(2'h3)] : reg2349[(4'h9):(3'h5)]);
                    end
                end
              for (forvar2353 = (1'h0); (forvar2353 < (1'h0)); forvar2353 = (forvar2353 + (1'h1)))
                begin
                  if ((((reg2098[(2'h2):(2'h2)] <<< {forvar2338}) ?
                      reg2261[(3'h4):(2'h3)] : reg2080[(3'h6):(3'h5)]) < (^~(reg2098 + (8'hb9)))))
                    begin
                      reg2354 <= $unsigned(reg2333);
                      reg2355 <= reg2250;
                      reg2356 <= $signed(reg2206);
                      reg2357 <= (reg2124[(1'h0):(1'h0)] >>> (({reg2121} || $unsigned((8'ha1))) | (((8'h9e) ?
                          reg2149 : (8'hb4)) >= $unsigned(reg2303))));
                    end
                  else
                    begin
                      reg2354 <= $signed($signed($signed($signed((8'had)))));
                      reg2355 <= (~^(^reg2287[(2'h3):(2'h3)]));
                      reg2356 <= ((&$unsigned((forvar2326 ?
                          reg2094 : reg2232))) || {((-reg2313) ^~ reg2302)});
                    end
                  if (reg2268[(3'h5):(3'h4)])
                    begin
                      reg2358 <= (~|{reg2301[(3'h5):(3'h4)]});
                    end
                  else
                    begin
                      reg2358 <= $unsigned((8'hba));
                    end
                  if (reg2088[(3'h5):(1'h0)])
                    begin
                      reg2359 <= ($unsigned(reg2356[(2'h2):(1'h1)]) || $signed(reg2155));
                      reg2360 <= reg2244[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2359 <= reg2190[(3'h4):(1'h1)];
                      reg2360 <= $signed($unsigned(((~|reg2275) ?
                          {reg2183} : reg2324)));
                      reg2361 <= reg2274[(2'h3):(2'h3)];
                      reg2362 <= {reg2328};
                    end
                end
              for (forvar2363 = (1'h0); (forvar2363 < (2'h3)); forvar2363 = (forvar2363 + (1'h1)))
                begin
                  for (forvar2364 = (1'h0); (forvar2364 < (2'h3)); forvar2364 = (forvar2364 + (1'h1)))
                    begin
                      reg2365 <= (reg2269[(3'h6):(2'h3)] ?
                          {(-{reg2263})} : reg2337[(3'h4):(1'h0)]);
                    end
                  for (forvar2366 = (1'h0); (forvar2366 < (1'h1)); forvar2366 = (forvar2366 + (1'h1)))
                    begin
                      reg2367 <= $signed($unsigned({(forvar2341 ?
                              reg2300 : reg2188)}));
                      reg2368 <= $signed({(~^reg2313)});
                      reg2369 <= reg2148;
                      reg2370 <= (wire2044 ?
                          (!(!$unsigned((8'hb2)))) : reg2175);
                    end
                  for (forvar2371 = (1'h0); (forvar2371 < (2'h2)); forvar2371 = (forvar2371 + (1'h1)))
                    begin
                      reg2372 <= (~|$signed(((reg2108 ? reg2046 : reg2183) ?
                          (~reg2137) : (~reg2098))));
                      reg2373 <= (!reg2076);
                      reg2374 <= {(&$signed({(8'ha6)}))};
                      reg2375 <= reg2193;
                    end
                  if (reg2095)
                    begin
                      reg2376 <= reg2103;
                      reg2377 <= (8'hb5);
                      reg2378 <= {$signed(((^reg2242) ?
                              ((8'hb8) ^ (8'h9c)) : $signed((8'hb9))))};
                      reg2379 <= (reg2156 ?
                          ($unsigned($signed(reg2173)) ?
                              (-reg2154) : ($unsigned(reg2150) ?
                                  $signed(reg2336) : (reg2064 || reg2285))) : (8'haf));
                    end
                  else
                    begin
                      reg2376 <= reg2222;
                    end
                end
            end
          if ({reg2253})
            begin
              for (forvar2380 = (1'h0); (forvar2380 < (1'h1)); forvar2380 = (forvar2380 + (1'h1)))
                begin
                  if ((^~reg2148))
                    begin
                      reg2381 <= reg2085;
                      reg2382 <= reg2177[(2'h2):(2'h2)];
                      reg2383 <= (^({$unsigned(reg2072)} ?
                          $unsigned($signed(reg2218)) : ($unsigned(reg2280) >= $unsigned(reg2177))));
                    end
                  else
                    begin
                      reg2381 <= (reg2215 ?
                          $unsigned(reg2151[(1'h0):(1'h0)]) : {$signed($unsigned(reg2072))});
                    end
                end
            end
          else
            begin
              for (forvar2380 = (1'h0); (forvar2380 < (1'h1)); forvar2380 = (forvar2380 + (1'h1)))
                begin
                  for (forvar2381 = (1'h0); (forvar2381 < (2'h2)); forvar2381 = (forvar2381 + (1'h1)))
                    begin
                      reg2382 <= (~|reg2383[(1'h1):(1'h1)]);
                      reg2383 <= ((&(reg2144[(4'hc):(3'h5)] ?
                          (^~reg2097) : (reg2273 ?
                              reg2372 : reg2316))) & reg2071[(4'hd):(4'hc)]);
                      reg2384 <= reg2152;
                    end
                  if ($signed($unsigned((+(reg2296 << reg2096)))))
                    begin
                      reg2385 <= (^reg2286);
                      reg2386 <= $signed(reg2242);
                      reg2387 <= ($signed(({reg2300} ?
                              reg2279 : $unsigned(reg2375))) ?
                          $unsigned(wire2234) : reg2348);
                      reg2388 <= $signed({reg2077[(4'ha):(1'h1)]});
                    end
                  else
                    begin
                      reg2385 <= {$unsigned((~|$unsigned((8'had))))};
                      reg2386 <= ($unsigned(reg2311[(4'h9):(2'h3)]) >= $unsigned(($unsigned(reg2146) ?
                          $unsigned(reg2376) : reg2066)));
                    end
                  reg2389 <= (reg2170 ~^ reg2144[(2'h3):(2'h3)]);
                  for (forvar2390 = (1'h0); (forvar2390 < (2'h3)); forvar2390 = (forvar2390 + (1'h1)))
                    begin
                      reg2391 <= reg2097[(4'hf):(4'hc)];
                      reg2392 <= ($unsigned(reg2109[(3'h5):(2'h3)]) ?
                          reg2223 : reg2331);
                    end
                end
            end
        end
    end
  module2393 #() modinst2503 (.wire2394(reg2251), .wire2395(reg2289), .wire2396(reg2094), .clk(clk), .wire2397(reg2154), .wire2398(reg2198), .y(wire2502));
  assign wire2504 = reg2233[(2'h3):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar2505 = (1'h0); (forvar2505 < (2'h3)); forvar2505 = (forvar2505 + (1'h1)))
        begin
          if (reg2199)
            begin
              for (forvar2506 = (1'h0); (forvar2506 < (2'h3)); forvar2506 = (forvar2506 + (1'h1)))
                begin
                  if ((-{$signed(reg2156[(4'hd):(4'ha)])}))
                    begin
                      reg2507 <= {reg2198[(3'h5):(3'h5)]};
                      reg2508 <= $signed({reg2206[(1'h1):(1'h1)]});
                      reg2509 <= $signed((+(~^reg2152[(1'h1):(1'h0)])));
                      reg2510 <= reg2232[(4'he):(1'h0)];
                    end
                  else
                    begin
                      reg2507 <= ({{(reg2315 ~^ reg2277)}} ?
                          {reg2186} : $signed((&(reg2183 ?
                              reg2306 : (8'hb6)))));
                    end
                  for (forvar2511 = (1'h0); (forvar2511 < (2'h3)); forvar2511 = (forvar2511 + (1'h1)))
                    begin
                      reg2512 <= $unsigned((~reg2281[(1'h1):(1'h1)]));
                      reg2513 <= (reg2348[(2'h2):(2'h2)] ? reg2249 : reg2306);
                    end
                end
              reg2514 <= ($signed(reg2307) ?
                  $unsigned($signed(reg2156)) : reg2228);
              for (forvar2515 = (1'h0); (forvar2515 < (2'h3)); forvar2515 = (forvar2515 + (1'h1)))
                begin
                  for (forvar2516 = (1'h0); (forvar2516 < (2'h3)); forvar2516 = (forvar2516 + (1'h1)))
                    begin
                      reg2517 <= reg2258;
                      reg2518 <= ({$unsigned(reg2309[(1'h0):(1'h0)])} ?
                          reg2264 : $signed(reg2367[(3'h4):(2'h2)]));
                    end
                end
            end
          else
            begin
              for (forvar2506 = (1'h0); (forvar2506 < (2'h3)); forvar2506 = (forvar2506 + (1'h1)))
                begin
                  if (reg2262[(3'h6):(2'h3)])
                    begin
                      reg2507 <= {$signed(reg2064)};
                      reg2508 <= (+(|($signed(reg2132) ?
                          reg2354 : (!reg2313))));
                    end
                  else
                    begin
                      reg2507 <= ($signed($unsigned($unsigned(reg2275))) ~^ (8'h9f));
                      reg2508 <= reg2130;
                      reg2509 <= ($signed((-$unsigned(reg2096))) ?
                          (reg2327 == reg2222[(2'h3):(2'h3)]) : $signed($unsigned(((8'ha5) <<< reg2286))));
                    end
                  reg2510 <= reg2130[(4'h8):(3'h5)];
                end
              for (forvar2511 = (1'h0); (forvar2511 < (1'h1)); forvar2511 = (forvar2511 + (1'h1)))
                begin
                  for (forvar2512 = (1'h0); (forvar2512 < (1'h0)); forvar2512 = (forvar2512 + (1'h1)))
                    begin
                      reg2513 <= ({{reg2324}} & (^~(+(reg2389 != reg2229))));
                    end
                  for (forvar2514 = (1'h0); (forvar2514 < (1'h1)); forvar2514 = (forvar2514 + (1'h1)))
                    begin
                      reg2515 <= ($signed((reg2249 > $unsigned(reg2386))) ?
                          ({{reg2291}} ^ reg2283) : ($signed(((8'hba) ?
                                  reg2382 : reg2251)) ?
                              {((8'hb2) >= reg2313)} : $unsigned($signed(reg2386))));
                    end
                  for (forvar2516 = (1'h0); (forvar2516 < (2'h2)); forvar2516 = (forvar2516 + (1'h1)))
                    begin
                      reg2517 <= reg2274;
                      reg2518 <= ($unsigned(({reg2077} << $unsigned(reg2107))) * (^$unsigned((reg2144 > (8'ha8)))));
                      reg2519 <= (|((~^(reg2301 ? reg2267 : wire2040)) ?
                          reg2319[(2'h2):(1'h0)] : $signed(reg2115)));
                      reg2520 <= reg2178[(1'h0):(1'h0)];
                    end
                end
              if ($signed((~^$unsigned($signed((8'hb4))))))
                begin
                  for (forvar2521 = (1'h0); (forvar2521 < (2'h3)); forvar2521 = (forvar2521 + (1'h1)))
                    begin
                      reg2522 <= {$unsigned(reg2257[(1'h1):(1'h1)])};
                      reg2523 <= $signed(reg2345[(1'h0):(1'h0)]);
                      reg2524 <= {$unsigned($unsigned(reg2387))};
                      reg2525 <= ({{reg2175}} ?
                          {$signed(reg2156)} : ((reg2197[(2'h2):(1'h0)] ?
                              $signed(reg2391) : (&reg2079)) >= $signed((reg2173 ?
                              reg2282 : reg2152))));
                    end
                end
              else
                begin
                  reg2521 <= $signed(reg2508[(1'h0):(1'h0)]);
                  reg2522 <= (((-reg2262) ?
                          $signed((reg2376 ? reg2077 : reg2121)) : (-reg2377)) ?
                      (((reg2156 ? (8'ha9) : reg2052) || $signed(reg2383)) ?
                          ((reg2152 << reg2249) ?
                              (reg2245 || reg2195) : (reg2209 ?
                                  reg2056 : reg2293)) : $unsigned((reg2081 >= (8'had)))) : $signed((8'hb4)));
                end
            end
        end
      for (forvar2526 = (1'h0); (forvar2526 < (1'h1)); forvar2526 = (forvar2526 + (1'h1)))
        begin
          if ($unsigned(reg2372[(3'h6):(1'h1)]))
            begin
              if (($signed(reg2130) ?
                  $unsigned((8'hb7)) : (^($unsigned(reg2083) >>> (reg2123 ?
                      reg2129 : (8'had))))))
                begin
                  for (forvar2527 = (1'h0); (forvar2527 < (2'h2)); forvar2527 = (forvar2527 + (1'h1)))
                    begin
                      reg2528 <= (forvar2505[(3'h4):(2'h3)] * reg2142);
                    end
                  if (reg2155)
                    begin
                      reg2529 <= $unsigned(((~^reg2271) | $signed({(8'hac)})));
                      reg2530 <= $signed(wire2234);
                    end
                  else
                    begin
                      reg2529 <= {$unsigned(reg2048[(3'h4):(1'h1)])};
                    end
                  for (forvar2531 = (1'h0); (forvar2531 < (2'h3)); forvar2531 = (forvar2531 + (1'h1)))
                    begin
                      reg2532 <= reg2524;
                    end
                end
              else
                begin
                  reg2527 <= reg2328;
                  if ((~$unsigned($unsigned((reg2518 ? reg2051 : reg2201)))))
                    begin
                      reg2528 <= reg2108;
                      reg2529 <= $signed(((!reg2085[(2'h2):(1'h0)]) ?
                          reg2241[(3'h7):(1'h0)] : reg2201));
                      reg2530 <= reg2324[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2528 <= $signed((+($unsigned(reg2280) ?
                          (reg2532 ? reg2194 : reg2050) : (reg2508 ?
                              reg2185 : reg2076))));
                      reg2529 <= (($signed($unsigned(reg2276)) >>> reg2370[(1'h0):(1'h0)]) ?
                          $signed((reg2334 ?
                              $unsigned(reg2283) : (reg2278 + reg2169))) : (&(~|reg2509[(3'h7):(3'h4)])));
                      reg2530 <= (-((((8'hb1) ^ reg2100) ?
                              ((8'h9f) <= reg2154) : (reg2183 ?
                                  (8'ha7) : reg2232)) ?
                          (|reg2179[(4'ha):(3'h4)]) : ($signed(reg2524) ?
                              (forvar2521 ?
                                  reg2339 : reg2316) : reg2057[(1'h0):(1'h0)])));
                    end
                  if (({reg2129} ?
                      {$unsigned(reg2149[(3'h4):(1'h1)])} : $unsigned((8'hac))))
                    begin
                      reg2531 <= reg2241;
                    end
                  else
                    begin
                      reg2531 <= reg2312;
                    end
                  if ($unsigned({{(^reg2315)}}))
                    begin
                      reg2532 <= forvar2511;
                      reg2533 <= {($signed($unsigned(reg2071)) ?
                              reg2144 : {$signed((8'h9c))})};
                      reg2534 <= $signed($unsigned((-{reg2140})));
                      reg2535 <= ((~|reg2186[(3'h5):(3'h4)]) ~^ ((reg2350 != $signed((8'ha6))) ?
                          reg2311 : {reg2147[(2'h3):(2'h2)]}));
                    end
                  else
                    begin
                      reg2532 <= ((reg2293 ?
                          (reg2071 ?
                              (reg2355 ?
                                  reg2260 : reg2519) : reg2509) : wire2044) <= reg2244[(4'ha):(1'h1)]);
                      reg2533 <= $unsigned({($signed((8'ha8)) ?
                              (reg2065 * reg2389) : $signed((8'ha2)))});
                      reg2534 <= $signed($signed($signed((+reg2308))));
                    end
                end
              if (reg2145)
                begin
                  if ((|(((forvar2527 ?
                      reg2120 : reg2286) >= reg2210) && reg2346[(2'h2):(2'h2)])))
                    begin
                      reg2536 <= reg2074;
                      reg2537 <= reg2085;
                      reg2538 <= reg2142;
                      reg2539 <= $unsigned(reg2272);
                    end
                  else
                    begin
                      reg2536 <= reg2260;
                      reg2537 <= $signed(reg2155[(2'h2):(1'h1)]);
                    end
                end
              else
                begin
                  if ($unsigned($unsigned({$signed(reg2523)})))
                    begin
                      reg2536 <= $signed($unsigned(reg2266[(2'h2):(2'h2)]));
                      reg2537 <= {(-reg2268)};
                    end
                  else
                    begin
                      reg2536 <= $signed(($unsigned($unsigned(reg2259)) * ($signed((8'hae)) < reg2383)));
                      reg2537 <= (wire2235 ?
                          reg2514[(3'h5):(2'h2)] : $unsigned(((forvar2526 ?
                                  (8'hb0) : (8'haf)) ?
                              $signed(reg2226) : {reg2300})));
                    end
                  if ($signed((reg2174[(1'h1):(1'h1)] ?
                      $unsigned($unsigned(reg2214)) : $signed({wire2502}))))
                    begin
                      reg2538 <= ((forvar2505[(2'h2):(2'h2)] ?
                              ((-(8'ha9)) ?
                                  (reg2049 - reg2059) : {reg2276}) : reg2349[(1'h1):(1'h1)]) ?
                          ((~^(reg2288 ? reg2508 : reg2194)) ?
                              reg2113[(3'h7):(3'h4)] : $signed({reg2082})) : (reg2129[(2'h3):(1'h1)] ?
                              reg2319 : wire2235[(3'h4):(2'h2)]));
                      reg2539 <= $unsigned((!($unsigned(reg2072) == $signed(reg2389))));
                    end
                  else
                    begin
                      reg2538 <= (($signed($signed(reg2509)) <= reg2356) <= reg2327[(3'h4):(3'h4)]);
                      reg2539 <= (|$unsigned((reg2109 ?
                          {reg2517} : reg2055[(3'h5):(2'h3)])));
                      reg2540 <= $unsigned((reg2307 >= (!reg2061[(2'h3):(1'h1)])));
                      reg2541 <= reg2308[(2'h2):(1'h1)];
                    end
                  for (forvar2542 = (1'h0); (forvar2542 < (2'h2)); forvar2542 = (forvar2542 + (1'h1)))
                    begin
                      reg2543 <= $signed(reg2340[(3'h4):(2'h2)]);
                      reg2544 <= (reg2132[(2'h2):(2'h2)] <<< reg2538);
                      reg2545 <= (reg2265[(1'h1):(1'h1)] >>> ((reg2311 ?
                              (~|reg2199) : $unsigned(reg2307)) ?
                          reg2281 : (reg2293[(4'hd):(4'h9)] ?
                              {(8'h9d)} : $signed(reg2387))));
                    end
                  if ($signed(reg2166[(2'h3):(2'h2)]))
                    begin
                      reg2546 <= reg2229;
                      reg2547 <= $unsigned((reg2276 * (+$signed(reg2545))));
                      reg2548 <= reg2216;
                    end
                  else
                    begin
                      reg2546 <= (!(reg2282[(3'h4):(1'h1)] ^~ reg2269[(3'h6):(3'h5)]));
                      reg2547 <= $signed((reg2094 >>> (!(-(8'hae)))));
                      reg2548 <= ((8'h9e) ?
                          reg2339 : (reg2154 ^ $unsigned((reg2238 + reg2213))));
                      reg2549 <= ($signed((reg2324 ?
                          (reg2065 ? wire2043 : reg2529) : (reg2385 ?
                              reg2201 : (8'haa)))) * reg2180);
                    end
                end
            end
          else
            begin
              for (forvar2527 = (1'h0); (forvar2527 < (2'h3)); forvar2527 = (forvar2527 + (1'h1)))
                begin
                  for (forvar2528 = (1'h0); (forvar2528 < (1'h0)); forvar2528 = (forvar2528 + (1'h1)))
                    begin
                      reg2529 <= ((reg2256 ?
                              $unsigned(reg2531) : reg2059[(4'hc):(4'hb)]) ?
                          (forvar2531 - (8'h9d)) : reg2093);
                      reg2530 <= reg2122;
                    end
                  if (((8'ha9) ?
                      ((8'h9c) ?
                          (^(reg2288 ?
                              reg2106 : forvar2526)) : (8'ha8)) : $unsigned(reg2261)))
                    begin
                      reg2531 <= (8'h9c);
                      reg2532 <= $unsigned((~|$signed((reg2183 << reg2169))));
                      reg2533 <= ($signed($signed((reg2238 ?
                              reg2146 : reg2523))) ?
                          wire2235[(1'h1):(1'h1)] : (^~((reg2356 >>> reg2313) ?
                              $signed((8'hb3)) : $signed(reg2116))));
                    end
                  else
                    begin
                      reg2531 <= (-(8'ha7));
                      reg2532 <= ($signed({$signed(reg2188)}) & forvar2527[(3'h4):(1'h0)]);
                      reg2533 <= $signed(reg2199[(4'hd):(3'h7)]);
                    end
                  if (reg2255[(3'h4):(2'h3)])
                    begin
                      reg2534 <= reg2286;
                      reg2535 <= $signed(($unsigned((reg2183 ?
                              reg2316 : reg2191)) ?
                          {{reg2248}} : reg2335));
                      reg2536 <= $signed($signed($signed($unsigned((8'h9f)))));
                      reg2537 <= ($signed($unsigned((reg2373 ?
                          reg2528 : reg2302))) <<< (((reg2275 <<< reg2331) ?
                          (reg2096 > reg2534) : (|reg2152)) != (reg2328[(4'h9):(4'h8)] < $signed((8'ha5)))));
                    end
                  else
                    begin
                      reg2534 <= reg2244;
                      reg2535 <= ((((reg2382 ?
                              reg2142 : reg2109) != reg2099[(1'h1):(1'h0)]) <<< $unsigned((~&reg2335))) ?
                          ((reg2202 << (reg2060 ? (8'hb2) : (8'ha7))) ?
                              ((8'ha0) & $unsigned(reg2133)) : ($unsigned((8'ha7)) ?
                                  {reg2258} : $unsigned(reg2169))) : $unsigned($signed((reg2212 >= reg2280))));
                      reg2536 <= $signed((!$unsigned((!reg2281))));
                    end
                end
              reg2538 <= $unsigned((~^(wire2042[(2'h3):(1'h0)] ?
                  reg2541[(1'h1):(1'h1)] : (^~reg2085))));
              for (forvar2539 = (1'h0); (forvar2539 < (1'h0)); forvar2539 = (forvar2539 + (1'h1)))
                begin
                  if ((reg2183 ? reg2121 : reg2177))
                    begin
                      reg2540 <= (reg2247[(1'h1):(1'h1)] ?
                          (((!reg2117) >> (reg2386 ? reg2114 : reg2079)) ?
                              (~^((8'hb4) & (8'hb4))) : $unsigned($unsigned(reg2077))) : $unsigned((~&$unsigned(reg2185))));
                    end
                  else
                    begin
                      reg2540 <= reg2194;
                      reg2541 <= ((reg2376[(1'h0):(1'h0)] ?
                              (|reg2180) : {(+reg2266)}) ?
                          (reg2521 <<< (!(~|forvar2514))) : reg2146);
                      reg2542 <= $signed($unsigned($signed(reg2188[(3'h4):(2'h2)])));
                      reg2543 <= (~^(~(-(+reg2507))));
                    end
                  if (reg2376)
                    begin
                      reg2544 <= reg2312[(3'h6):(2'h2)];
                      reg2545 <= $unsigned(($unsigned((reg2358 ~^ reg2389)) > {(reg2151 ?
                              reg2218 : reg2277)}));
                      reg2546 <= $signed(reg2233[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg2544 <= $unsigned(reg2227);
                      reg2545 <= reg2047;
                      reg2546 <= (($unsigned((|reg2132)) ~^ $signed($signed(reg2197))) ?
                          $signed({$signed(reg2541)}) : {reg2160[(1'h0):(1'h0)]});
                    end
                  for (forvar2547 = (1'h0); (forvar2547 < (1'h0)); forvar2547 = (forvar2547 + (1'h1)))
                    begin
                      reg2548 <= reg2308[(4'he):(4'he)];
                    end
                end
              for (forvar2549 = (1'h0); (forvar2549 < (2'h2)); forvar2549 = (forvar2549 + (1'h1)))
                begin
                  if ((reg2064 <<< reg2057))
                    begin
                      reg2550 <= $unsigned((-(8'h9f)));
                      reg2551 <= $unsigned($signed(($unsigned(reg2183) > (reg2524 ~^ reg2264))));
                      reg2552 <= $signed($signed($signed(reg2302[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg2550 <= (~|($signed((reg2112 ?
                          reg2125 : reg2107)) < $unsigned(reg2251[(3'h4):(1'h1)])));
                    end
                  for (forvar2553 = (1'h0); (forvar2553 < (1'h1)); forvar2553 = (forvar2553 + (1'h1)))
                    begin
                      reg2554 <= reg2141[(3'h4):(3'h4)];
                    end
                end
            end
          for (forvar2555 = (1'h0); (forvar2555 < (1'h0)); forvar2555 = (forvar2555 + (1'h1)))
            begin
              if (((!(~|reg2387)) <= ((reg2180[(2'h2):(2'h2)] ?
                      $unsigned(reg2194) : (reg2527 & reg2093)) ?
                  (8'h9e) : (reg2554 ? (reg2242 <<< reg2277) : (8'hb4)))))
                begin
                  for (forvar2556 = (1'h0); (forvar2556 < (2'h3)); forvar2556 = (forvar2556 + (1'h1)))
                    begin
                      reg2557 <= (|$unsigned(forvar2505));
                      reg2558 <= $unsigned((~|$signed((reg2340 ?
                          (8'ha1) : reg2523))));
                      reg2559 <= $unsigned($unsigned(reg2116[(1'h1):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar2556 = (1'h0); (forvar2556 < (2'h3)); forvar2556 = (forvar2556 + (1'h1)))
                    begin
                      reg2557 <= (reg2115[(4'hc):(4'h8)] ?
                          $unsigned(reg2509[(2'h2):(1'h1)]) : (~^$unsigned((reg2146 <= reg2066))));
                      reg2558 <= {reg2216};
                    end
                  if ($signed(reg2348[(1'h1):(1'h0)]))
                    begin
                      reg2559 <= $signed(((reg2202 ?
                              {reg2128} : (reg2092 ? reg2066 : reg2123)) ?
                          $unsigned($unsigned(reg2287)) : (reg2349[(4'hb):(4'ha)] + (~|reg2294))));
                      reg2560 <= reg2160;
                    end
                  else
                    begin
                      reg2559 <= $signed($unsigned((reg2533[(1'h1):(1'h0)] - reg2299)));
                      reg2560 <= $unsigned(((^reg2333) ?
                          (reg2268[(2'h2):(1'h1)] ?
                              reg2051 : (reg2088 == reg2384)) : (~^reg2113[(4'ha):(4'h9)])));
                    end
                end
              for (forvar2561 = (1'h0); (forvar2561 < (1'h0)); forvar2561 = (forvar2561 + (1'h1)))
                begin
                  if ($unsigned({($signed(reg2149) < reg2336[(1'h1):(1'h1)])}))
                    begin
                      reg2562 <= reg2101[(1'h1):(1'h1)];
                      reg2563 <= reg2378;
                      reg2564 <= $signed((reg2557[(2'h2):(1'h0)] ?
                          (-reg2255[(4'hb):(4'hb)]) : $unsigned((8'hb4))));
                    end
                  else
                    begin
                      reg2562 <= (reg2544[(3'h4):(3'h4)] != (reg2212 & reg2560));
                    end
                end
              for (forvar2565 = (1'h0); (forvar2565 < (2'h2)); forvar2565 = (forvar2565 + (1'h1)))
                begin
                  for (forvar2566 = (1'h0); (forvar2566 < (2'h3)); forvar2566 = (forvar2566 + (1'h1)))
                    begin
                      reg2567 <= ((((+reg2528) ?
                          $signed((8'hb1)) : (~|reg2517)) | reg2362[(3'h4):(1'h1)]) - $unsigned(reg2292));
                    end
                end
              for (forvar2568 = (1'h0); (forvar2568 < (1'h1)); forvar2568 = (forvar2568 + (1'h1)))
                begin
                  reg2569 <= reg2550;
                  if (reg2513)
                    begin
                      reg2570 <= reg2224[(1'h1):(1'h1)];
                      reg2571 <= {reg2339};
                    end
                  else
                    begin
                      reg2570 <= $signed(reg2548[(3'h4):(3'h4)]);
                      reg2571 <= $unsigned($signed(($unsigned((8'ha9)) ?
                          reg2365[(1'h0):(1'h0)] : reg2145)));
                      reg2572 <= $unsigned(reg2316);
                    end
                  for (forvar2573 = (1'h0); (forvar2573 < (2'h3)); forvar2573 = (forvar2573 + (1'h1)))
                    begin
                      reg2574 <= (~reg2194[(4'hc):(3'h5)]);
                      reg2575 <= (((reg2232[(4'hb):(1'h0)] ?
                              reg2255[(3'h4):(3'h4)] : reg2283[(3'h4):(3'h4)]) ?
                          ((reg2217 ?
                              (8'hba) : reg2266) && forvar2573) : ((wire2235 ~^ (8'hb2)) ?
                              (reg2531 >>> reg2247) : (8'haa))) >= (&((^wire2042) ?
                          (reg2336 || reg2077) : reg2348)));
                      reg2576 <= {(~(reg2348 ?
                              reg2359[(4'h9):(4'h8)] : {reg2314}))};
                      reg2577 <= reg2100[(4'hb):(3'h6)];
                    end
                end
            end
        end
    end
  assign wire2578 = reg2114[(4'h8):(4'h8)];
  module2579 #() modinst3040 (.wire2581(reg2525), .wire2580(reg2367), .y(wire3039), .wire2583(reg2082), .wire2582(reg2269), .clk(clk));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2579  (y, clk, wire2583, wire2582, wire2581, wire2580);
  output wire [(32'h1496):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire2583;
  input wire [(4'hb):(1'h0)] wire2582;
  input wire signed [(2'h2):(1'h0)] wire2581;
  input wire signed [(4'he):(1'h0)] wire2580;
  wire signed [(4'hc):(1'h0)] wire3038;
  wire signed [(4'he):(1'h0)] wire2673;
  wire signed [(3'h4):(1'h0)] wire2672;
  wire [(3'h5):(1'h0)] wire2671;
  wire signed [(4'h8):(1'h0)] wire2670;
  wire signed [(3'h5):(1'h0)] wire2669;
  wire signed [(5'h10):(1'h0)] wire2668;
  wire signed [(2'h2):(1'h0)] wire2585;
  wire signed [(4'h8):(1'h0)] wire2584;
  reg [(4'hf):(1'h0)] reg3025 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3017 = (1'h0);
  reg [(2'h2):(1'h0)] reg3037 = (1'h0);
  reg [(2'h3):(1'h0)] reg3036 = (1'h0);
  reg [(3'h6):(1'h0)] reg3035 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3030 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3034 = (1'h0);
  reg [(4'hd):(1'h0)] reg3033 = (1'h0);
  reg [(4'h9):(1'h0)] reg3032 = (1'h0);
  reg [(4'hc):(1'h0)] reg3031 = (1'h0);
  reg [(2'h3):(1'h0)] reg3029 = (1'h0);
  reg [(4'hc):(1'h0)] reg3028 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3027 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3026 = (1'h0);
  reg [(5'h10):(1'h0)] reg3024 = (1'h0);
  reg [(3'h7):(1'h0)] reg3023 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3022 = (1'h0);
  reg [(4'ha):(1'h0)] reg3021 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3020 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3019 = (1'h0);
  reg [(2'h2):(1'h0)] reg3018 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3016 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3015 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3014 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3013 = (1'h0);
  reg [(3'h5):(1'h0)] reg2996 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2995 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2987 = (1'h0);
  reg [(4'h8):(1'h0)] reg2976 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3010 = (1'h0);
  reg [(4'hc):(1'h0)] reg3009 = (1'h0);
  reg [(3'h4):(1'h0)] reg3008 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3007 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3005 = (1'h0);
  reg [(4'h9):(1'h0)] reg3004 = (1'h0);
  reg [(4'ha):(1'h0)] reg3003 = (1'h0);
  reg [(4'he):(1'h0)] reg3002 = (1'h0);
  reg [(5'h10):(1'h0)] reg3001 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2999 = (1'h0);
  reg [(4'h8):(1'h0)] reg2998 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2997 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2994 = (1'h0);
  reg [(3'h5):(1'h0)] reg2993 = (1'h0);
  reg [(4'hb):(1'h0)] reg2992 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2991 = (1'h0);
  reg [(4'hf):(1'h0)] reg2990 = (1'h0);
  reg [(4'ha):(1'h0)] reg2989 = (1'h0);
  reg [(2'h2):(1'h0)] reg2988 = (1'h0);
  reg [(2'h2):(1'h0)] reg2986 = (1'h0);
  reg [(4'he):(1'h0)] reg2985 = (1'h0);
  reg [(3'h6):(1'h0)] reg2984 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2983 = (1'h0);
  reg [(4'hf):(1'h0)] reg2982 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2981 = (1'h0);
  reg [(4'h8):(1'h0)] reg2980 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2978 = (1'h0);
  reg [(3'h7):(1'h0)] reg2977 = (1'h0);
  reg [(4'hb):(1'h0)] reg2975 = (1'h0);
  reg [(4'hc):(1'h0)] reg2973 = (1'h0);
  reg [(3'h6):(1'h0)] reg2972 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2971 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2965 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2970 = (1'h0);
  reg [(4'hb):(1'h0)] reg2969 = (1'h0);
  reg [(4'hc):(1'h0)] reg2968 = (1'h0);
  reg [(4'h8):(1'h0)] reg2967 = (1'h0);
  reg [(2'h2):(1'h0)] reg2966 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2963 = (1'h0);
  reg [(4'hb):(1'h0)] reg2962 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2961 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2960 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2959 = (1'h0);
  reg [(4'hb):(1'h0)] reg2958 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2957 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2956 = (1'h0);
  reg [(4'hf):(1'h0)] reg2955 = (1'h0);
  reg [(2'h2):(1'h0)] reg2954 = (1'h0);
  reg [(4'hc):(1'h0)] reg2948 = (1'h0);
  reg [(4'ha):(1'h0)] reg2952 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2951 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2950 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2949 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2946 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2943 = (1'h0);
  reg [(4'hc):(1'h0)] reg2932 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2923 = (1'h0);
  reg [(3'h4):(1'h0)] reg2922 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2947 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2945 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2944 = (1'h0);
  reg [(2'h3):(1'h0)] reg2942 = (1'h0);
  reg [(4'hb):(1'h0)] reg2941 = (1'h0);
  reg [(4'ha):(1'h0)] reg2940 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2939 = (1'h0);
  reg [(3'h4):(1'h0)] reg2938 = (1'h0);
  reg [(4'h9):(1'h0)] reg2928 = (1'h0);
  reg [(2'h2):(1'h0)] reg2937 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2936 = (1'h0);
  reg [(4'h9):(1'h0)] reg2935 = (1'h0);
  reg [(3'h4):(1'h0)] reg2934 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2933 = (1'h0);
  reg [(2'h2):(1'h0)] reg2931 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2930 = (1'h0);
  reg [(3'h4):(1'h0)] reg2929 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2927 = (1'h0);
  reg [(3'h6):(1'h0)] reg2926 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2925 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2924 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2921 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2920 = (1'h0);
  reg [(3'h5):(1'h0)] reg2919 = (1'h0);
  reg [(2'h3):(1'h0)] reg2918 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2917 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2916 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2915 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2914 = (1'h0);
  reg [(2'h3):(1'h0)] reg2913 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2912 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2911 = (1'h0);
  reg [(3'h6):(1'h0)] reg2910 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2909 = (1'h0);
  reg [(4'ha):(1'h0)] reg2908 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2907 = (1'h0);
  reg [(3'h4):(1'h0)] reg2906 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2904 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2902 = (1'h0);
  reg [(3'h5):(1'h0)] reg2901 = (1'h0);
  reg [(4'hc):(1'h0)] reg2899 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2898 = (1'h0);
  reg [(4'hb):(1'h0)] reg2897 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2896 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2895 = (1'h0);
  reg [(4'hd):(1'h0)] reg2893 = (1'h0);
  reg [(4'h8):(1'h0)] reg2892 = (1'h0);
  reg [(4'he):(1'h0)] reg2891 = (1'h0);
  reg [(4'hb):(1'h0)] reg2890 = (1'h0);
  reg [(4'hf):(1'h0)] reg2887 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2886 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2885 = (1'h0);
  reg [(5'h10):(1'h0)] reg2884 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2881 = (1'h0);
  reg [(4'h9):(1'h0)] reg2867 = (1'h0);
  reg [(4'hb):(1'h0)] reg2865 = (1'h0);
  reg [(5'h10):(1'h0)] reg2862 = (1'h0);
  reg [(5'h10):(1'h0)] reg2853 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2852 = (1'h0);
  reg [(3'h4):(1'h0)] reg2847 = (1'h0);
  reg [(3'h6):(1'h0)] reg2826 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2820 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2812 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2807 = (1'h0);
  reg [(4'hc):(1'h0)] reg2782 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2879 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2878 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2877 = (1'h0);
  reg [(4'h8):(1'h0)] reg2876 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2874 = (1'h0);
  reg [(4'hc):(1'h0)] reg2873 = (1'h0);
  reg [(4'hf):(1'h0)] reg2872 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2871 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2869 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2868 = (1'h0);
  reg [(4'ha):(1'h0)] reg2866 = (1'h0);
  reg [(3'h7):(1'h0)] reg2863 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2861 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2860 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2859 = (1'h0);
  reg [(4'he):(1'h0)] reg2857 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2858 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2856 = (1'h0);
  reg [(4'h9):(1'h0)] reg2855 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2854 = (1'h0);
  reg [(2'h2):(1'h0)] reg2851 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2850 = (1'h0);
  reg [(4'hd):(1'h0)] reg2849 = (1'h0);
  reg [(4'ha):(1'h0)] reg2848 = (1'h0);
  reg [(3'h5):(1'h0)] reg2846 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2845 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2844 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2840 = (1'h0);
  reg [(4'ha):(1'h0)] reg2837 = (1'h0);
  reg [(2'h3):(1'h0)] reg2843 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2842 = (1'h0);
  reg [(3'h7):(1'h0)] reg2841 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2839 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2838 = (1'h0);
  reg [(3'h4):(1'h0)] reg2836 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2835 = (1'h0);
  reg [(4'ha):(1'h0)] reg2834 = (1'h0);
  reg [(4'h8):(1'h0)] reg2833 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2832 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2831 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2830 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2829 = (1'h0);
  reg [(3'h4):(1'h0)] reg2828 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2821 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2827 = (1'h0);
  reg [(3'h4):(1'h0)] reg2825 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2824 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2823 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2822 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2819 = (1'h0);
  reg [(3'h5):(1'h0)] reg2777 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2818 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2817 = (1'h0);
  reg [(4'hc):(1'h0)] reg2816 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2815 = (1'h0);
  reg [(4'hb):(1'h0)] reg2814 = (1'h0);
  reg [(4'ha):(1'h0)] reg2813 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2811 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2810 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2809 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2808 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2806 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2805 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2804 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2803 = (1'h0);
  reg [(4'hc):(1'h0)] reg2802 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2801 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2796 = (1'h0);
  reg [(2'h2):(1'h0)] reg2800 = (1'h0);
  reg [(3'h5):(1'h0)] reg2799 = (1'h0);
  reg [(3'h7):(1'h0)] reg2798 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2797 = (1'h0);
  reg [(2'h3):(1'h0)] reg2795 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2794 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2793 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2792 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2791 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2790 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2789 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2788 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2787 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2786 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2785 = (1'h0);
  reg [(4'h8):(1'h0)] reg2784 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2783 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2781 = (1'h0);
  reg [(3'h5):(1'h0)] reg2780 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2779 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2778 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2776 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2775 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2774 = (1'h0);
  reg [(4'he):(1'h0)] reg2773 = (1'h0);
  reg [(3'h6):(1'h0)] reg2772 = (1'h0);
  reg [(4'he):(1'h0)] reg2771 = (1'h0);
  reg [(3'h7):(1'h0)] reg2770 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2768 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2767 = (1'h0);
  reg [(4'ha):(1'h0)] reg2766 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2765 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2751 = (1'h0);
  reg [(4'hc):(1'h0)] reg2750 = (1'h0);
  reg [(5'h10):(1'h0)] reg2763 = (1'h0);
  reg [(4'ha):(1'h0)] reg2761 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2759 = (1'h0);
  reg [(4'h9):(1'h0)] reg2762 = (1'h0);
  reg [(4'hb):(1'h0)] reg2760 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2758 = (1'h0);
  reg [(3'h5):(1'h0)] reg2757 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2756 = (1'h0);
  reg [(5'h10):(1'h0)] reg2755 = (1'h0);
  reg [(4'hd):(1'h0)] reg2754 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2753 = (1'h0);
  reg [(4'h9):(1'h0)] reg2752 = (1'h0);
  reg [(3'h4):(1'h0)] reg2749 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2748 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2747 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2743 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2746 = (1'h0);
  reg [(4'hc):(1'h0)] reg2745 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2744 = (1'h0);
  reg [(4'hd):(1'h0)] reg2742 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2741 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2740 = (1'h0);
  reg [(4'he):(1'h0)] reg2739 = (1'h0);
  reg [(4'ha):(1'h0)] reg2738 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2737 = (1'h0);
  reg [(4'h8):(1'h0)] reg2736 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2735 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2734 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2733 = (1'h0);
  reg [(2'h2):(1'h0)] reg2731 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2730 = (1'h0);
  reg [(3'h7):(1'h0)] reg2729 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2700 = (1'h0);
  reg [(5'h10):(1'h0)] reg2707 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2704 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2701 = (1'h0);
  reg [(4'hc):(1'h0)] reg2698 = (1'h0);
  reg [(4'h9):(1'h0)] reg2694 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2692 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2728 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2727 = (1'h0);
  reg [(4'he):(1'h0)] reg2726 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2725 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2724 = (1'h0);
  reg [(4'hf):(1'h0)] reg2718 = (1'h0);
  reg [(2'h3):(1'h0)] reg2706 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2712 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2723 = (1'h0);
  reg [(3'h4):(1'h0)] reg2722 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2721 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2720 = (1'h0);
  reg [(4'h9):(1'h0)] reg2719 = (1'h0);
  reg [(4'ha):(1'h0)] reg2717 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2716 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2715 = (1'h0);
  reg [(4'h8):(1'h0)] reg2714 = (1'h0);
  reg [(3'h5):(1'h0)] reg2713 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2711 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2710 = (1'h0);
  reg [(4'h8):(1'h0)] reg2709 = (1'h0);
  reg [(4'ha):(1'h0)] reg2708 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2705 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2703 = (1'h0);
  reg [(3'h7):(1'h0)] reg2702 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2699 = (1'h0);
  reg [(2'h3):(1'h0)] reg2697 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2696 = (1'h0);
  reg [(3'h6):(1'h0)] reg2695 = (1'h0);
  reg [(4'he):(1'h0)] reg2693 = (1'h0);
  reg [(4'h8):(1'h0)] reg2684 = (1'h0);
  reg [(4'hc):(1'h0)] reg2691 = (1'h0);
  reg [(2'h2):(1'h0)] reg2690 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2687 = (1'h0);
  reg [(3'h5):(1'h0)] reg2686 = (1'h0);
  reg [(4'hf):(1'h0)] reg2685 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2683 = (1'h0);
  reg [(4'hc):(1'h0)] reg2682 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2681 = (1'h0);
  reg [(2'h3):(1'h0)] reg2678 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2667 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2666 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2661 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2664 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2663 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2662 = (1'h0);
  reg [(4'h9):(1'h0)] reg2660 = (1'h0);
  reg [(4'h8):(1'h0)] reg2659 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2658 = (1'h0);
  reg [(4'ha):(1'h0)] reg2650 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2657 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2656 = (1'h0);
  reg [(3'h4):(1'h0)] reg2655 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2654 = (1'h0);
  reg [(4'he):(1'h0)] reg2653 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2652 = (1'h0);
  reg [(2'h3):(1'h0)] reg2651 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2649 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2648 = (1'h0);
  reg [(4'ha):(1'h0)] reg2646 = (1'h0);
  reg [(4'hd):(1'h0)] reg2645 = (1'h0);
  reg [(4'h9):(1'h0)] reg2644 = (1'h0);
  reg [(2'h3):(1'h0)] reg2642 = (1'h0);
  reg [(3'h6):(1'h0)] reg2641 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2640 = (1'h0);
  reg [(4'hd):(1'h0)] reg2639 = (1'h0);
  reg [(3'h7):(1'h0)] reg2636 = (1'h0);
  reg [(2'h3):(1'h0)] reg2635 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2634 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2633 = (1'h0);
  reg [(3'h7):(1'h0)] reg2632 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2631 = (1'h0);
  reg [(4'h9):(1'h0)] reg2630 = (1'h0);
  reg [(2'h2):(1'h0)] reg2629 = (1'h0);
  reg [(4'hb):(1'h0)] reg2628 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2627 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2625 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2623 = (1'h0);
  reg [(3'h4):(1'h0)] reg2622 = (1'h0);
  reg [(4'h9):(1'h0)] reg2621 = (1'h0);
  reg [(4'hc):(1'h0)] reg2620 = (1'h0);
  reg [(2'h2):(1'h0)] reg2619 = (1'h0);
  reg [(4'hc):(1'h0)] reg2618 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2616 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2609 = (1'h0);
  reg [(4'he):(1'h0)] reg2604 = (1'h0);
  reg [(4'hc):(1'h0)] reg2602 = (1'h0);
  reg [(4'hb):(1'h0)] reg2617 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2615 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2614 = (1'h0);
  reg [(4'ha):(1'h0)] reg2613 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2612 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2611 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2610 = (1'h0);
  reg [(5'h10):(1'h0)] reg2608 = (1'h0);
  reg [(3'h5):(1'h0)] reg2607 = (1'h0);
  reg [(4'hc):(1'h0)] reg2606 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2605 = (1'h0);
  reg [(4'hd):(1'h0)] reg2603 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2600 = (1'h0);
  reg [(5'h10):(1'h0)] reg2599 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2598 = (1'h0);
  reg [(4'hf):(1'h0)] reg2597 = (1'h0);
  reg [(2'h2):(1'h0)] reg2596 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2595 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2594 = (1'h0);
  reg [(4'hb):(1'h0)] reg2593 = (1'h0);
  reg [(4'hf):(1'h0)] reg2592 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2591 = (1'h0);
  reg [(2'h2):(1'h0)] reg2590 = (1'h0);
  reg [(3'h4):(1'h0)] reg2589 = (1'h0);
  reg [(4'h9):(1'h0)] reg2588 = (1'h0);
  reg [(2'h3):(1'h0)] reg2587 = (1'h0);
  reg [(2'h3):(1'h0)] reg2586 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3026 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3021 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3016 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3015 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3034 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3030 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3025 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3017 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3012 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3011 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2994 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2989 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2988 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2975 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3006 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3000 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2996 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2995 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2987 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2979 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2976 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2974 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2966 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2968 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2965 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2964 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2953 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2948 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2944 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2942 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2938 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2945 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2941 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2935 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2925 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2929 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2918 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2917 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2911 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2946 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2943 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2936 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2934 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2927 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2932 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2928 = (1'h0);
  reg [(4'he):(1'h0)] forvar2923 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2922 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2915 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2905 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2903 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2900 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2894 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2889 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2888 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2883 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2882 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2880 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2859 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2854 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2849 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2843 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2834 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2833 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2816 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2813 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2811 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2827 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2818 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2805 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2814 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2809 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2803 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2800 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2793 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2789 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2784 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2779 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2877 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2875 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2870 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2867 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2865 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2864 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2862 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2858 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2857 = (1'h0);
  reg [(4'he):(1'h0)] forvar2853 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2852 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2847 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2841 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2840 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2837 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2822 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2826 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2821 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2820 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2774 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2773 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2812 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2807 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2799 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2796 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2792 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2790 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2787 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2782 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2777 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2769 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2764 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2760 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2754 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2753 = (1'h0);
  reg [(4'he):(1'h0)] forvar2761 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2759 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2751 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2750 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2740 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2743 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2732 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2727 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2726 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2725 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2722 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2720 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2709 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2705 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2696 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2714 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2710 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2703 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2702 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2697 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2693 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2719 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2716 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2711 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2718 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2712 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2707 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2706 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2704 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2701 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2700 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2698 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2694 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2692 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2689 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2688 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2684 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2680 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2679 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2677 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2676 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2675 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2674 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2596 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2591 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2588 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2665 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2660 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2661 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2653 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2648 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2650 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2647 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2643 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2638 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2637 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2626 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2624 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2615 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2605 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2600 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2616 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2609 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2604 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2602 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2601 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2595 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2594 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2586 = (1'h0);
  assign y = {wire3038,
                 wire2673,
                 wire2672,
                 wire2671,
                 wire2670,
                 wire2669,
                 wire2668,
                 wire2585,
                 wire2584,
                 reg3025,
                 reg3017,
                 reg3037,
                 reg3036,
                 reg3035,
                 reg3030,
                 reg3034,
                 reg3033,
                 reg3032,
                 reg3031,
                 reg3029,
                 reg3028,
                 reg3027,
                 reg3026,
                 reg3024,
                 reg3023,
                 reg3022,
                 reg3021,
                 reg3020,
                 reg3019,
                 reg3018,
                 reg3016,
                 reg3015,
                 reg3014,
                 reg3013,
                 reg2996,
                 reg2995,
                 reg2987,
                 reg2976,
                 reg3010,
                 reg3009,
                 reg3008,
                 reg3007,
                 reg3005,
                 reg3004,
                 reg3003,
                 reg3002,
                 reg3001,
                 reg2999,
                 reg2998,
                 reg2997,
                 reg2994,
                 reg2993,
                 reg2992,
                 reg2991,
                 reg2990,
                 reg2989,
                 reg2988,
                 reg2986,
                 reg2985,
                 reg2984,
                 reg2983,
                 reg2982,
                 reg2981,
                 reg2980,
                 reg2978,
                 reg2977,
                 reg2975,
                 reg2973,
                 reg2972,
                 reg2971,
                 reg2965,
                 reg2970,
                 reg2969,
                 reg2968,
                 reg2967,
                 reg2966,
                 reg2963,
                 reg2962,
                 reg2961,
                 reg2960,
                 reg2959,
                 reg2958,
                 reg2957,
                 reg2956,
                 reg2955,
                 reg2954,
                 reg2948,
                 reg2952,
                 reg2951,
                 reg2950,
                 reg2949,
                 reg2946,
                 reg2943,
                 reg2932,
                 reg2923,
                 reg2922,
                 reg2947,
                 reg2945,
                 reg2944,
                 reg2942,
                 reg2941,
                 reg2940,
                 reg2939,
                 reg2938,
                 reg2928,
                 reg2937,
                 reg2936,
                 reg2935,
                 reg2934,
                 reg2933,
                 reg2931,
                 reg2930,
                 reg2929,
                 reg2927,
                 reg2926,
                 reg2925,
                 reg2924,
                 reg2921,
                 reg2920,
                 reg2919,
                 reg2918,
                 reg2917,
                 reg2916,
                 reg2915,
                 reg2914,
                 reg2913,
                 reg2912,
                 reg2911,
                 reg2910,
                 reg2909,
                 reg2908,
                 reg2907,
                 reg2906,
                 reg2904,
                 reg2902,
                 reg2901,
                 reg2899,
                 reg2898,
                 reg2897,
                 reg2896,
                 reg2895,
                 reg2893,
                 reg2892,
                 reg2891,
                 reg2890,
                 reg2887,
                 reg2886,
                 reg2885,
                 reg2884,
                 reg2881,
                 reg2867,
                 reg2865,
                 reg2862,
                 reg2853,
                 reg2852,
                 reg2847,
                 reg2826,
                 reg2820,
                 reg2812,
                 reg2807,
                 reg2782,
                 reg2879,
                 reg2878,
                 reg2877,
                 reg2876,
                 reg2874,
                 reg2873,
                 reg2872,
                 reg2871,
                 reg2869,
                 reg2868,
                 reg2866,
                 reg2863,
                 reg2861,
                 reg2860,
                 reg2859,
                 reg2857,
                 reg2858,
                 reg2856,
                 reg2855,
                 reg2854,
                 reg2851,
                 reg2850,
                 reg2849,
                 reg2848,
                 reg2846,
                 reg2845,
                 reg2844,
                 reg2840,
                 reg2837,
                 reg2843,
                 reg2842,
                 reg2841,
                 reg2839,
                 reg2838,
                 reg2836,
                 reg2835,
                 reg2834,
                 reg2833,
                 reg2832,
                 reg2831,
                 reg2830,
                 reg2829,
                 reg2828,
                 reg2821,
                 reg2827,
                 reg2825,
                 reg2824,
                 reg2823,
                 reg2822,
                 reg2819,
                 reg2777,
                 reg2818,
                 reg2817,
                 reg2816,
                 reg2815,
                 reg2814,
                 reg2813,
                 reg2811,
                 reg2810,
                 reg2809,
                 reg2808,
                 reg2806,
                 reg2805,
                 reg2804,
                 reg2803,
                 reg2802,
                 reg2801,
                 reg2796,
                 reg2800,
                 reg2799,
                 reg2798,
                 reg2797,
                 reg2795,
                 reg2794,
                 reg2793,
                 reg2792,
                 reg2791,
                 reg2790,
                 reg2789,
                 reg2788,
                 reg2787,
                 reg2786,
                 reg2785,
                 reg2784,
                 reg2783,
                 reg2781,
                 reg2780,
                 reg2779,
                 reg2778,
                 reg2776,
                 reg2775,
                 reg2774,
                 reg2773,
                 reg2772,
                 reg2771,
                 reg2770,
                 reg2768,
                 reg2767,
                 reg2766,
                 reg2765,
                 reg2751,
                 reg2750,
                 reg2763,
                 reg2761,
                 reg2759,
                 reg2762,
                 reg2760,
                 reg2758,
                 reg2757,
                 reg2756,
                 reg2755,
                 reg2754,
                 reg2753,
                 reg2752,
                 reg2749,
                 reg2748,
                 reg2747,
                 reg2743,
                 reg2746,
                 reg2745,
                 reg2744,
                 reg2742,
                 reg2741,
                 reg2740,
                 reg2739,
                 reg2738,
                 reg2737,
                 reg2736,
                 reg2735,
                 reg2734,
                 reg2733,
                 reg2731,
                 reg2730,
                 reg2729,
                 reg2700,
                 reg2707,
                 reg2704,
                 reg2701,
                 reg2698,
                 reg2694,
                 reg2692,
                 reg2728,
                 reg2727,
                 reg2726,
                 reg2725,
                 reg2724,
                 reg2718,
                 reg2706,
                 reg2712,
                 reg2723,
                 reg2722,
                 reg2721,
                 reg2720,
                 reg2719,
                 reg2717,
                 reg2716,
                 reg2715,
                 reg2714,
                 reg2713,
                 reg2711,
                 reg2710,
                 reg2709,
                 reg2708,
                 reg2705,
                 reg2703,
                 reg2702,
                 reg2699,
                 reg2697,
                 reg2696,
                 reg2695,
                 reg2693,
                 reg2684,
                 reg2691,
                 reg2690,
                 reg2687,
                 reg2686,
                 reg2685,
                 reg2683,
                 reg2682,
                 reg2681,
                 reg2678,
                 reg2667,
                 reg2666,
                 reg2661,
                 reg2664,
                 reg2663,
                 reg2662,
                 reg2660,
                 reg2659,
                 reg2658,
                 reg2650,
                 reg2657,
                 reg2656,
                 reg2655,
                 reg2654,
                 reg2653,
                 reg2652,
                 reg2651,
                 reg2649,
                 reg2648,
                 reg2646,
                 reg2645,
                 reg2644,
                 reg2642,
                 reg2641,
                 reg2640,
                 reg2639,
                 reg2636,
                 reg2635,
                 reg2634,
                 reg2633,
                 reg2632,
                 reg2631,
                 reg2630,
                 reg2629,
                 reg2628,
                 reg2627,
                 reg2625,
                 reg2623,
                 reg2622,
                 reg2621,
                 reg2620,
                 reg2619,
                 reg2618,
                 reg2616,
                 reg2609,
                 reg2604,
                 reg2602,
                 reg2617,
                 reg2615,
                 reg2614,
                 reg2613,
                 reg2612,
                 reg2611,
                 reg2610,
                 reg2608,
                 reg2607,
                 reg2606,
                 reg2605,
                 reg2603,
                 reg2600,
                 reg2599,
                 reg2598,
                 reg2597,
                 reg2596,
                 reg2595,
                 reg2594,
                 reg2593,
                 reg2592,
                 reg2591,
                 reg2590,
                 reg2589,
                 reg2588,
                 reg2587,
                 reg2586,
                 forvar3026,
                 forvar3021,
                 forvar3016,
                 forvar3015,
                 forvar3034,
                 forvar3030,
                 forvar3025,
                 forvar3017,
                 forvar3012,
                 forvar3011,
                 forvar2994,
                 forvar2989,
                 forvar2988,
                 forvar2975,
                 forvar3006,
                 forvar3000,
                 forvar2996,
                 forvar2995,
                 forvar2987,
                 forvar2979,
                 forvar2976,
                 forvar2974,
                 forvar2966,
                 forvar2968,
                 forvar2965,
                 forvar2964,
                 forvar2953,
                 forvar2948,
                 forvar2944,
                 forvar2942,
                 forvar2938,
                 forvar2945,
                 forvar2941,
                 forvar2935,
                 forvar2925,
                 forvar2929,
                 forvar2918,
                 forvar2917,
                 forvar2911,
                 forvar2946,
                 forvar2943,
                 forvar2936,
                 forvar2934,
                 forvar2927,
                 forvar2932,
                 forvar2928,
                 forvar2923,
                 forvar2922,
                 forvar2915,
                 forvar2905,
                 forvar2903,
                 forvar2900,
                 forvar2894,
                 forvar2889,
                 forvar2888,
                 forvar2883,
                 forvar2882,
                 forvar2880,
                 forvar2859,
                 forvar2854,
                 forvar2849,
                 forvar2843,
                 forvar2834,
                 forvar2833,
                 forvar2816,
                 forvar2813,
                 forvar2811,
                 forvar2827,
                 forvar2818,
                 forvar2805,
                 forvar2814,
                 forvar2809,
                 forvar2803,
                 forvar2800,
                 forvar2793,
                 forvar2789,
                 forvar2784,
                 forvar2779,
                 forvar2877,
                 forvar2875,
                 forvar2870,
                 forvar2867,
                 forvar2865,
                 forvar2864,
                 forvar2862,
                 forvar2858,
                 forvar2857,
                 forvar2853,
                 forvar2852,
                 forvar2847,
                 forvar2841,
                 forvar2840,
                 forvar2837,
                 forvar2822,
                 forvar2826,
                 forvar2821,
                 forvar2820,
                 forvar2774,
                 forvar2773,
                 forvar2812,
                 forvar2807,
                 forvar2799,
                 forvar2796,
                 forvar2792,
                 forvar2790,
                 forvar2787,
                 forvar2782,
                 forvar2777,
                 forvar2769,
                 forvar2764,
                 forvar2760,
                 forvar2754,
                 forvar2753,
                 forvar2761,
                 forvar2759,
                 forvar2751,
                 forvar2750,
                 forvar2740,
                 forvar2743,
                 forvar2732,
                 forvar2727,
                 forvar2726,
                 forvar2725,
                 forvar2722,
                 forvar2720,
                 forvar2709,
                 forvar2705,
                 forvar2696,
                 forvar2714,
                 forvar2710,
                 forvar2703,
                 forvar2702,
                 forvar2697,
                 forvar2693,
                 forvar2719,
                 forvar2716,
                 forvar2711,
                 forvar2718,
                 forvar2712,
                 forvar2707,
                 forvar2706,
                 forvar2704,
                 forvar2701,
                 forvar2700,
                 forvar2698,
                 forvar2694,
                 forvar2692,
                 forvar2689,
                 forvar2688,
                 forvar2684,
                 forvar2680,
                 forvar2679,
                 forvar2677,
                 forvar2676,
                 forvar2675,
                 forvar2674,
                 forvar2596,
                 forvar2591,
                 forvar2588,
                 forvar2665,
                 forvar2660,
                 forvar2661,
                 forvar2653,
                 forvar2648,
                 forvar2650,
                 forvar2647,
                 forvar2643,
                 forvar2638,
                 forvar2637,
                 forvar2626,
                 forvar2624,
                 forvar2615,
                 forvar2605,
                 forvar2600,
                 forvar2616,
                 forvar2609,
                 forvar2604,
                 forvar2602,
                 forvar2601,
                 forvar2595,
                 forvar2594,
                 forvar2586,
                 (1'h0)};
  assign wire2584 = (|wire2581);
  assign wire2585 = (~wire2580[(4'hc):(4'hc)]);
  always
    @(posedge clk) begin
      if ($unsigned((+$signed({(8'ha6)}))))
        begin
          if ($signed({((&wire2582) || $unsigned((8'hba)))}))
            begin
              if (wire2584)
                begin
                  if ($unsigned($unsigned($signed(wire2581))))
                    begin
                      reg2586 <= (^~{$unsigned(wire2584[(2'h2):(1'h0)])});
                      reg2587 <= (wire2581[(2'h2):(1'h0)] ?
                          wire2584[(1'h0):(1'h0)] : $signed(wire2584[(3'h4):(2'h3)]));
                      reg2588 <= $unsigned((wire2585[(1'h0):(1'h0)] ?
                          ($unsigned(wire2581) ?
                              $signed(wire2581) : (wire2582 ?
                                  wire2584 : wire2581)) : ((reg2587 ?
                              (8'hb7) : wire2585) || $unsigned(wire2581))));
                    end
                  else
                    begin
                      reg2586 <= $signed(wire2582);
                      reg2587 <= ((8'hb4) ?
                          ($signed(wire2580[(4'ha):(3'h6)]) - $unsigned(reg2588[(1'h0):(1'h0)])) : ((~|wire2583[(1'h1):(1'h0)]) ?
                              reg2588[(3'h6):(2'h2)] : ((~&wire2584) && (~reg2587))));
                    end
                  if ((-$unsigned($signed((wire2581 ? wire2580 : (8'hb6))))))
                    begin
                      reg2589 <= (~({(reg2586 * wire2584)} ?
                          ((wire2584 ?
                              wire2583 : wire2584) - reg2587) : reg2588[(1'h0):(1'h0)]));
                      reg2590 <= $unsigned($signed($unsigned((8'hb1))));
                    end
                  else
                    begin
                      reg2589 <= ({((wire2585 ?
                              (8'hba) : wire2580) * $unsigned(wire2585))} || $signed({wire2581[(1'h1):(1'h1)]}));
                      reg2590 <= ((((reg2589 ? wire2582 : reg2587) ?
                          $signed(wire2581) : {wire2581}) ~^ $signed((~|reg2589))) * $signed((wire2583[(2'h3):(1'h0)] ?
                          $signed(wire2584) : (!reg2590))));
                      reg2591 <= (reg2589[(2'h3):(2'h2)] | (reg2586 || {reg2588[(3'h5):(1'h1)]}));
                    end
                  if ((^((~^(~|reg2588)) ?
                      ((wire2580 >= reg2586) ^ reg2589) : {(wire2580 ?
                              reg2587 : reg2587)})))
                    begin
                      reg2592 <= $signed(reg2586);
                      reg2593 <= (reg2592 * wire2581);
                    end
                  else
                    begin
                      reg2592 <= $unsigned((-(8'hb9)));
                      reg2593 <= ((+((-reg2588) + wire2580[(4'he):(1'h0)])) && $unsigned((((8'ha8) || reg2586) ?
                          (reg2587 & wire2583) : $unsigned(reg2587))));
                      reg2594 <= reg2589[(2'h3):(1'h0)];
                      reg2595 <= $unsigned($unsigned((((8'ha4) ?
                              wire2585 : (8'hb2)) ?
                          (reg2586 ? wire2581 : reg2590) : {reg2590})));
                    end
                end
              else
                begin
                  reg2586 <= (-(~^(~|$unsigned(reg2595))));
                end
            end
          else
            begin
              for (forvar2586 = (1'h0); (forvar2586 < (1'h1)); forvar2586 = (forvar2586 + (1'h1)))
                begin
                  if ($unsigned(wire2583[(1'h0):(1'h0)]))
                    begin
                      reg2587 <= $signed($unsigned((reg2587[(1'h1):(1'h1)] ?
                          {reg2587} : $signed((8'hba)))));
                      reg2588 <= ($signed($signed($unsigned(wire2582))) ?
                          $unsigned({{wire2582}}) : $unsigned(wire2581[(1'h0):(1'h0)]));
                      reg2589 <= (($unsigned((~forvar2586)) >>> (wire2583[(2'h3):(1'h0)] >= $unsigned(wire2585))) << reg2587[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg2587 <= reg2591[(1'h1):(1'h1)];
                    end
                  if ((~|reg2589[(2'h3):(2'h3)]))
                    begin
                      reg2590 <= $unsigned(reg2588[(1'h0):(1'h0)]);
                      reg2591 <= {(^~forvar2586[(4'he):(3'h4)])};
                      reg2592 <= ((8'haa) ?
                          reg2592[(1'h1):(1'h0)] : forvar2586);
                    end
                  else
                    begin
                      reg2590 <= $unsigned($signed(($unsigned(wire2582) != (+reg2594))));
                      reg2591 <= (-reg2589[(2'h3):(2'h3)]);
                      reg2592 <= $signed($signed(reg2593[(4'ha):(3'h7)]));
                      reg2593 <= wire2583;
                    end
                end
              for (forvar2594 = (1'h0); (forvar2594 < (1'h1)); forvar2594 = (forvar2594 + (1'h1)))
                begin
                  for (forvar2595 = (1'h0); (forvar2595 < (2'h2)); forvar2595 = (forvar2595 + (1'h1)))
                    begin
                      reg2596 <= reg2589[(1'h0):(1'h0)];
                    end
                  if (($unsigned(reg2596) ^~ (&$unsigned({(8'ha9)}))))
                    begin
                      reg2597 <= reg2590[(1'h1):(1'h1)];
                      reg2598 <= reg2591[(4'hb):(3'h5)];
                      reg2599 <= reg2593[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg2597 <= forvar2595;
                      reg2598 <= reg2587;
                    end
                end
            end
          if ($signed($unsigned(($signed(wire2585) << (wire2585 ?
              forvar2595 : reg2592)))))
            begin
              reg2600 <= {(($signed(reg2591) ?
                      (~reg2599) : reg2593) ^ $signed((reg2596 ?
                      reg2594 : reg2593)))};
              for (forvar2601 = (1'h0); (forvar2601 < (1'h0)); forvar2601 = (forvar2601 + (1'h1)))
                begin
                  for (forvar2602 = (1'h0); (forvar2602 < (1'h1)); forvar2602 = (forvar2602 + (1'h1)))
                    begin
                      reg2603 <= {reg2592[(4'ha):(3'h4)]};
                    end
                  for (forvar2604 = (1'h0); (forvar2604 < (2'h2)); forvar2604 = (forvar2604 + (1'h1)))
                    begin
                      reg2605 <= $signed($unsigned(wire2581));
                      reg2606 <= $unsigned(reg2600[(2'h2):(1'h0)]);
                      reg2607 <= $signed((^~(~^(reg2594 ?
                          forvar2595 : reg2587))));
                    end
                end
              reg2608 <= forvar2586[(3'h6):(2'h2)];
              for (forvar2609 = (1'h0); (forvar2609 < (2'h2)); forvar2609 = (forvar2609 + (1'h1)))
                begin
                  reg2610 <= reg2603;
                  if (((+forvar2601[(4'h9):(3'h6)]) > $signed($unsigned((wire2580 ?
                      reg2607 : reg2599)))))
                    begin
                      reg2611 <= reg2605[(3'h5):(3'h5)];
                      reg2612 <= $unsigned((+($unsigned(reg2606) | (^~(8'hb6)))));
                      reg2613 <= $unsigned({({forvar2609} <= (wire2583 - wire2583))});
                    end
                  else
                    begin
                      reg2611 <= reg2607[(2'h3):(2'h2)];
                      reg2612 <= (($unsigned($signed((8'hab))) < (reg2591[(1'h1):(1'h0)] << {(8'ha1)})) ?
                          (((reg2599 ? forvar2595 : reg2598) ?
                              {reg2612} : (reg2593 ~^ reg2597)) * ((wire2583 - reg2600) ?
                              (reg2605 ? forvar2586 : (8'ha6)) : (reg2591 ?
                                  (8'had) : reg2592))) : reg2589);
                      reg2613 <= $unsigned($unsigned((^~(reg2594 ?
                          (8'hb3) : forvar2609))));
                    end
                  if ((|reg2587))
                    begin
                      reg2614 <= {$unsigned({$signed(forvar2595)})};
                    end
                  else
                    begin
                      reg2614 <= $signed((8'ha6));
                      reg2615 <= reg2589;
                    end
                  for (forvar2616 = (1'h0); (forvar2616 < (2'h2)); forvar2616 = (forvar2616 + (1'h1)))
                    begin
                      reg2617 <= $signed(reg2595);
                    end
                end
            end
          else
            begin
              for (forvar2600 = (1'h0); (forvar2600 < (2'h3)); forvar2600 = (forvar2600 + (1'h1)))
                begin
                  for (forvar2601 = (1'h0); (forvar2601 < (2'h2)); forvar2601 = (forvar2601 + (1'h1)))
                    begin
                      reg2602 <= $unsigned($signed($unsigned($signed(reg2607))));
                      reg2603 <= ($unsigned(reg2598[(4'h9):(2'h2)]) | ((-$unsigned(reg2598)) << (~|(reg2610 != wire2584))));
                      reg2604 <= $signed(wire2584);
                    end
                  for (forvar2605 = (1'h0); (forvar2605 < (1'h1)); forvar2605 = (forvar2605 + (1'h1)))
                    begin
                      reg2606 <= reg2595[(4'h8):(3'h6)];
                      reg2607 <= reg2606[(1'h1):(1'h0)];
                    end
                  if (forvar2616[(1'h1):(1'h0)])
                    begin
                      reg2608 <= wire2580;
                      reg2609 <= $unsigned(($signed((^reg2593)) || forvar2600));
                      reg2610 <= ($unsigned(({forvar2594} - (~forvar2604))) >>> {$signed((reg2614 >= forvar2604))});
                    end
                  else
                    begin
                      reg2608 <= ($unsigned(((|reg2596) | reg2598[(1'h1):(1'h0)])) == (((~reg2593) ?
                          reg2614 : (reg2586 == reg2589)) >= $signed(forvar2594[(3'h5):(2'h2)])));
                    end
                  if ($signed((reg2599 >>> ((reg2593 >> reg2614) ?
                      (-forvar2586) : $signed(forvar2586)))))
                    begin
                      reg2611 <= $unsigned($signed((wire2583 & (forvar2594 ?
                          reg2617 : reg2592))));
                      reg2612 <= ($signed($unsigned((reg2595 ?
                          reg2598 : reg2602))) ~^ (reg2590 && $unsigned($signed(forvar2586))));
                    end
                  else
                    begin
                      reg2611 <= {(!reg2587)};
                      reg2612 <= $signed((^$signed((wire2584 ?
                          (8'h9e) : reg2604))));
                      reg2613 <= reg2593;
                      reg2614 <= (({wire2585} ?
                          ((~wire2581) <<< $signed(reg2611)) : ($signed(forvar2595) > (wire2582 ?
                              reg2604 : reg2590))) | reg2615[(4'h8):(3'h4)]);
                    end
                end
              if ($signed(((reg2600[(3'h4):(1'h0)] - $unsigned(reg2600)) - reg2609[(2'h2):(1'h0)])))
                begin
                  for (forvar2615 = (1'h0); (forvar2615 < (1'h1)); forvar2615 = (forvar2615 + (1'h1)))
                    begin
                      reg2616 <= reg2589;
                      reg2617 <= $signed((wire2581[(1'h0):(1'h0)] ?
                          $unsigned(reg2589[(2'h2):(1'h1)]) : $signed($signed((8'ha6)))));
                      reg2618 <= (~|reg2617);
                      reg2619 <= reg2592;
                    end
                  if ((($signed((^~reg2588)) ?
                      (|$signed(forvar2586)) : (wire2583[(2'h2):(1'h1)] * (forvar2601 ^~ reg2615))) * $signed(reg2597[(4'hc):(4'hc)])))
                    begin
                      reg2620 <= $unsigned($signed($signed({reg2614})));
                      reg2621 <= reg2592[(3'h5):(1'h1)];
                      reg2622 <= $signed($signed((forvar2595 ?
                          (+forvar2616) : (+reg2614))));
                      reg2623 <= wire2584[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg2620 <= $unsigned(reg2608);
                      reg2621 <= wire2583;
                    end
                end
              else
                begin
                  reg2615 <= ((~|$signed((~^(8'hab)))) <= $unsigned($unsigned(reg2589[(2'h2):(2'h2)])));
                  for (forvar2616 = (1'h0); (forvar2616 < (2'h3)); forvar2616 = (forvar2616 + (1'h1)))
                    begin
                      reg2617 <= ((-$signed((&(8'hb0)))) ?
                          ($unsigned((reg2621 ? reg2623 : reg2616)) ?
                              $unsigned({reg2596}) : $signed(wire2581[(1'h1):(1'h0)])) : $signed($signed((reg2611 + (8'ha7)))));
                      reg2618 <= $signed((reg2596 ^ ((&forvar2594) ?
                          $unsigned(reg2586) : (reg2614 && reg2588))));
                    end
                  if (forvar2602[(2'h3):(2'h2)])
                    begin
                      reg2619 <= (|((~|reg2595) ~^ $signed(reg2603[(4'hb):(2'h2)])));
                      reg2620 <= ((8'h9c) ^ $signed($signed({reg2623})));
                    end
                  else
                    begin
                      reg2619 <= (8'ha3);
                      reg2620 <= ((~$signed(((8'ha4) ? wire2584 : reg2588))) ?
                          {forvar2609[(4'h8):(2'h2)]} : {forvar2586[(1'h0):(1'h0)]});
                      reg2621 <= $unsigned((~^forvar2595[(3'h6):(2'h3)]));
                    end
                end
              for (forvar2624 = (1'h0); (forvar2624 < (1'h0)); forvar2624 = (forvar2624 + (1'h1)))
                begin
                  reg2625 <= $unsigned((reg2599 ^ $unsigned(reg2612[(4'ha):(1'h1)])));
                  for (forvar2626 = (1'h0); (forvar2626 < (2'h2)); forvar2626 = (forvar2626 + (1'h1)))
                    begin
                      reg2627 <= $unsigned(($unsigned(reg2614) & (forvar2594[(2'h3):(2'h3)] >= ((8'hb4) <<< reg2594))));
                      reg2628 <= {(((reg2610 < (8'ha3)) ?
                                  wire2585[(1'h1):(1'h0)] : (forvar2602 + (8'ha0))) ?
                              $unsigned((reg2591 ^ reg2596)) : ((reg2606 ^~ (8'ha7)) != $unsigned((8'h9c))))};
                      reg2629 <= ((wire2584 ?
                          (+$unsigned(reg2602)) : $signed($signed(reg2628))) >> reg2599);
                      reg2630 <= $signed((({forvar2624} ~^ forvar2600) ?
                          ((reg2612 ?
                              reg2621 : reg2605) <<< $unsigned(reg2596)) : ((!reg2614) ?
                              reg2620 : (-reg2594))));
                    end
                  if ($signed((~^(+(reg2599 ? forvar2605 : reg2600)))))
                    begin
                      reg2631 <= reg2596[(2'h2):(2'h2)];
                      reg2632 <= {(!$unsigned({reg2605}))};
                    end
                  else
                    begin
                      reg2631 <= $signed($unsigned(reg2602));
                      reg2632 <= reg2595;
                    end
                  if ($signed((wire2581 ^~ (reg2587 ?
                      (wire2580 ? (8'hb1) : forvar2615) : (+wire2582)))))
                    begin
                      reg2633 <= (!$unsigned({((8'ha3) ? (8'hae) : reg2615)}));
                      reg2634 <= (($unsigned(reg2617[(2'h2):(2'h2)]) >>> reg2587[(2'h2):(2'h2)]) ?
                          (reg2590[(1'h1):(1'h0)] & $signed((reg2612 ?
                              reg2617 : reg2597))) : reg2598);
                      reg2635 <= {$signed($signed(((8'hac) ?
                              reg2628 : reg2631)))};
                      reg2636 <= ($signed(($unsigned((8'hb1)) ?
                          (reg2631 <<< (8'hb3)) : $signed(reg2596))) == {$unsigned((reg2590 + reg2609))});
                    end
                  else
                    begin
                      reg2633 <= (-{$signed(reg2635[(2'h3):(2'h2)])});
                      reg2634 <= $unsigned((($unsigned(wire2585) < $signed(reg2596)) ^ reg2634[(3'h4):(2'h2)]));
                    end
                end
              for (forvar2637 = (1'h0); (forvar2637 < (1'h0)); forvar2637 = (forvar2637 + (1'h1)))
                begin
                  for (forvar2638 = (1'h0); (forvar2638 < (1'h0)); forvar2638 = (forvar2638 + (1'h1)))
                    begin
                      reg2639 <= forvar2595;
                      reg2640 <= reg2610[(4'hf):(3'h5)];
                    end
                  if ((8'h9c))
                    begin
                      reg2641 <= ((&(~^reg2592[(3'h5):(3'h5)])) >>> $unsigned(((reg2623 ?
                          forvar2601 : reg2625) - {reg2602})));
                      reg2642 <= ((forvar2601[(4'hb):(1'h0)] > reg2595) ?
                          (reg2612 >>> $signed($signed(forvar2586))) : $unsigned(reg2600[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg2641 <= wire2585[(1'h1):(1'h1)];
                      reg2642 <= (reg2605 ? (-reg2614) : reg2593);
                    end
                  for (forvar2643 = (1'h0); (forvar2643 < (2'h3)); forvar2643 = (forvar2643 + (1'h1)))
                    begin
                      reg2644 <= ({((reg2622 <<< wire2581) ?
                              forvar2643[(4'h9):(3'h5)] : {reg2592})} ^ $unsigned($unsigned($signed((8'had)))));
                      reg2645 <= $signed((forvar2604 | (wire2582[(1'h1):(1'h0)] ?
                          {reg2613} : (+reg2630))));
                      reg2646 <= (8'hb3);
                    end
                end
            end
          for (forvar2647 = (1'h0); (forvar2647 < (1'h0)); forvar2647 = (forvar2647 + (1'h1)))
            begin
              if ((8'haa))
                begin
                  if (($unsigned($unsigned((reg2603 ? reg2608 : reg2596))) ?
                      $unsigned($signed(((8'h9f) - reg2632))) : ($unsigned(forvar2615) ?
                          (8'hb9) : wire2583[(2'h2):(2'h2)])))
                    begin
                      reg2648 <= reg2641[(3'h4):(1'h1)];
                      reg2649 <= (~&wire2580[(4'hb):(1'h0)]);
                    end
                  else
                    begin
                      reg2648 <= ($unsigned($unsigned($signed((8'ha1)))) ?
                          (((&(8'hb3)) + $signed(reg2646)) ^~ $unsigned(reg2640[(2'h3):(1'h0)])) : (-{((8'hb5) ?
                                  reg2611 : reg2604)}));
                    end
                  for (forvar2650 = (1'h0); (forvar2650 < (2'h2)); forvar2650 = (forvar2650 + (1'h1)))
                    begin
                      reg2651 <= (!reg2588[(3'h4):(1'h0)]);
                      reg2652 <= ({$unsigned(forvar2594)} - {$unsigned((reg2603 | reg2645))});
                      reg2653 <= reg2604[(1'h1):(1'h1)];
                    end
                  if (((wire2580 ^ (&(reg2608 ? forvar2595 : reg2589))) ?
                      $signed(reg2609) : $unsigned(wire2581[(1'h1):(1'h0)])))
                    begin
                      reg2654 <= (|$unsigned($unsigned(reg2613)));
                      reg2655 <= (reg2627 ?
                          (^~$unsigned((reg2594 ?
                              (8'hb9) : reg2591))) : $signed(((^~reg2616) ?
                              (reg2589 ? reg2615 : (8'hba)) : reg2614)));
                      reg2656 <= ((forvar2595[(1'h1):(1'h1)] ?
                              ((reg2594 ?
                                  wire2582 : reg2617) == wire2580[(2'h3):(1'h0)]) : ((reg2608 * (8'ha2)) != (8'h9f))) ?
                          reg2644 : (reg2629 >>> $unsigned(forvar2600)));
                      reg2657 <= reg2651[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg2654 <= reg2617[(3'h6):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar2648 = (1'h0); (forvar2648 < (1'h0)); forvar2648 = (forvar2648 + (1'h1)))
                    begin
                      reg2649 <= $signed($unsigned($signed((forvar2594 < (8'ha1)))));
                      reg2650 <= reg2636[(3'h5):(3'h4)];
                      reg2651 <= $unsigned(($unsigned(((8'h9d) >>> (8'h9e))) ?
                          (^~reg2598[(4'hd):(4'h9)]) : forvar2609));
                      reg2652 <= forvar2609;
                    end
                  for (forvar2653 = (1'h0); (forvar2653 < (1'h1)); forvar2653 = (forvar2653 + (1'h1)))
                    begin
                      reg2654 <= $unsigned(($signed((reg2597 ?
                              (8'hab) : (8'haf))) ?
                          reg2646[(3'h7):(2'h2)] : ($unsigned(reg2587) | $signed((8'haf)))));
                      reg2655 <= (~^reg2635[(1'h0):(1'h0)]);
                      reg2656 <= $signed((forvar2594 ?
                          forvar2624[(2'h2):(1'h0)] : $signed(reg2625[(3'h6):(3'h5)])));
                      reg2657 <= (^$signed({((8'ha2) + reg2588)}));
                    end
                  reg2658 <= (~|reg2594[(2'h2):(1'h0)]);
                end
              reg2659 <= reg2629[(2'h2):(2'h2)];
              if ($unsigned($unsigned((^~(reg2658 <<< reg2634)))))
                begin
                  reg2660 <= $signed($signed(reg2639));
                  for (forvar2661 = (1'h0); (forvar2661 < (1'h0)); forvar2661 = (forvar2661 + (1'h1)))
                    begin
                      reg2662 <= ($unsigned($unsigned($signed(reg2614))) ?
                          forvar2661 : (|(8'ha4)));
                      reg2663 <= ($unsigned(((reg2652 ? reg2662 : reg2622) ?
                              (8'hb1) : reg2625)) ?
                          ((~|(reg2622 >> forvar2586)) > ((8'had) ?
                              $unsigned(forvar2595) : forvar2594)) : $signed((~$signed((8'h9f)))));
                      reg2664 <= ({reg2655} ?
                          (-({forvar2600} >> reg2657)) : (+forvar2638[(4'hb):(3'h5)]));
                    end
                end
              else
                begin
                  for (forvar2660 = (1'h0); (forvar2660 < (1'h1)); forvar2660 = (forvar2660 + (1'h1)))
                    begin
                      reg2661 <= reg2595[(4'h9):(4'h9)];
                    end
                  reg2662 <= $unsigned(({(reg2628 + reg2646)} ?
                      $signed((reg2623 ?
                          reg2636 : (8'h9c))) : (~reg2642[(2'h2):(1'h0)])));
                end
              for (forvar2665 = (1'h0); (forvar2665 < (2'h3)); forvar2665 = (forvar2665 + (1'h1)))
                begin
                  if (forvar2665)
                    begin
                      reg2666 <= $signed((^{$signed(reg2650)}));
                      reg2667 <= $unsigned($signed($unsigned((forvar2638 >= reg2618))));
                    end
                  else
                    begin
                      reg2666 <= wire2583;
                    end
                end
            end
        end
      else
        begin
          for (forvar2586 = (1'h0); (forvar2586 < (2'h2)); forvar2586 = (forvar2586 + (1'h1)))
            begin
              if ($signed($unsigned($signed({(8'hb3)}))))
                begin
                  if (reg2589[(2'h3):(1'h0)])
                    begin
                      reg2587 <= (wire2581 ?
                          $unsigned(reg2609[(1'h0):(1'h0)]) : ((reg2598 | reg2661) != $signed(((8'hb2) - forvar2638))));
                    end
                  else
                    begin
                      reg2587 <= {forvar2616[(2'h3):(1'h0)]};
                    end
                  for (forvar2588 = (1'h0); (forvar2588 < (2'h2)); forvar2588 = (forvar2588 + (1'h1)))
                    begin
                      reg2589 <= $unsigned($unsigned(forvar2653));
                      reg2590 <= $unsigned((reg2614 ?
                          ((reg2651 - reg2658) < wire2584[(4'h8):(4'h8)]) : {(reg2659 ?
                                  reg2658 : wire2580)}));
                    end
                  for (forvar2591 = (1'h0); (forvar2591 < (2'h2)); forvar2591 = (forvar2591 + (1'h1)))
                    begin
                      reg2592 <= ((~^forvar2615[(3'h4):(3'h4)]) ?
                          $unsigned($signed($signed(reg2597))) : $signed(forvar2647[(3'h5):(1'h0)]));
                      reg2593 <= ((reg2654[(1'h0):(1'h0)] >> (reg2645 < (~forvar2601))) ^ $signed({(~&reg2667)}));
                    end
                end
              else
                begin
                  if ((~$unsigned(reg2622[(2'h2):(2'h2)])))
                    begin
                      reg2587 <= $unsigned(reg2644);
                      reg2588 <= reg2633;
                      reg2589 <= (~^(((&reg2651) ^ reg2587) ?
                          wire2585 : reg2667));
                      reg2590 <= {forvar2588};
                    end
                  else
                    begin
                      reg2587 <= $signed((($unsigned(forvar2650) >>> (|reg2644)) + ({reg2634} ?
                          (reg2586 ? reg2655 : forvar2653) : (forvar2647 ?
                              wire2585 : (8'hb8)))));
                      reg2588 <= ($unsigned((~&(~|(8'haf)))) ^~ forvar2605[(4'ha):(4'ha)]);
                      reg2589 <= reg2648[(4'hc):(1'h0)];
                    end
                  if ({(+(reg2614[(4'h9):(3'h4)] ?
                          {forvar2624} : $unsigned(reg2620)))})
                    begin
                      reg2591 <= reg2588[(1'h1):(1'h1)];
                      reg2592 <= (|((reg2588 ?
                          ((8'ha8) ?
                              forvar2594 : reg2633) : forvar2616[(2'h3):(1'h0)]) == (+(&reg2648))));
                      reg2593 <= {reg2650};
                      reg2594 <= ({$signed(forvar2616)} ?
                          ($signed((reg2595 >> reg2650)) <= reg2649[(1'h0):(1'h0)]) : $signed($signed(((8'had) != reg2617))));
                    end
                  else
                    begin
                      reg2591 <= forvar2602[(1'h0):(1'h0)];
                      reg2592 <= (reg2618 - (((reg2646 & reg2634) < (~&reg2608)) ?
                          (forvar2660 ?
                              $unsigned(reg2617) : (reg2639 < wire2584)) : (~&{reg2617})));
                    end
                  reg2595 <= $unsigned((+(+(forvar2665 != forvar2594))));
                  for (forvar2596 = (1'h0); (forvar2596 < (1'h0)); forvar2596 = (forvar2596 + (1'h1)))
                    begin
                      reg2597 <= (~$signed(($unsigned(reg2645) || (reg2652 ?
                          forvar2586 : (8'ha3)))));
                      reg2598 <= (~|forvar2594);
                    end
                end
            end
        end
    end
  assign wire2668 = reg2588[(3'h7):(2'h2)];
  assign wire2669 = {reg2604};
  assign wire2670 = {reg2595};
  assign wire2671 = $unsigned((reg2623 + $signed(reg2625[(1'h1):(1'h1)])));
  assign wire2672 = reg2612[(4'hb):(4'h9)];
  assign wire2673 = reg2617[(4'hb):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar2674 = (1'h0); (forvar2674 < (2'h3)); forvar2674 = (forvar2674 + (1'h1)))
        begin
          for (forvar2675 = (1'h0); (forvar2675 < (1'h1)); forvar2675 = (forvar2675 + (1'h1)))
            begin
              for (forvar2676 = (1'h0); (forvar2676 < (2'h2)); forvar2676 = (forvar2676 + (1'h1)))
                begin
                  for (forvar2677 = (1'h0); (forvar2677 < (2'h3)); forvar2677 = (forvar2677 + (1'h1)))
                    begin
                      reg2678 <= wire2585;
                    end
                end
              for (forvar2679 = (1'h0); (forvar2679 < (2'h3)); forvar2679 = (forvar2679 + (1'h1)))
                begin
                  for (forvar2680 = (1'h0); (forvar2680 < (2'h2)); forvar2680 = (forvar2680 + (1'h1)))
                    begin
                      reg2681 <= $unsigned((~|{reg2598}));
                      reg2682 <= forvar2679;
                    end
                  reg2683 <= {(((-wire2670) << $signed(reg2596)) ?
                          ($signed(reg2611) ?
                              (-reg2598) : reg2644) : ((8'ha9) ~^ (reg2623 - reg2602)))};
                end
            end
          if (reg2596[(1'h1):(1'h1)])
            begin
              if ((reg2593 ?
                  reg2616[(1'h0):(1'h0)] : (wire2668[(3'h4):(2'h2)] ?
                      reg2662[(1'h1):(1'h1)] : reg2639[(3'h6):(1'h0)])))
                begin
                  for (forvar2684 = (1'h0); (forvar2684 < (2'h2)); forvar2684 = (forvar2684 + (1'h1)))
                    begin
                      reg2685 <= (((wire2673[(4'ha):(4'h9)] ?
                                  (reg2590 >= reg2589) : (reg2615 ?
                                      reg2651 : (8'had))) ?
                              wire2670[(4'h8):(1'h1)] : reg2613) ?
                          {($unsigned(forvar2676) ?
                                  (reg2598 > reg2666) : reg2617)} : reg2598[(1'h1):(1'h1)]);
                      reg2686 <= (($signed($unsigned((8'ha3))) ?
                              wire2672[(2'h2):(1'h0)] : $unsigned((reg2602 | reg2612))) ?
                          ((reg2589[(1'h0):(1'h0)] | (+wire2671)) & $unsigned((reg2625 ?
                              reg2630 : wire2583))) : $signed(((reg2627 ?
                              (8'hb9) : reg2610) >= $signed(reg2594))));
                      reg2687 <= ($unsigned({(!reg2589)}) <<< (-(~|(wire2580 ?
                          reg2593 : forvar2674))));
                    end
                end
              else
                begin
                  for (forvar2684 = (1'h0); (forvar2684 < (1'h0)); forvar2684 = (forvar2684 + (1'h1)))
                    begin
                      reg2685 <= (8'ha0);
                      reg2686 <= reg2652[(3'h6):(3'h5)];
                      reg2687 <= ((reg2663[(2'h3):(1'h1)] ?
                              reg2608[(4'hb):(4'h8)] : (reg2604 ?
                                  $signed((8'had)) : (wire2673 <<< wire2671))) ?
                          (~(~&$signed(reg2622))) : reg2655[(1'h1):(1'h1)]);
                    end
                end
              for (forvar2688 = (1'h0); (forvar2688 < (1'h0)); forvar2688 = (forvar2688 + (1'h1)))
                begin
                  for (forvar2689 = (1'h0); (forvar2689 < (1'h0)); forvar2689 = (forvar2689 + (1'h1)))
                    begin
                      reg2690 <= (reg2640[(3'h7):(3'h5)] | reg2648[(4'ha):(1'h1)]);
                      reg2691 <= $signed(reg2588[(3'h4):(1'h0)]);
                    end
                end
            end
          else
            begin
              reg2684 <= {{{(reg2648 & forvar2680)}}};
              reg2685 <= (((~^(!reg2657)) != ((8'had) ?
                  $unsigned(reg2667) : reg2607)) < $signed($unsigned(reg2691[(3'h5):(1'h0)])));
            end
        end
      if ((($unsigned((reg2648 && reg2662)) ?
              reg2607 : $signed($unsigned((8'hae)))) ?
          {(reg2586 && reg2613)} : $signed(((reg2592 > reg2628) >> reg2635))))
        begin
          for (forvar2692 = (1'h0); (forvar2692 < (2'h3)); forvar2692 = (forvar2692 + (1'h1)))
            begin
              if (wire2585)
                begin
                  reg2693 <= reg2630;
                  for (forvar2694 = (1'h0); (forvar2694 < (1'h0)); forvar2694 = (forvar2694 + (1'h1)))
                    begin
                      reg2695 <= (8'had);
                      reg2696 <= (8'haf);
                      reg2697 <= reg2614;
                    end
                  for (forvar2698 = (1'h0); (forvar2698 < (2'h2)); forvar2698 = (forvar2698 + (1'h1)))
                    begin
                      reg2699 <= $signed($unsigned(reg2613));
                    end
                end
              else
                begin
                  reg2693 <= reg2614;
                end
              for (forvar2700 = (1'h0); (forvar2700 < (1'h1)); forvar2700 = (forvar2700 + (1'h1)))
                begin
                  for (forvar2701 = (1'h0); (forvar2701 < (2'h2)); forvar2701 = (forvar2701 + (1'h1)))
                    begin
                      reg2702 <= $unsigned(reg2654);
                      reg2703 <= reg2609;
                    end
                end
            end
          for (forvar2704 = (1'h0); (forvar2704 < (1'h0)); forvar2704 = (forvar2704 + (1'h1)))
            begin
              reg2705 <= {{{(reg2642 ? reg2682 : wire2672)}}};
            end
          if (($unsigned(($signed(wire2673) ? $signed(forvar2700) : (8'hb9))) ?
              (reg2639 ?
                  $unsigned($signed(reg2703)) : $unsigned((reg2590 ?
                      reg2696 : reg2599))) : $signed(wire2671[(1'h0):(1'h0)])))
            begin
              for (forvar2706 = (1'h0); (forvar2706 < (1'h0)); forvar2706 = (forvar2706 + (1'h1)))
                begin
                  for (forvar2707 = (1'h0); (forvar2707 < (1'h1)); forvar2707 = (forvar2707 + (1'h1)))
                    begin
                      reg2708 <= (({(reg2634 - reg2655)} ?
                          (8'h9f) : {$signed((8'hac))}) != ((+forvar2706[(1'h1):(1'h0)]) != ($unsigned(wire2672) != (!reg2588))));
                      reg2709 <= (^~((+reg2617) ?
                          reg2684 : $unsigned($unsigned(reg2662))));
                      reg2710 <= $unsigned({(((8'ha7) ? (8'h9c) : reg2702) ?
                              reg2616[(4'h8):(3'h6)] : (reg2627 ?
                                  wire2671 : reg2687))});
                      reg2711 <= {reg2683[(1'h0):(1'h0)]};
                    end
                end
              if ((~(!(reg2667 ? reg2640 : $signed(reg2610)))))
                begin
                  for (forvar2712 = (1'h0); (forvar2712 < (1'h1)); forvar2712 = (forvar2712 + (1'h1)))
                    begin
                      reg2713 <= reg2621[(3'h7):(1'h1)];
                    end
                  if (($unsigned($signed(reg2713[(3'h5):(1'h1)])) >>> (($signed((8'hba)) ?
                      $signed(reg2699) : (+(8'hb1))) <= (^~(reg2597 ?
                      reg2635 : reg2616)))))
                    begin
                      reg2714 <= (forvar2700[(2'h3):(2'h2)] ?
                          $unsigned($unsigned({reg2598})) : $signed((((8'ha4) & (8'ha5)) & reg2633[(3'h4):(2'h2)])));
                      reg2715 <= (^(~^(~^forvar2689)));
                      reg2716 <= (wire2582[(2'h2):(2'h2)] ?
                          ((reg2655[(3'h4):(1'h0)] ?
                              {reg2590} : $unsigned((8'haf))) > ({forvar2698} ?
                              ((8'ha1) ?
                                  reg2592 : (8'haa)) : wire2580)) : reg2666);
                      reg2717 <= (8'ha6);
                    end
                  else
                    begin
                      reg2714 <= {$signed(((forvar2712 ? reg2656 : reg2699) ?
                              (reg2633 * wire2583) : reg2667))};
                      reg2715 <= {$unsigned(reg2713[(3'h5):(1'h1)])};
                      reg2716 <= ((8'hae) ?
                          (((^~reg2606) ? (reg2703 < (8'ha1)) : (&reg2593)) ?
                              ((~reg2658) < (^~reg2687)) : $unsigned((reg2654 ?
                                  reg2629 : reg2682))) : $unsigned($unsigned({reg2702})));
                      reg2717 <= reg2708[(3'h5):(1'h0)];
                    end
                  for (forvar2718 = (1'h0); (forvar2718 < (2'h3)); forvar2718 = (forvar2718 + (1'h1)))
                    begin
                      reg2719 <= (((~^(reg2655 + reg2661)) < $signed(reg2604)) + reg2703);
                    end
                  if (reg2703[(3'h4):(1'h0)])
                    begin
                      reg2720 <= $unsigned((!((~|(8'h9f)) >>> $unsigned(reg2589))));
                    end
                  else
                    begin
                      reg2720 <= $signed((((~|reg2629) ?
                              (reg2666 ? reg2603 : forvar2684) : (reg2708 ?
                                  (8'ha2) : reg2635)) ?
                          $signed(reg2589[(2'h2):(1'h1)]) : (|$signed(reg2717))));
                      reg2721 <= ((&forvar2684) <= $unsigned($unsigned({reg2659})));
                      reg2722 <= ({$signed({reg2683})} ?
                          reg2623 : (((~wire2670) ?
                              (~(8'hb8)) : (reg2586 ^ reg2610)) <<< {reg2627[(1'h0):(1'h0)]}));
                      reg2723 <= ($signed((reg2654 ^ (reg2617 ?
                          reg2696 : forvar2692))) > $unsigned(reg2684[(2'h2):(2'h2)]));
                    end
                end
              else
                begin
                  reg2712 <= (+$unsigned({reg2609[(4'he):(3'h4)]}));
                  if ((((|$unsigned(reg2696)) ?
                          (|(reg2720 <<< (8'h9c))) : (reg2608 | (8'ha7))) ?
                      reg2610 : (|((reg2598 ~^ forvar2674) ?
                          (reg2682 >> forvar2704) : (wire2584 >>> forvar2689)))))
                    begin
                      reg2713 <= $unsigned((($signed(reg2613) + reg2634[(3'h4):(3'h4)]) + ($unsigned((8'hac)) ?
                          $signed(reg2604) : (forvar2689 ?
                              (8'hb3) : (8'hb3)))));
                      reg2714 <= $unsigned((^~reg2592));
                    end
                  else
                    begin
                      reg2713 <= $signed((^$unsigned($unsigned((8'h9e)))));
                    end
                  reg2715 <= (wire2582[(2'h3):(1'h0)] * $signed((8'had)));
                end
            end
          else
            begin
              reg2706 <= {$signed(reg2720[(1'h0):(1'h0)])};
              for (forvar2707 = (1'h0); (forvar2707 < (1'h0)); forvar2707 = (forvar2707 + (1'h1)))
                begin
                  if ($unsigned(($unsigned((&wire2669)) ?
                      ({reg2599} ^ reg2633) : forvar2700[(3'h4):(2'h2)])))
                    begin
                      reg2708 <= reg2663[(3'h4):(3'h4)];
                      reg2709 <= (8'haf);
                      reg2710 <= (8'hb1);
                    end
                  else
                    begin
                      reg2708 <= (!(!{(reg2713 != (8'hb4))}));
                      reg2709 <= forvar2679;
                      reg2710 <= (~&(^~wire2582));
                    end
                  for (forvar2711 = (1'h0); (forvar2711 < (1'h1)); forvar2711 = (forvar2711 + (1'h1)))
                    begin
                      reg2712 <= ((reg2715[(3'h4):(3'h4)] ~^ reg2661) <<< $signed((-wire2671)));
                      reg2713 <= $signed($signed(reg2684[(3'h7):(2'h2)]));
                      reg2714 <= wire2671;
                      reg2715 <= {(~$signed($signed(reg2627)))};
                    end
                  for (forvar2716 = (1'h0); (forvar2716 < (1'h0)); forvar2716 = (forvar2716 + (1'h1)))
                    begin
                      reg2717 <= ((8'hb2) ? (8'ha4) : reg2649[(2'h2):(1'h0)]);
                      reg2718 <= reg2660[(2'h2):(1'h1)];
                    end
                end
              if (($signed(forvar2677) + (((reg2594 ?
                      reg2652 : (8'ha5)) ^~ reg2609) ?
                  {reg2636} : $unsigned({(8'hae)}))))
                begin
                  for (forvar2719 = (1'h0); (forvar2719 < (2'h3)); forvar2719 = (forvar2719 + (1'h1)))
                    begin
                      reg2720 <= ((^~(~|(^~forvar2716))) ^~ reg2664[(3'h6):(3'h5)]);
                      reg2721 <= reg2682[(4'hc):(4'h9)];
                      reg2722 <= ((reg2714 + forvar2680[(4'h9):(3'h6)]) ?
                          (($unsigned(reg2607) <<< (~|reg2618)) ?
                              $unsigned((reg2621 ?
                                  reg2699 : reg2640)) : ($signed(reg2615) ?
                                  reg2713 : $unsigned(reg2645))) : ($signed(reg2587) << ((reg2695 ?
                                  forvar2680 : reg2605) ?
                              $unsigned(forvar2680) : (reg2605 ?
                                  reg2586 : reg2599))));
                    end
                  reg2723 <= $unsigned(forvar2688[(4'hb):(2'h3)]);
                  if ($unsigned((~&($signed(reg2709) ?
                      $signed(reg2642) : wire2581))))
                    begin
                      reg2724 <= (reg2690[(1'h1):(1'h1)] >>> $signed(wire2670[(3'h4):(2'h2)]));
                      reg2725 <= wire2671;
                      reg2726 <= reg2682[(4'ha):(4'h9)];
                    end
                  else
                    begin
                      reg2724 <= (+($signed((reg2725 ? reg2648 : reg2721)) ?
                          $unsigned(reg2655) : $signed({reg2702})));
                    end
                end
              else
                begin
                  reg2719 <= (reg2606[(3'h4):(1'h1)] ?
                      reg2606[(1'h0):(1'h0)] : ((|(reg2710 ?
                          wire2585 : forvar2688)) && $unsigned((reg2598 >>> reg2586))));
                  if (({{{reg2605}}} ?
                      {((+wire2583) ?
                              wire2584 : $unsigned(reg2649))} : forvar2688[(3'h5):(3'h5)]))
                    begin
                      reg2720 <= $signed((~&(8'ha9)));
                      reg2721 <= $unsigned($signed((&reg2725[(3'h4):(1'h1)])));
                      reg2722 <= (^~reg2686);
                      reg2723 <= forvar2701;
                    end
                  else
                    begin
                      reg2720 <= reg2619;
                      reg2721 <= $signed(reg2617);
                    end
                  reg2724 <= reg2655[(1'h1):(1'h0)];
                end
              reg2727 <= $signed(($unsigned($signed(wire2584)) ~^ ($signed(reg2641) ?
                  (-forvar2704) : reg2641)));
            end
          reg2728 <= $signed(forvar2675[(4'hf):(1'h1)]);
        end
      else
        begin
          reg2692 <= (&$unsigned(reg2623));
          if ((reg2617[(2'h3):(2'h2)] ?
              ({(~|reg2606)} + $unsigned(reg2718[(4'h9):(3'h4)])) : reg2609))
            begin
              for (forvar2693 = (1'h0); (forvar2693 < (1'h1)); forvar2693 = (forvar2693 + (1'h1)))
                begin
                  if ({(((reg2592 ?
                              forvar2700 : reg2636) == $unsigned(wire2580)) ?
                          $signed((reg2605 ?
                              reg2603 : reg2659)) : wire2582[(1'h0):(1'h0)])})
                    begin
                      reg2694 <= {$signed(wire2585[(2'h2):(2'h2)])};
                      reg2695 <= $signed(reg2708);
                      reg2696 <= (reg2653[(2'h2):(2'h2)] << reg2711[(3'h6):(3'h5)]);
                    end
                  else
                    begin
                      reg2694 <= $unsigned($signed(($signed(reg2657) == reg2657[(4'h9):(1'h0)])));
                      reg2695 <= $signed($signed(reg2630));
                      reg2696 <= $signed(reg2617[(2'h3):(1'h1)]);
                    end
                  for (forvar2697 = (1'h0); (forvar2697 < (1'h1)); forvar2697 = (forvar2697 + (1'h1)))
                    begin
                      reg2698 <= $unsigned(reg2726);
                      reg2699 <= reg2612[(2'h3):(1'h1)];
                    end
                  for (forvar2700 = (1'h0); (forvar2700 < (1'h0)); forvar2700 = (forvar2700 + (1'h1)))
                    begin
                      reg2701 <= (~&(~^(((8'hac) ? reg2651 : forvar2719) ?
                          (^~(8'ha4)) : {reg2709})));
                    end
                end
              for (forvar2702 = (1'h0); (forvar2702 < (2'h3)); forvar2702 = (forvar2702 + (1'h1)))
                begin
                  for (forvar2703 = (1'h0); (forvar2703 < (2'h3)); forvar2703 = (forvar2703 + (1'h1)))
                    begin
                      reg2704 <= ($unsigned(($signed(forvar2677) ?
                              reg2678 : $signed((8'ha9)))) ?
                          reg2695 : $unsigned((~|reg2712)));
                    end
                  if (($signed({(^~reg2694)}) ?
                      ((^~$unsigned(reg2725)) != $unsigned($unsigned(reg2625))) : forvar2692))
                    begin
                      reg2705 <= (-$signed(reg2593[(3'h6):(3'h5)]));
                      reg2706 <= $unsigned(reg2692);
                      reg2707 <= ((8'h9c) ^~ (wire2581[(2'h2):(2'h2)] <<< ($unsigned(reg2725) ?
                          reg2628[(2'h2):(1'h1)] : wire2581)));
                    end
                  else
                    begin
                      reg2705 <= (reg2713 + $unsigned(((8'haf) > (-reg2697))));
                      reg2706 <= $signed((^~(~^(^~reg2639))));
                      reg2707 <= reg2727;
                      reg2708 <= $unsigned(reg2716[(4'ha):(2'h2)]);
                    end
                  reg2709 <= (-forvar2698[(2'h2):(2'h2)]);
                end
              for (forvar2710 = (1'h0); (forvar2710 < (1'h0)); forvar2710 = (forvar2710 + (1'h1)))
                begin
                  for (forvar2711 = (1'h0); (forvar2711 < (2'h2)); forvar2711 = (forvar2711 + (1'h1)))
                    begin
                      reg2712 <= (^~reg2648[(4'hd):(2'h3)]);
                      reg2713 <= reg2644;
                    end
                end
              for (forvar2714 = (1'h0); (forvar2714 < (2'h2)); forvar2714 = (forvar2714 + (1'h1)))
                begin
                  if ({(^$unsigned(forvar2689))})
                    begin
                      reg2715 <= (~|((forvar2710 * (reg2721 ?
                          reg2706 : wire2581)) <= (8'h9f)));
                      reg2716 <= reg2649[(2'h3):(2'h3)];
                      reg2717 <= (&$unsigned({$unsigned((8'hac))}));
                      reg2718 <= $unsigned(reg2590);
                    end
                  else
                    begin
                      reg2715 <= forvar2674;
                      reg2716 <= (reg2609 ?
                          {reg2631[(1'h0):(1'h0)]} : (forvar2688[(4'hc):(3'h5)] ?
                              reg2660 : $signed($unsigned(reg2596))));
                      reg2717 <= reg2684;
                    end
                  if ((forvar2692[(1'h1):(1'h1)] ?
                      reg2693 : $unsigned(reg2618[(3'h4):(1'h0)])))
                    begin
                      reg2719 <= $signed(reg2642[(2'h3):(1'h0)]);
                      reg2720 <= ($signed({((8'hb7) <<< reg2640)}) <= {reg2610});
                      reg2721 <= ($unsigned(reg2598[(4'he):(3'h6)]) ?
                          $signed(forvar2702) : forvar2704[(3'h6):(1'h0)]);
                    end
                  else
                    begin
                      reg2719 <= $signed((^({reg2663} > (~&(8'ha4)))));
                      reg2720 <= (-(!($unsigned((8'haf)) ?
                          reg2625 : (forvar2719 || reg2710))));
                      reg2721 <= ({forvar2684} && ($unsigned((~&reg2655)) < reg2723));
                      reg2722 <= (~^(((reg2645 < (8'ha0)) ?
                              (^~reg2612) : $unsigned(reg2608)) ?
                          reg2604[(4'hd):(3'h5)] : $unsigned((forvar2703 ?
                              (8'hae) : reg2693))));
                    end
                end
            end
          else
            begin
              if (reg2667[(3'h4):(2'h2)])
                begin
                  reg2693 <= $signed($unsigned($unsigned({(8'ha6)})));
                  if ($signed((~&reg2704)))
                    begin
                      reg2694 <= reg2653;
                      reg2695 <= reg2685[(4'h9):(2'h2)];
                    end
                  else
                    begin
                      reg2694 <= {reg2629[(1'h0):(1'h0)]};
                      reg2695 <= {reg2644[(2'h2):(1'h1)]};
                    end
                  for (forvar2696 = (1'h0); (forvar2696 < (2'h2)); forvar2696 = (forvar2696 + (1'h1)))
                    begin
                      reg2697 <= reg2604[(4'hd):(3'h7)];
                      reg2698 <= (+reg2709[(3'h5):(1'h1)]);
                      reg2699 <= (reg2718 ?
                          ($signed({reg2620}) <= (&(reg2650 && (8'hab)))) : reg2695[(3'h4):(1'h1)]);
                      reg2700 <= {($unsigned(reg2724[(4'h8):(3'h5)]) >>> (8'hb3))};
                    end
                  if (reg2636)
                    begin
                      reg2701 <= (reg2681 || {(8'h9e)});
                      reg2702 <= (&reg2710[(4'h8):(3'h4)]);
                    end
                  else
                    begin
                      reg2701 <= reg2662[(1'h0):(1'h0)];
                      reg2702 <= forvar2694[(4'h8):(3'h6)];
                      reg2703 <= $signed(((~&(forvar2696 | forvar2711)) == (8'hb4)));
                      reg2704 <= (wire2673[(4'hd):(4'hd)] - forvar2703);
                    end
                end
              else
                begin
                  for (forvar2693 = (1'h0); (forvar2693 < (1'h0)); forvar2693 = (forvar2693 + (1'h1)))
                    begin
                      reg2694 <= reg2703[(3'h7):(3'h5)];
                    end
                end
              for (forvar2705 = (1'h0); (forvar2705 < (1'h0)); forvar2705 = (forvar2705 + (1'h1)))
                begin
                  if (forvar2716)
                    begin
                      reg2706 <= (|$unsigned(reg2633[(2'h2):(2'h2)]));
                      reg2707 <= ((forvar2714 ^ reg2720[(2'h2):(1'h1)]) ?
                          {wire2580[(4'h9):(4'h9)]} : $unsigned((~reg2712[(2'h2):(1'h1)])));
                      reg2708 <= (~^$signed((reg2696 ?
                          ((8'ha2) ^~ forvar2706) : $unsigned((8'hb8)))));
                    end
                  else
                    begin
                      reg2706 <= (forvar2719 ?
                          ($unsigned((reg2704 >= reg2667)) << (reg2726 < $unsigned(forvar2676))) : (^($unsigned(reg2662) <= reg2654)));
                      reg2707 <= ((~|(reg2588[(3'h4):(1'h1)] ?
                              (^~wire2581) : $unsigned(reg2723))) ?
                          (forvar2698[(1'h0):(1'h0)] & (reg2606[(3'h7):(3'h6)] <<< (forvar2674 ?
                              reg2631 : wire2669))) : (~^reg2710[(3'h4):(1'h1)]));
                      reg2708 <= $signed($unsigned($signed($unsigned(reg2627))));
                    end
                  for (forvar2709 = (1'h0); (forvar2709 < (1'h0)); forvar2709 = (forvar2709 + (1'h1)))
                    begin
                      reg2710 <= (((forvar2716[(2'h3):(1'h0)] ?
                                  {reg2607} : (reg2723 ?
                                      forvar2712 : (8'hb3))) ?
                              {(-(8'hb1))} : {forvar2701}) ?
                          (reg2604[(3'h5):(1'h0)] ?
                              $unsigned((+reg2704)) : (forvar2716 ?
                                  (|reg2636) : forvar2719)) : ((8'hb8) ?
                              reg2718[(1'h0):(1'h0)] : ((wire2670 ?
                                      reg2726 : forvar2710) ?
                                  (+reg2654) : (8'h9c))));
                      reg2711 <= ((($unsigned((8'ha9)) ?
                          reg2704[(1'h0):(1'h0)] : (|reg2664)) && $unsigned(reg2702)) | (((reg2618 || reg2616) < $unsigned((8'h9c))) ?
                          {(^reg2707)} : {reg2712}));
                      reg2712 <= reg2717;
                      reg2713 <= ($signed((~|(8'hba))) ?
                          (+$signed((-reg2607))) : (reg2636 ~^ ($signed(reg2613) ?
                              forvar2707 : (reg2650 <<< (8'hb8)))));
                    end
                  for (forvar2714 = (1'h0); (forvar2714 < (1'h1)); forvar2714 = (forvar2714 + (1'h1)))
                    begin
                      reg2715 <= (^~(!$signed($unsigned(forvar2694))));
                    end
                  if ((8'hb8))
                    begin
                      reg2716 <= {(|((forvar2704 & reg2614) ?
                              (|reg2707) : (~&(8'ha2))))};
                      reg2717 <= (^~reg2633);
                      reg2718 <= (~reg2697);
                      reg2719 <= ($signed((reg2593 ?
                              wire2668 : $signed((8'hb6)))) ?
                          (~&$signed(((8'ha8) ?
                              reg2699 : reg2685))) : $unsigned($unsigned((reg2610 ?
                              forvar2712 : reg2642))));
                    end
                  else
                    begin
                      reg2716 <= $unsigned(reg2695);
                      reg2717 <= (~$unsigned(((reg2714 ?
                          reg2613 : wire2582) & ((8'ha0) || reg2724))));
                      reg2718 <= wire2584;
                    end
                end
              if ((reg2708 <<< (!(((8'hb6) & (8'ha0)) ?
                  (reg2692 + reg2684) : (reg2641 && forvar2697)))))
                begin
                  reg2720 <= {(({reg2653} ?
                              $signed(reg2617) : forvar2693[(1'h0):(1'h0)]) ?
                          ($unsigned(reg2683) ^~ (reg2631 ?
                              reg2657 : reg2625)) : $signed(reg2697))};
                end
              else
                begin
                  for (forvar2720 = (1'h0); (forvar2720 < (2'h3)); forvar2720 = (forvar2720 + (1'h1)))
                    begin
                      reg2721 <= $unsigned({(|(~|reg2704))});
                    end
                  for (forvar2722 = (1'h0); (forvar2722 < (2'h3)); forvar2722 = (forvar2722 + (1'h1)))
                    begin
                      reg2723 <= (((forvar2706[(1'h1):(1'h0)] ?
                          $signed(reg2698) : $unsigned(reg2646)) ^~ reg2698[(4'h9):(3'h6)]) > reg2654[(1'h0):(1'h0)]);
                      reg2724 <= (reg2650[(4'h9):(4'h8)] ?
                          $unsigned((forvar2700 ?
                              $unsigned((8'hb6)) : wire2668[(3'h7):(3'h5)])) : (reg2588 - (+(wire2668 >> reg2699))));
                    end
                end
            end
          for (forvar2725 = (1'h0); (forvar2725 < (1'h1)); forvar2725 = (forvar2725 + (1'h1)))
            begin
              for (forvar2726 = (1'h0); (forvar2726 < (1'h0)); forvar2726 = (forvar2726 + (1'h1)))
                begin
                  for (forvar2727 = (1'h0); (forvar2727 < (2'h3)); forvar2727 = (forvar2727 + (1'h1)))
                    begin
                      reg2728 <= ({reg2720} >> $signed(reg2589[(3'h4):(2'h3)]));
                      reg2729 <= $unsigned(((reg2604 >= (|(8'ha7))) ?
                          ($signed((8'hb3)) != reg2609[(4'h8):(2'h3)]) : (reg2684 ?
                              $unsigned(reg2639) : (8'ha8))));
                      reg2730 <= ($signed(((reg2620 == reg2619) ?
                          reg2591[(4'h8):(3'h7)] : forvar2700)) && $signed($signed($signed(reg2607))));
                      reg2731 <= reg2620[(4'h9):(4'h9)];
                    end
                  for (forvar2732 = (1'h0); (forvar2732 < (1'h1)); forvar2732 = (forvar2732 + (1'h1)))
                    begin
                      reg2733 <= ($unsigned((~&(forvar2703 ~^ reg2594))) ?
                          ($signed((&reg2586)) >= (((8'hac) ?
                              forvar2714 : reg2654) == $signed(reg2725))) : (!$unsigned($unsigned(reg2617))));
                      reg2734 <= ((-(~&$unsigned(reg2627))) ?
                          $signed(reg2700) : ((+wire2583) * reg2596));
                      reg2735 <= reg2721[(1'h1):(1'h1)];
                    end
                end
              if (wire2583[(2'h2):(1'h0)])
                begin
                  if (reg2666)
                    begin
                      reg2736 <= (~&((|reg2614) <= $unsigned(forvar2689)));
                      reg2737 <= ((^~((reg2727 ?
                              forvar2705 : (8'ha6)) >>> $unsigned(forvar2725))) ?
                          reg2691 : (forvar2700[(1'h0):(1'h0)] ?
                              (~$signed(reg2623)) : ($signed(forvar2709) * reg2634)));
                    end
                  else
                    begin
                      reg2736 <= ((~^($signed(reg2685) ?
                              (^~reg2687) : reg2707[(3'h6):(1'h1)])) ?
                          (|(~^{(8'had)})) : (^~forvar2710[(3'h7):(1'h0)]));
                      reg2737 <= ((reg2594[(2'h3):(1'h1)] ?
                          reg2597[(3'h6):(3'h4)] : $unsigned(reg2661[(1'h1):(1'h1)])) ^ $unsigned($signed(((8'hb5) >> reg2727))));
                      reg2738 <= (forvar2693 ?
                          reg2592[(4'he):(3'h5)] : {reg2598});
                    end
                  if (reg2724)
                    begin
                      reg2739 <= {(+reg2709[(3'h4):(1'h1)])};
                      reg2740 <= $unsigned({(8'ha5)});
                    end
                  else
                    begin
                      reg2739 <= reg2710[(3'h6):(1'h0)];
                      reg2740 <= reg2723;
                      reg2741 <= reg2603;
                      reg2742 <= {$signed((~wire2582[(3'h7):(1'h1)]))};
                    end
                  for (forvar2743 = (1'h0); (forvar2743 < (2'h2)); forvar2743 = (forvar2743 + (1'h1)))
                    begin
                      reg2744 <= (~&(&reg2655));
                      reg2745 <= forvar2707[(4'h8):(1'h0)];
                      reg2746 <= wire2580[(4'he):(3'h7)];
                    end
                end
              else
                begin
                  if (((reg2597 ?
                      (~(forvar2727 ?
                          forvar2727 : reg2656)) : $signed($signed(reg2659))) | (reg2654[(2'h3):(1'h0)] ?
                      $signed(reg2717) : (~(reg2727 | reg2596)))))
                    begin
                      reg2736 <= reg2635;
                      reg2737 <= reg2723;
                      reg2738 <= (-reg2657[(4'hc):(2'h2)]);
                    end
                  else
                    begin
                      reg2736 <= ({forvar2719} >>> (8'hb7));
                      reg2737 <= $signed((reg2662 ?
                          reg2716[(4'h8):(2'h2)] : reg2631));
                      reg2738 <= (|reg2666[(2'h2):(1'h1)]);
                      reg2739 <= $unsigned(reg2592);
                    end
                  for (forvar2740 = (1'h0); (forvar2740 < (1'h1)); forvar2740 = (forvar2740 + (1'h1)))
                    begin
                      reg2741 <= ((~&$signed({reg2698})) + (&$signed(forvar2719)));
                    end
                  if ((~|reg2641[(1'h1):(1'h1)]))
                    begin
                      reg2742 <= ($unsigned((|{reg2588})) ^ ({reg2712[(3'h4):(2'h3)]} ?
                          $signed((|forvar2732)) : (~&$signed(reg2712))));
                      reg2743 <= reg2650[(4'ha):(1'h1)];
                      reg2744 <= $unsigned({$signed({reg2743})});
                      reg2745 <= (reg2737 != reg2617);
                    end
                  else
                    begin
                      reg2742 <= $signed($unsigned(forvar2688[(4'hb):(4'ha)]));
                    end
                  if ({$signed(reg2617[(4'h9):(3'h7)])})
                    begin
                      reg2746 <= (~^reg2712);
                      reg2747 <= reg2725[(1'h0):(1'h0)];
                      reg2748 <= reg2663;
                    end
                  else
                    begin
                      reg2746 <= ($signed((~$signed(reg2683))) ?
                          (^{$unsigned((8'hb2))}) : (forvar2725 ?
                              reg2602[(4'hc):(1'h1)] : reg2687));
                      reg2747 <= {$unsigned($unsigned(reg2652[(1'h1):(1'h0)]))};
                      reg2748 <= reg2719[(1'h1):(1'h1)];
                      reg2749 <= (!$unsigned(reg2587));
                    end
                end
            end
          if (forvar2693[(3'h5):(1'h0)])
            begin
              for (forvar2750 = (1'h0); (forvar2750 < (1'h1)); forvar2750 = (forvar2750 + (1'h1)))
                begin
                  for (forvar2751 = (1'h0); (forvar2751 < (1'h1)); forvar2751 = (forvar2751 + (1'h1)))
                    begin
                      reg2752 <= (wire2581 ?
                          (((^reg2652) <= (~|reg2602)) << reg2608[(2'h2):(1'h0)]) : (8'hab));
                    end
                  if ({reg2728})
                    begin
                      reg2753 <= $signed((^$unsigned((~reg2653))));
                    end
                  else
                    begin
                      reg2753 <= wire2669;
                      reg2754 <= $unsigned((+forvar2732));
                      reg2755 <= ((8'hb4) ?
                          (((~&forvar2703) ? reg2692 : (8'hba)) ?
                              forvar2692 : (~&(wire2580 ?
                                  reg2609 : reg2753))) : ((+(reg2600 ?
                                  (8'hb2) : wire2582)) ?
                              (forvar2709[(5'h10):(1'h1)] ^~ (reg2696 ?
                                  wire2580 : (8'h9d))) : $unsigned(forvar2712[(4'hb):(4'h8)])));
                    end
                  if ($unsigned((|((reg2702 ? forvar2674 : reg2633) ?
                      reg2691[(4'hc):(4'h8)] : ((8'hb8) ? (8'h9d) : reg2603)))))
                    begin
                      reg2756 <= $unsigned($unsigned(forvar2720[(2'h3):(2'h3)]));
                      reg2757 <= reg2708;
                      reg2758 <= forvar2719[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg2756 <= $signed({reg2657});
                      reg2757 <= ({$signed((reg2704 ?
                              reg2610 : reg2724))} ^~ (forvar2707 ?
                          ((|reg2736) ?
                              $unsigned(reg2687) : {reg2639}) : $unsigned((8'hb6))));
                      reg2758 <= $signed((&(8'ha8)));
                    end
                end
              if ($unsigned((8'hb9)))
                begin
                  for (forvar2759 = (1'h0); (forvar2759 < (2'h2)); forvar2759 = (forvar2759 + (1'h1)))
                    begin
                      reg2760 <= $signed((((forvar2679 ?
                                  forvar2707 : forvar2743) ?
                              (reg2657 ? wire2581 : reg2712) : forvar2698) ?
                          $signed(forvar2676) : reg2757[(1'h1):(1'h0)]));
                    end
                  for (forvar2761 = (1'h0); (forvar2761 < (1'h1)); forvar2761 = (forvar2761 + (1'h1)))
                    begin
                      reg2762 <= ((~&($unsigned(reg2640) ?
                          (^~reg2619) : reg2616[(1'h1):(1'h1)])) < (!$signed({reg2749})));
                    end
                end
              else
                begin
                  reg2759 <= $unsigned(((~|(forvar2677 ?
                      forvar2707 : reg2610)) ^ $signed($signed((8'ha2)))));
                  if ((~|$signed($signed((reg2596 ? reg2633 : reg2654)))))
                    begin
                      reg2760 <= (($unsigned(reg2736[(2'h3):(2'h3)]) ?
                              ((forvar2676 && (8'ha9)) != reg2724[(3'h5):(3'h4)]) : (&$signed(reg2631))) ?
                          reg2682[(1'h1):(1'h0)] : (reg2695 ~^ $signed((forvar2696 ~^ (8'haf)))));
                      reg2761 <= (~^(-$unsigned({reg2610})));
                      reg2762 <= {reg2620[(2'h3):(2'h3)]};
                    end
                  else
                    begin
                      reg2760 <= ((forvar2725 ?
                          (&(reg2684 ? reg2599 : forvar2751)) : ((reg2698 ?
                              reg2705 : reg2660) - $unsigned(reg2614))) << {((forvar2707 ?
                                  (8'ha0) : reg2633) ?
                              $unsigned(reg2701) : (reg2599 >>> reg2705))});
                      reg2761 <= forvar2680;
                      reg2762 <= $unsigned($signed((reg2652[(1'h0):(1'h0)] ?
                          $signed(reg2630) : reg2723)));
                      reg2763 <= $signed({$signed($unsigned(reg2640))});
                    end
                end
            end
          else
            begin
              if ($unsigned((&reg2729[(3'h7):(2'h2)])))
                begin
                  if (($unsigned($unsigned(reg2627[(3'h4):(2'h3)])) << $unsigned($signed($signed(forvar2676)))))
                    begin
                      reg2750 <= $unsigned((wire2582 ^~ forvar2705));
                      reg2751 <= {$unsigned($signed({reg2693}))};
                      reg2752 <= reg2655;
                    end
                  else
                    begin
                      reg2750 <= $signed(reg2714[(3'h4):(1'h1)]);
                      reg2751 <= ($signed(((reg2613 ? reg2603 : (8'hb6)) ?
                          (&reg2694) : $unsigned(reg2755))) ^ $signed($signed((!reg2697))));
                    end
                  for (forvar2753 = (1'h0); (forvar2753 < (2'h3)); forvar2753 = (forvar2753 + (1'h1)))
                    begin
                      reg2754 <= reg2587[(1'h0):(1'h0)];
                      reg2755 <= ((~&(reg2597[(3'h6):(3'h6)] ?
                              reg2635 : (forvar2693 ~^ forvar2677))) ?
                          ((~|(!(8'hb1))) <= reg2617[(3'h6):(3'h5)]) : forvar2720);
                      reg2756 <= ((^~reg2639) ?
                          ($signed((reg2746 ?
                              wire2584 : (8'ha7))) * (8'hb7)) : (|$signed($unsigned((8'ha6)))));
                    end
                end
              else
                begin
                  if (reg2726[(4'ha):(4'h8)])
                    begin
                      reg2750 <= $unsigned($unsigned($signed((~(8'ha0)))));
                      reg2751 <= $unsigned(($signed($unsigned(reg2644)) ?
                          {(&reg2658)} : (reg2623 ?
                              $unsigned((8'hb3)) : {(8'h9d)})));
                    end
                  else
                    begin
                      reg2750 <= (($signed(((8'ha5) ?
                          (8'hb3) : (8'hb7))) | (8'h9f)) >> wire2670);
                      reg2751 <= $signed((^$signed((!reg2610))));
                      reg2752 <= $unsigned((|$unsigned(reg2632)));
                      reg2753 <= (-(((~reg2761) >= (forvar2675 == reg2592)) ?
                          reg2742[(3'h7):(3'h6)] : $unsigned((reg2725 + reg2707))));
                    end
                  for (forvar2754 = (1'h0); (forvar2754 < (1'h1)); forvar2754 = (forvar2754 + (1'h1)))
                    begin
                      reg2755 <= reg2739;
                      reg2756 <= $signed((reg2632[(2'h3):(1'h0)] <<< reg2710));
                      reg2757 <= {$unsigned((~&forvar2693[(4'hb):(4'h8)]))};
                    end
                  if (((reg2639 - reg2600) ?
                      {$unsigned($signed(reg2720))} : $unsigned(((reg2653 ?
                              reg2742 : (8'ha4)) ?
                          $unsigned(reg2690) : {reg2709}))))
                    begin
                      reg2758 <= (!(8'hac));
                    end
                  else
                    begin
                      reg2758 <= (+wire2580[(4'h8):(2'h3)]);
                      reg2759 <= ($signed(reg2627) >> {{$unsigned((8'h9c))}});
                    end
                end
              for (forvar2760 = (1'h0); (forvar2760 < (2'h3)); forvar2760 = (forvar2760 + (1'h1)))
                begin
                  if (({$unsigned((reg2630 ? (8'haa) : reg2761))} == reg2634))
                    begin
                      reg2761 <= reg2738;
                      reg2762 <= ($unsigned($unsigned((reg2739 || forvar2714))) ?
                          (8'hb0) : (reg2714[(4'h8):(2'h2)] & (|$signed(reg2661))));
                      reg2763 <= reg2752;
                    end
                  else
                    begin
                      reg2761 <= reg2594;
                      reg2762 <= (reg2693[(4'ha):(1'h0)] ?
                          (^~$signed((reg2629 ?
                              (8'hb4) : forvar2698))) : (reg2608 ?
                              reg2751[(4'h8):(1'h1)] : forvar2720[(4'h9):(3'h5)]));
                    end
                  for (forvar2764 = (1'h0); (forvar2764 < (2'h2)); forvar2764 = (forvar2764 + (1'h1)))
                    begin
                      reg2765 <= (($signed((reg2636 ? (8'hb1) : reg2630)) ?
                          (^~$signed((8'h9e))) : (8'haa)) >= $unsigned(reg2640));
                      reg2766 <= (~&$unsigned($signed(reg2608)));
                      reg2767 <= $unsigned(((forvar2693 ?
                              (reg2737 ?
                                  forvar2689 : reg2684) : reg2685[(1'h1):(1'h0)]) ?
                          (^~(8'haa)) : $signed(((8'ha3) ?
                              reg2751 : wire2582))));
                      reg2768 <= forvar2764[(3'h4):(3'h4)];
                    end
                  for (forvar2769 = (1'h0); (forvar2769 < (1'h1)); forvar2769 = (forvar2769 + (1'h1)))
                    begin
                      reg2770 <= $unsigned(((8'hb5) ?
                          ((forvar2697 ? forvar2753 : (8'hba)) ?
                              $signed(forvar2689) : (~|forvar2697)) : ($unsigned(reg2588) != reg2631)));
                      reg2771 <= $signed(((forvar2718[(2'h3):(2'h3)] ?
                              $unsigned(forvar2700) : reg2648) ?
                          {$unsigned(forvar2679)} : (~&((8'hb0) ?
                              reg2686 : reg2723))));
                    end
                end
              reg2772 <= $unsigned(reg2744);
            end
        end
    end
  always
    @(posedge clk) begin
      if ((($signed((reg2757 ?
          reg2716 : reg2664)) >= $signed({reg2586})) >> ({(~&(8'ha4))} < ($unsigned((8'hb6)) | $unsigned(reg2657)))))
        begin
          if ({($signed(reg2681) ?
                  (reg2631[(2'h3):(2'h2)] * reg2733[(1'h0):(1'h0)]) : $signed({(8'hb3)}))})
            begin
              if (reg2745)
                begin
                  if ((&(reg2693 ?
                      (~{reg2749}) : $unsigned((reg2657 ? reg2630 : (8'ha8))))))
                    begin
                      reg2773 <= $unsigned({$unsigned($unsigned(reg2697))});
                    end
                  else
                    begin
                      reg2773 <= (reg2698 + wire2670);
                      reg2774 <= reg2763;
                      reg2775 <= {(((reg2606 >> reg2739) > reg2587[(1'h1):(1'h0)]) ?
                              reg2642[(1'h0):(1'h0)] : reg2594)};
                      reg2776 <= ($unsigned({$unsigned(reg2629)}) ?
                          reg2747[(2'h2):(2'h2)] : (&reg2618));
                    end
                  for (forvar2777 = (1'h0); (forvar2777 < (1'h1)); forvar2777 = (forvar2777 + (1'h1)))
                    begin
                      reg2778 <= {((8'ha0) ? $signed((|reg2629)) : (8'h9e))};
                      reg2779 <= (-reg2654);
                      reg2780 <= (-$unsigned((reg2690 ?
                          $signed(reg2714) : reg2690[(1'h1):(1'h0)])));
                      reg2781 <= (!reg2756);
                    end
                  for (forvar2782 = (1'h0); (forvar2782 < (2'h2)); forvar2782 = (forvar2782 + (1'h1)))
                    begin
                      reg2783 <= reg2667;
                      reg2784 <= (-$signed({reg2620[(4'hb):(1'h0)]}));
                      reg2785 <= reg2656;
                    end
                end
              else
                begin
                  if (($signed((~^reg2761[(3'h6):(3'h6)])) <<< reg2649[(2'h3):(1'h0)]))
                    begin
                      reg2773 <= {((reg2635 ?
                                  {reg2733} : (reg2734 ? wire2581 : (8'ha9))) ?
                              (8'hab) : (8'hb1))};
                      reg2774 <= {$signed(reg2639)};
                    end
                  else
                    begin
                      reg2773 <= ((&$signed(reg2741)) != ((+reg2596[(1'h1):(1'h1)]) * {reg2738}));
                    end
                end
              if ((reg2705[(1'h1):(1'h0)] ?
                  $signed(wire2671) : ($signed($signed(reg2714)) | $signed(wire2672[(1'h1):(1'h0)]))))
                begin
                  if ($signed(($unsigned((^reg2716)) ?
                      reg2635[(1'h1):(1'h1)] : ((8'ha8) ~^ $signed(reg2756)))))
                    begin
                      reg2786 <= reg2648;
                      reg2787 <= (^~reg2748[(4'ha):(2'h2)]);
                      reg2788 <= (!(+reg2742[(4'hb):(3'h7)]));
                    end
                  else
                    begin
                      reg2786 <= (reg2703[(1'h1):(1'h0)] && ((~&((8'ha7) ?
                          reg2646 : reg2613)) >> ($unsigned(reg2714) ?
                          $signed(reg2594) : (reg2786 >> reg2678))));
                      reg2787 <= (^(((reg2698 ? reg2650 : reg2615) ?
                          $signed(reg2712) : (^~reg2783)) >> $unsigned(reg2707[(3'h6):(1'h0)])));
                      reg2788 <= $signed(reg2700[(4'h8):(1'h1)]);
                      reg2789 <= {(($signed(reg2592) < reg2627) ?
                              reg2758 : $signed($unsigned(reg2603)))};
                    end
                  reg2790 <= $unsigned({$unsigned((reg2743 ?
                          reg2622 : reg2602))});
                  if (reg2751[(2'h3):(1'h0)])
                    begin
                      reg2791 <= ($unsigned(reg2742) ?
                          $signed(reg2657) : ({$signed(reg2768)} <<< $signed(reg2685[(2'h2):(2'h2)])));
                      reg2792 <= reg2664;
                      reg2793 <= (((|$unsigned(reg2593)) & $signed({reg2609})) ^~ reg2607[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg2791 <= $unsigned(({reg2790} ?
                          $unsigned((!reg2722)) : {reg2592}));
                      reg2792 <= $unsigned($signed((reg2609 ~^ $unsigned(reg2598))));
                      reg2793 <= ({reg2758} ?
                          {reg2793} : ((((8'h9f) > reg2743) != (reg2726 ~^ reg2644)) < (reg2605[(3'h7):(3'h7)] - (reg2602 ?
                              reg2776 : reg2771))));
                    end
                end
              else
                begin
                  reg2786 <= (((~^reg2641) ?
                          reg2651[(2'h3):(1'h0)] : ((reg2632 || reg2743) << reg2661)) ?
                      (reg2597[(1'h0):(1'h0)] ?
                          $signed(((8'hae) <<< reg2631)) : reg2786) : (8'hb0));
                  for (forvar2787 = (1'h0); (forvar2787 < (1'h0)); forvar2787 = (forvar2787 + (1'h1)))
                    begin
                      reg2788 <= reg2627[(3'h4):(1'h0)];
                      reg2789 <= ($unsigned({$unsigned((8'ha7))}) ?
                          wire2581 : {((reg2714 ?
                                  reg2772 : reg2656) | reg2727)});
                    end
                  for (forvar2790 = (1'h0); (forvar2790 < (2'h3)); forvar2790 = (forvar2790 + (1'h1)))
                    begin
                      reg2791 <= $signed((~^reg2775[(2'h2):(1'h0)]));
                    end
                  for (forvar2792 = (1'h0); (forvar2792 < (2'h3)); forvar2792 = (forvar2792 + (1'h1)))
                    begin
                      reg2793 <= reg2743;
                      reg2794 <= $unsigned(((!{reg2704}) >> {(^~(8'ha5))}));
                    end
                end
              if ({(((reg2726 ? reg2602 : reg2692) ?
                      (8'ha6) : {(8'ha9)}) != ((+wire2668) & reg2757[(1'h1):(1'h0)]))})
                begin
                  reg2795 <= (~reg2741[(1'h1):(1'h0)]);
                  for (forvar2796 = (1'h0); (forvar2796 < (2'h3)); forvar2796 = (forvar2796 + (1'h1)))
                    begin
                      reg2797 <= (reg2743[(3'h4):(2'h2)] - $signed($unsigned(reg2644[(1'h0):(1'h0)])));
                    end
                  if ((~&$unsigned((reg2687 ? (+(8'haa)) : {reg2711}))))
                    begin
                      reg2798 <= ((reg2604 == reg2773[(3'h6):(1'h0)]) ?
                          (8'hae) : (wire2671[(1'h0):(1'h0)] ?
                              reg2748[(2'h3):(1'h1)] : (!(reg2697 <= reg2772))));
                      reg2799 <= reg2709;
                    end
                  else
                    begin
                      reg2798 <= $signed(reg2757[(2'h2):(1'h1)]);
                      reg2799 <= ({$unsigned(reg2605[(4'h8):(2'h2)])} ^~ reg2628[(3'h6):(1'h1)]);
                      reg2800 <= $unsigned(reg2633);
                    end
                end
              else
                begin
                  if ($signed(reg2652))
                    begin
                      reg2795 <= ($unsigned((reg2757[(2'h2):(2'h2)] < {reg2682})) ?
                          (8'ha7) : (^~((&reg2696) < $signed(forvar2790))));
                      reg2796 <= reg2591[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg2795 <= (+{((reg2784 ?
                              reg2693 : reg2645) ^~ $signed((8'haf)))});
                      reg2796 <= (reg2721[(2'h2):(2'h2)] < (~^($unsigned(reg2703) ?
                          $signed(reg2778) : reg2654)));
                      reg2797 <= reg2590;
                      reg2798 <= forvar2792[(4'h8):(1'h1)];
                    end
                  for (forvar2799 = (1'h0); (forvar2799 < (1'h1)); forvar2799 = (forvar2799 + (1'h1)))
                    begin
                      reg2800 <= wire2580[(2'h2):(1'h0)];
                      reg2801 <= reg2748;
                      reg2802 <= (^reg2687);
                      reg2803 <= ((-($unsigned(reg2702) | (reg2773 ?
                          reg2737 : reg2623))) <<< (((-reg2742) ?
                          (|reg2623) : reg2590) & ($unsigned((8'hae)) ?
                          $signed(wire2583) : (reg2617 ? reg2613 : reg2597))));
                    end
                  if ({reg2796})
                    begin
                      reg2804 <= (~|$unsigned($signed({(8'hb9)})));
                      reg2805 <= reg2763[(2'h2):(1'h1)];
                      reg2806 <= (~&reg2788);
                    end
                  else
                    begin
                      reg2804 <= reg2602[(4'hb):(2'h3)];
                      reg2805 <= reg2709;
                    end
                  for (forvar2807 = (1'h0); (forvar2807 < (2'h3)); forvar2807 = (forvar2807 + (1'h1)))
                    begin
                      reg2808 <= (+reg2706);
                      reg2809 <= reg2622;
                      reg2810 <= reg2701[(4'hd):(4'h8)];
                      reg2811 <= (reg2608[(2'h3):(2'h3)] >>> (8'ha0));
                    end
                end
              for (forvar2812 = (1'h0); (forvar2812 < (1'h1)); forvar2812 = (forvar2812 + (1'h1)))
                begin
                  if ($signed(($unsigned((~|reg2713)) ? reg2587 : wire2583)))
                    begin
                      reg2813 <= ($unsigned(((^reg2704) && reg2648)) ?
                          reg2695[(2'h3):(1'h1)] : ($unsigned(reg2706[(1'h0):(1'h0)]) >> ((8'haf) && reg2758[(2'h3):(1'h0)])));
                      reg2814 <= $unsigned($unsigned(reg2720[(2'h2):(1'h0)]));
                      reg2815 <= reg2783;
                      reg2816 <= {$signed(({reg2610} ?
                              (reg2813 >>> reg2789) : $signed(reg2791)))};
                    end
                  else
                    begin
                      reg2813 <= $signed($signed(($signed(reg2641) ?
                          $signed(reg2757) : $unsigned(reg2686))));
                      reg2814 <= (reg2803 ?
                          reg2794[(4'hc):(2'h2)] : (wire2669 >>> (8'ha6)));
                    end
                  if (wire2668[(4'h9):(4'h8)])
                    begin
                      reg2817 <= ((&reg2663) <= $unsigned({(reg2708 ?
                              (8'hb2) : reg2786)}));
                      reg2818 <= $signed((~^(|(reg2622 > (8'hb4)))));
                    end
                  else
                    begin
                      reg2817 <= $signed(reg2633[(2'h3):(2'h2)]);
                      reg2818 <= reg2768[(2'h2):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar2773 = (1'h0); (forvar2773 < (1'h0)); forvar2773 = (forvar2773 + (1'h1)))
                begin
                  for (forvar2774 = (1'h0); (forvar2774 < (2'h2)); forvar2774 = (forvar2774 + (1'h1)))
                    begin
                      reg2775 <= $signed({{(forvar2812 >>> reg2783)}});
                      reg2776 <= $signed((~(~|$signed((8'ha9)))));
                    end
                  reg2777 <= (forvar2773[(4'ha):(2'h3)] ?
                      ($unsigned((|reg2618)) >= forvar2777[(2'h3):(1'h1)]) : ($signed($signed(reg2655)) ?
                          ({wire2582} >> (reg2635 ?
                              reg2602 : (8'ha7))) : reg2805[(4'h8):(3'h5)]));
                  reg2778 <= (8'h9c);
                end
            end
          reg2819 <= reg2752[(4'h8):(3'h6)];
          for (forvar2820 = (1'h0); (forvar2820 < (2'h2)); forvar2820 = (forvar2820 + (1'h1)))
            begin
              if (($unsigned($unsigned((~^reg2783))) ^~ $unsigned($unsigned(reg2738[(3'h4):(3'h4)]))))
                begin
                  for (forvar2821 = (1'h0); (forvar2821 < (1'h1)); forvar2821 = (forvar2821 + (1'h1)))
                    begin
                      reg2822 <= ($signed(reg2735) ?
                          ((&$unsigned(reg2775)) > $unsigned({reg2690})) : ({(reg2621 ?
                                  reg2799 : (8'had))} << $signed((^(8'hb4)))));
                      reg2823 <= $unsigned((({(8'h9d)} || {(8'ha8)}) | ((reg2818 ?
                          reg2619 : reg2771) >>> $signed((8'ha9)))));
                      reg2824 <= ((($signed(reg2649) ^~ $signed(reg2631)) ?
                              (~|$unsigned(reg2641)) : ((~&reg2604) >= $unsigned(reg2605))) ?
                          (-wire2669[(3'h5):(1'h0)]) : reg2725[(3'h6):(3'h6)]);
                    end
                  reg2825 <= (wire2583[(1'h1):(1'h1)] < $unsigned(reg2817));
                  for (forvar2826 = (1'h0); (forvar2826 < (1'h0)); forvar2826 = (forvar2826 + (1'h1)))
                    begin
                      reg2827 <= reg2693;
                    end
                end
              else
                begin
                  reg2821 <= ((^(|(reg2754 == reg2609))) - {reg2765});
                  for (forvar2822 = (1'h0); (forvar2822 < (2'h3)); forvar2822 = (forvar2822 + (1'h1)))
                    begin
                      reg2823 <= (reg2657[(1'h0):(1'h0)] != (!($unsigned((8'hb5)) ?
                          (!(8'hb1)) : $unsigned(reg2706))));
                      reg2824 <= reg2704[(1'h1):(1'h1)];
                      reg2825 <= (((~$signed((8'ha1))) ?
                          ($signed(reg2659) ?
                              (reg2729 ?
                                  reg2682 : reg2711) : reg2666[(4'hc):(1'h1)]) : (+reg2592[(4'ha):(3'h7)])) >= (8'ha9));
                    end
                  for (forvar2826 = (1'h0); (forvar2826 < (2'h2)); forvar2826 = (forvar2826 + (1'h1)))
                    begin
                      reg2827 <= reg2797;
                      reg2828 <= (reg2683[(3'h6):(3'h4)] ?
                          $signed({{reg2651}}) : (reg2784[(1'h1):(1'h0)] ?
                              reg2724[(4'h9):(1'h0)] : {(reg2589 >= reg2787)}));
                      reg2829 <= ((reg2591[(4'hc):(4'hc)] ^ reg2686[(3'h5):(3'h4)]) && $unsigned(($signed((8'had)) != {reg2683})));
                    end
                end
              if ((-{reg2702[(1'h0):(1'h0)]}))
                begin
                  if ({(reg2740 ?
                          {(reg2741 != (8'h9c))} : ((~|reg2794) >= $unsigned(reg2651)))})
                    begin
                      reg2830 <= (((reg2681 ^ (wire2669 ? reg2744 : reg2768)) ?
                              $signed(reg2606[(4'h8):(3'h7)]) : reg2699) ?
                          (~$unsigned($unsigned((8'hb1)))) : reg2663);
                    end
                  else
                    begin
                      reg2830 <= (reg2712 << $unsigned(($unsigned(reg2779) >= (reg2622 ~^ reg2588))));
                      reg2831 <= {($unsigned($unsigned(reg2639)) || ($unsigned(reg2749) ?
                              (~&reg2799) : (^(8'hae))))};
                      reg2832 <= reg2703[(1'h0):(1'h0)];
                    end
                  if ((((-reg2629[(1'h0):(1'h0)]) | reg2823) ?
                      $unsigned($signed(reg2611)) : ((^reg2612) ?
                          $unsigned((^~forvar2790)) : (8'hb7))))
                    begin
                      reg2833 <= (reg2641 ?
                          (&reg2603[(4'hd):(3'h4)]) : (reg2783 ?
                              ((reg2829 ? reg2682 : reg2780) ?
                                  (!(8'hb4)) : reg2793[(3'h4):(2'h3)]) : ((reg2763 * reg2700) ~^ {reg2751})));
                    end
                  else
                    begin
                      reg2833 <= ({(reg2606 == (^~reg2614))} ?
                          (!(|(!forvar2807))) : reg2617[(3'h5):(1'h0)]);
                      reg2834 <= ($signed(((reg2589 << reg2810) ^ ((8'hb1) >>> (8'hba)))) * reg2590[(1'h1):(1'h0)]);
                      reg2835 <= $unsigned(reg2791);
                      reg2836 <= (reg2793 > forvar2796[(3'h6):(3'h4)]);
                    end
                end
              else
                begin
                  if ({reg2589})
                    begin
                      reg2830 <= $signed($signed($signed({(8'haa)})));
                      reg2831 <= {((reg2767 ?
                                  (reg2620 ? reg2646 : reg2752) : reg2619) ?
                              reg2742[(4'h9):(2'h2)] : {(8'hb4)})};
                    end
                  else
                    begin
                      reg2830 <= ((^~$unsigned((reg2663 ~^ (8'ha8)))) >>> (reg2622[(3'h4):(2'h2)] ?
                          (8'ha5) : $unsigned((|forvar2822))));
                    end
                end
              if (reg2818[(1'h1):(1'h1)])
                begin
                  for (forvar2837 = (1'h0); (forvar2837 < (2'h3)); forvar2837 = (forvar2837 + (1'h1)))
                    begin
                      reg2838 <= ((forvar2790 ?
                          reg2635 : $unsigned($unsigned(reg2830))) >> $signed(reg2750[(2'h2):(1'h1)]));
                    end
                  reg2839 <= (reg2710[(1'h0):(1'h0)] | $unsigned($signed((reg2814 < reg2805))));
                  for (forvar2840 = (1'h0); (forvar2840 < (1'h0)); forvar2840 = (forvar2840 + (1'h1)))
                    begin
                      reg2841 <= $signed(($signed($signed(reg2684)) == (((8'h9e) ?
                              reg2831 : reg2738) ?
                          $signed(reg2755) : (reg2721 ? wire2670 : reg2747))));
                      reg2842 <= $signed((!$unsigned((reg2789 ?
                          forvar2807 : (8'ha2)))));
                      reg2843 <= {({$unsigned(forvar2821)} ?
                              $signed($signed(reg2799)) : $signed($unsigned(reg2763)))};
                    end
                end
              else
                begin
                  if (({(^forvar2826[(1'h1):(1'h1)])} ?
                      reg2722 : (((~forvar2773) * $signed(wire2581)) <= (~^(reg2739 ?
                          reg2692 : (8'haf))))))
                    begin
                      reg2837 <= $unsigned((reg2589 & (~^(^~reg2799))));
                      reg2838 <= (wire2581[(1'h0):(1'h0)] ^ (({forvar2837} + reg2618[(4'h9):(3'h4)]) > reg2748));
                      reg2839 <= {reg2801};
                      reg2840 <= (forvar2820 ?
                          ($signed($signed(reg2736)) ^ $signed(reg2613)) : $unsigned($signed(((8'haf) > reg2597))));
                    end
                  else
                    begin
                      reg2837 <= ($signed(((8'hb5) ?
                              $unsigned(reg2746) : reg2648)) ?
                          ({reg2827} ?
                              {reg2815} : (wire2671[(1'h0):(1'h0)] > reg2761)) : (8'ha8));
                      reg2838 <= $unsigned(reg2678[(2'h2):(1'h0)]);
                      reg2839 <= (&((^~reg2778[(1'h1):(1'h1)]) ?
                          (-((8'ha8) & reg2659)) : ($signed(reg2759) ?
                              (~|reg2700) : (reg2791 ? reg2756 : reg2699))));
                    end
                  for (forvar2841 = (1'h0); (forvar2841 < (1'h1)); forvar2841 = (forvar2841 + (1'h1)))
                    begin
                      reg2842 <= (~|$signed({reg2593[(4'ha):(4'h9)]}));
                      reg2843 <= (!reg2811);
                    end
                  if (reg2795)
                    begin
                      reg2844 <= ($signed(((forvar2807 > reg2630) ?
                          (reg2757 ? reg2691 : reg2722) : (reg2700 ?
                              forvar2840 : reg2696))) >= (!$signed($unsigned(reg2825))));
                      reg2845 <= {reg2719};
                      reg2846 <= (~(~^reg2636));
                    end
                  else
                    begin
                      reg2844 <= (($signed(reg2802) < reg2775) << (($signed(reg2686) >>> reg2621) == reg2825));
                    end
                  for (forvar2847 = (1'h0); (forvar2847 < (1'h0)); forvar2847 = (forvar2847 + (1'h1)))
                    begin
                      reg2848 <= reg2657[(3'h6):(2'h2)];
                      reg2849 <= $signed(forvar2796[(3'h7):(3'h7)]);
                      reg2850 <= reg2608;
                      reg2851 <= (-{($unsigned((8'haf)) ?
                              (&(8'ha9)) : (|reg2823))});
                    end
                end
            end
          if ({(({(8'hae)} ~^ (8'ha9)) ?
                  ((forvar2787 >>> reg2612) < reg2765) : (!reg2779))})
            begin
              for (forvar2852 = (1'h0); (forvar2852 < (2'h2)); forvar2852 = (forvar2852 + (1'h1)))
                begin
                  for (forvar2853 = (1'h0); (forvar2853 < (2'h3)); forvar2853 = (forvar2853 + (1'h1)))
                    begin
                      reg2854 <= $signed($unsigned($unsigned((!reg2848))));
                      reg2855 <= {((~wire2580[(4'h8):(1'h0)]) ?
                              $signed(reg2771) : reg2681)};
                      reg2856 <= reg2831;
                    end
                  for (forvar2857 = (1'h0); (forvar2857 < (1'h0)); forvar2857 = (forvar2857 + (1'h1)))
                    begin
                      reg2858 <= $signed($signed(($unsigned(reg2792) ?
                          ((8'ha5) ?
                              reg2808 : reg2834) : (reg2796 == reg2739))));
                    end
                end
            end
          else
            begin
              for (forvar2852 = (1'h0); (forvar2852 < (1'h1)); forvar2852 = (forvar2852 + (1'h1)))
                begin
                  for (forvar2853 = (1'h0); (forvar2853 < (2'h3)); forvar2853 = (forvar2853 + (1'h1)))
                    begin
                      reg2854 <= ({$unsigned((reg2799 ?
                              reg2843 : forvar2826))} <= $unsigned($unsigned($signed(reg2759))));
                      reg2855 <= $unsigned($signed(wire2671[(1'h1):(1'h0)]));
                      reg2856 <= (^reg2608);
                      reg2857 <= $signed(reg2741[(4'h9):(2'h2)]);
                    end
                  for (forvar2858 = (1'h0); (forvar2858 < (1'h1)); forvar2858 = (forvar2858 + (1'h1)))
                    begin
                      reg2859 <= ((reg2833[(3'h7):(2'h3)] - reg2857) & ($unsigned((wire2581 + reg2765)) ?
                          reg2694[(2'h3):(2'h3)] : reg2712[(2'h2):(1'h1)]));
                      reg2860 <= reg2825;
                      reg2861 <= {(~(~^(^reg2715)))};
                    end
                end
              for (forvar2862 = (1'h0); (forvar2862 < (1'h1)); forvar2862 = (forvar2862 + (1'h1)))
                begin
                  reg2863 <= (reg2694 ?
                      (reg2627[(3'h4):(1'h1)] ^~ ((forvar2852 ?
                          reg2667 : reg2838) * $unsigned(reg2700))) : (8'ha8));
                end
              for (forvar2864 = (1'h0); (forvar2864 < (2'h2)); forvar2864 = (forvar2864 + (1'h1)))
                begin
                  for (forvar2865 = (1'h0); (forvar2865 < (2'h2)); forvar2865 = (forvar2865 + (1'h1)))
                    begin
                      reg2866 <= (8'ha1);
                    end
                  for (forvar2867 = (1'h0); (forvar2867 < (2'h3)); forvar2867 = (forvar2867 + (1'h1)))
                    begin
                      reg2868 <= (+reg2653);
                      reg2869 <= $signed(reg2789[(4'h8):(3'h5)]);
                    end
                  for (forvar2870 = (1'h0); (forvar2870 < (2'h3)); forvar2870 = (forvar2870 + (1'h1)))
                    begin
                      reg2871 <= {($unsigned((wire2584 < reg2861)) * (!$signed(reg2731)))};
                      reg2872 <= $unsigned((~($signed(reg2628) ?
                          reg2731[(1'h0):(1'h0)] : ((8'hb1) | reg2661))));
                      reg2873 <= {(^$signed($signed(reg2818)))};
                      reg2874 <= $signed(reg2740[(1'h0):(1'h0)]);
                    end
                end
              if ((-reg2777[(3'h4):(3'h4)]))
                begin
                  for (forvar2875 = (1'h0); (forvar2875 < (2'h2)); forvar2875 = (forvar2875 + (1'h1)))
                    begin
                      reg2876 <= (reg2635 ?
                          (~&((forvar2857 && reg2827) ?
                              (reg2739 & reg2809) : {reg2740})) : (~|((reg2808 > (8'ha8)) ?
                              (~reg2816) : ((8'h9e) ^ forvar2821))));
                      reg2877 <= reg2662;
                    end
                end
              else
                begin
                  for (forvar2875 = (1'h0); (forvar2875 < (2'h2)); forvar2875 = (forvar2875 + (1'h1)))
                    begin
                      reg2876 <= (8'ha3);
                    end
                  for (forvar2877 = (1'h0); (forvar2877 < (2'h3)); forvar2877 = (forvar2877 + (1'h1)))
                    begin
                      reg2878 <= $unsigned($signed(((reg2790 ?
                          reg2695 : reg2655) - $unsigned((8'hb1)))));
                    end
                  reg2879 <= forvar2840;
                end
            end
        end
      else
        begin
          for (forvar2773 = (1'h0); (forvar2773 < (1'h1)); forvar2773 = (forvar2773 + (1'h1)))
            begin
              for (forvar2774 = (1'h0); (forvar2774 < (1'h0)); forvar2774 = (forvar2774 + (1'h1)))
                begin
                  if (reg2650)
                    begin
                      reg2775 <= {$signed($signed(reg2725))};
                      reg2776 <= (((~(reg2618 ^ reg2866)) - reg2731[(1'h0):(1'h0)]) > $unsigned($unsigned((reg2731 ?
                          reg2832 : reg2588))));
                      reg2777 <= (&(reg2768[(4'hc):(3'h6)] ^ $signed(reg2617)));
                      reg2778 <= {reg2805[(1'h1):(1'h1)]};
                    end
                  else
                    begin
                      reg2775 <= (~&$signed(reg2808));
                      reg2776 <= reg2825[(2'h2):(2'h2)];
                    end
                  for (forvar2779 = (1'h0); (forvar2779 < (2'h3)); forvar2779 = (forvar2779 + (1'h1)))
                    begin
                      reg2780 <= reg2787[(3'h7):(2'h3)];
                      reg2781 <= $signed({reg2800[(1'h0):(1'h0)]});
                      reg2782 <= $signed((-(+(reg2604 ? reg2819 : reg2667))));
                      reg2783 <= (!($signed((reg2795 ? reg2879 : forvar2875)) ?
                          (((8'ha6) ?
                              reg2595 : (8'ha6)) < $unsigned(reg2782)) : $signed(((8'hb7) ?
                              forvar2790 : reg2773))));
                    end
                  for (forvar2784 = (1'h0); (forvar2784 < (2'h3)); forvar2784 = (forvar2784 + (1'h1)))
                    begin
                      reg2785 <= $unsigned($signed(((~|reg2691) << {forvar2862})));
                      reg2786 <= ($signed(wire2582) ?
                          {{(~reg2625)}} : $signed(reg2871));
                      reg2787 <= ($signed(($signed((8'ha3)) ?
                          (reg2796 && reg2681) : reg2828[(2'h3):(2'h2)])) && ($unsigned({reg2645}) == reg2845));
                    end
                end
              reg2788 <= reg2605;
              if ({$unsigned({{forvar2853}})})
                begin
                  for (forvar2789 = (1'h0); (forvar2789 < (1'h0)); forvar2789 = (forvar2789 + (1'h1)))
                    begin
                      reg2790 <= (~|(^~reg2660[(2'h2):(1'h1)]));
                      reg2791 <= (((~|(|reg2841)) >= reg2827) ?
                          $unsigned($unsigned((forvar2826 * reg2627))) : {forvar2782[(3'h5):(3'h4)]});
                      reg2792 <= reg2713[(3'h5):(2'h3)];
                    end
                  if ((reg2810[(3'h7):(3'h6)] ?
                      {$signed(forvar2777)} : forvar2784))
                    begin
                      reg2793 <= $unsigned(($unsigned($signed(reg2634)) & reg2748[(3'h5):(3'h5)]));
                      reg2794 <= reg2729;
                      reg2795 <= reg2784[(3'h6):(2'h3)];
                    end
                  else
                    begin
                      reg2793 <= reg2742;
                      reg2794 <= (($signed({reg2818}) || {(+reg2876)}) <<< {((~^forvar2787) ?
                              (reg2687 - reg2857) : (reg2756 || reg2608))});
                      reg2795 <= ((8'hb0) ?
                          {((reg2619 ?
                                  (8'hb6) : forvar2875) + $unsigned(reg2604))} : $signed((~&(~^forvar2790))));
                      reg2796 <= $unsigned((~&forvar2837[(3'h6):(3'h6)]));
                    end
                end
              else
                begin
                  if ((8'had))
                    begin
                      reg2789 <= ((|$signed($unsigned(reg2587))) ^~ reg2811[(4'h9):(3'h4)]);
                      reg2790 <= forvar2852;
                    end
                  else
                    begin
                      reg2789 <= (({$unsigned(reg2860)} << $unsigned((reg2618 >>> reg2641))) * $unsigned((|(8'h9e))));
                      reg2790 <= {(~(forvar2773 <= reg2779))};
                      reg2791 <= (^~$signed((!$signed(reg2749))));
                      reg2792 <= reg2718;
                    end
                  for (forvar2793 = (1'h0); (forvar2793 < (2'h3)); forvar2793 = (forvar2793 + (1'h1)))
                    begin
                      reg2794 <= wire2668[(3'h7):(3'h6)];
                      reg2795 <= $unsigned(reg2767[(4'h8):(1'h0)]);
                      reg2796 <= $signed(((((8'hb7) && reg2851) && $signed(reg2796)) ?
                          reg2614 : $unsigned(reg2810)));
                      reg2797 <= (reg2604[(3'h5):(3'h4)] ?
                          $unsigned((+{reg2851})) : reg2705);
                    end
                  if ((~^(^~((reg2589 ? (8'h9e) : reg2728) ?
                      $unsigned(reg2878) : $unsigned(reg2710)))))
                    begin
                      reg2798 <= reg2791[(1'h0):(1'h0)];
                      reg2799 <= (reg2701[(4'h8):(3'h5)] ?
                          ($signed((~|wire2669)) ^ ((reg2777 ^ (8'ha1)) ?
                              (forvar2812 ?
                                  reg2818 : (8'ha6)) : reg2739)) : {$signed((reg2877 ?
                                  forvar2774 : forvar2784))});
                    end
                  else
                    begin
                      reg2798 <= reg2623;
                    end
                  for (forvar2800 = (1'h0); (forvar2800 < (2'h2)); forvar2800 = (forvar2800 + (1'h1)))
                    begin
                      reg2801 <= {($signed((reg2861 ? (8'ha1) : (8'hb6))) ?
                              $signed($unsigned(reg2755)) : $unsigned({reg2873}))};
                      reg2802 <= $unsigned((^{reg2748[(3'h5):(2'h2)]}));
                    end
                end
              for (forvar2803 = (1'h0); (forvar2803 < (1'h1)); forvar2803 = (forvar2803 + (1'h1)))
                begin
                  reg2804 <= (reg2740[(1'h1):(1'h1)] ?
                      $unsigned((^$unsigned(forvar2877))) : ((!reg2758) >= forvar2841[(4'ha):(3'h7)]));
                end
            end
          if ($unsigned($unsigned((^reg2795))))
            begin
              if ((!$unsigned((reg2860[(4'hb):(1'h1)] ?
                  {reg2784} : $signed(reg2832)))))
                begin
                  reg2805 <= {reg2723[(1'h0):(1'h0)]};
                  if ((&{{(forvar2857 >> reg2781)}}))
                    begin
                      reg2806 <= ((+((8'hab) ?
                          wire2673 : reg2765)) && (~^{{reg2825}}));
                      reg2807 <= reg2791[(4'ha):(2'h3)];
                    end
                  else
                    begin
                      reg2806 <= {reg2798};
                      reg2807 <= $unsigned($unsigned((|reg2727)));
                      reg2808 <= $signed({(reg2717 ?
                              $signed((8'ha4)) : reg2589[(1'h0):(1'h0)])});
                    end
                  for (forvar2809 = (1'h0); (forvar2809 < (2'h2)); forvar2809 = (forvar2809 + (1'h1)))
                    begin
                      reg2810 <= $signed($unsigned($signed((reg2723 ?
                          reg2738 : reg2858))));
                      reg2811 <= ($signed((reg2606 | forvar2870[(3'h6):(2'h2)])) & reg2774[(2'h3):(2'h2)]);
                      reg2812 <= (reg2846 * ({(forvar2865 ~^ (8'had))} ?
                          reg2828[(1'h1):(1'h0)] : $unsigned((~&(8'had)))));
                      reg2813 <= reg2723[(1'h0):(1'h0)];
                    end
                  for (forvar2814 = (1'h0); (forvar2814 < (1'h0)); forvar2814 = (forvar2814 + (1'h1)))
                    begin
                      reg2815 <= $signed($unsigned($unsigned({reg2812})));
                      reg2816 <= (~$unsigned(({reg2809} ?
                          forvar2877 : reg2597)));
                      reg2817 <= $signed((~|{(8'ha0)}));
                    end
                end
              else
                begin
                  for (forvar2805 = (1'h0); (forvar2805 < (1'h0)); forvar2805 = (forvar2805 + (1'h1)))
                    begin
                      reg2806 <= reg2873;
                      reg2807 <= {$signed((8'ha8))};
                      reg2808 <= $signed($signed($unsigned((reg2729 < reg2777))));
                    end
                end
              if ($unsigned(reg2741[(4'ha):(2'h3)]))
                begin
                  for (forvar2818 = (1'h0); (forvar2818 < (2'h2)); forvar2818 = (forvar2818 + (1'h1)))
                    begin
                      reg2819 <= reg2803;
                      reg2820 <= {$unsigned((reg2834 ?
                              forvar2857 : $unsigned(reg2835)))};
                    end
                  reg2821 <= (reg2633[(1'h1):(1'h1)] ?
                      (+reg2741[(4'h8):(3'h5)]) : $signed((reg2730[(2'h2):(1'h1)] < $signed((8'hb3)))));
                  if (reg2833)
                    begin
                      reg2822 <= reg2759[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg2822 <= $signed(reg2698);
                      reg2823 <= (reg2863 < $signed(reg2733));
                    end
                  if ((reg2718[(3'h5):(1'h0)] ?
                      (^~$unsigned((^reg2823))) : (({(8'hb8)} - reg2658[(1'h0):(1'h0)]) == ((8'ha5) ?
                          $signed((8'hb0)) : {(8'hba)}))))
                    begin
                      reg2824 <= {($unsigned((reg2800 ?
                              reg2874 : (8'h9d))) >> (~(forvar2820 - wire2669)))};
                      reg2825 <= reg2650[(1'h1):(1'h1)];
                      reg2826 <= reg2620;
                    end
                  else
                    begin
                      reg2824 <= $unsigned($unsigned(((reg2818 <= reg2755) <= (~|reg2844))));
                    end
                end
              else
                begin
                  for (forvar2818 = (1'h0); (forvar2818 < (2'h2)); forvar2818 = (forvar2818 + (1'h1)))
                    begin
                      reg2819 <= {$signed((^~$signed(reg2717)))};
                      reg2820 <= (&(!reg2753));
                      reg2821 <= $unsigned((8'ha9));
                    end
                  for (forvar2822 = (1'h0); (forvar2822 < (2'h3)); forvar2822 = (forvar2822 + (1'h1)))
                    begin
                      reg2823 <= reg2648;
                    end
                  if (reg2681[(1'h0):(1'h0)])
                    begin
                      reg2824 <= $signed($unsigned(forvar2793));
                      reg2825 <= $unsigned($unsigned($unsigned((reg2656 ?
                          reg2704 : reg2868))));
                      reg2826 <= (forvar2777[(1'h1):(1'h1)] ?
                          $signed(((reg2685 ? reg2778 : wire2583) ?
                              ((8'ha3) >= (8'hb0)) : $unsigned(reg2771))) : $unsigned(((-forvar2837) ?
                              {reg2607} : {reg2837})));
                    end
                  else
                    begin
                      reg2824 <= reg2856;
                      reg2825 <= (^~{$signed(reg2845[(3'h6):(1'h1)])});
                    end
                  for (forvar2827 = (1'h0); (forvar2827 < (1'h1)); forvar2827 = (forvar2827 + (1'h1)))
                    begin
                      reg2828 <= $signed((($unsigned(reg2685) ?
                              (!forvar2773) : (reg2845 ? reg2683 : reg2596)) ?
                          reg2758[(2'h3):(1'h0)] : ((^~reg2825) ?
                              ((8'ha9) + reg2815) : (reg2718 || reg2615))));
                      reg2829 <= reg2587[(1'h1):(1'h0)];
                      reg2830 <= {$unsigned((+wire2583[(1'h1):(1'h1)]))};
                    end
                end
              reg2831 <= reg2707[(3'h6):(2'h2)];
              reg2832 <= (8'hb4);
            end
          else
            begin
              if ((~^wire2673[(4'hc):(3'h7)]))
                begin
                  if ($signed({(reg2840 ?
                          (reg2597 != reg2784) : ((8'ha5) <<< reg2644))}))
                    begin
                      reg2805 <= (~^reg2686[(3'h4):(2'h2)]);
                      reg2806 <= reg2617;
                    end
                  else
                    begin
                      reg2805 <= $unsigned(reg2778[(1'h0):(1'h0)]);
                      reg2806 <= reg2770;
                    end
                  if (reg2595)
                    begin
                      reg2807 <= {$signed((reg2838[(4'h8):(1'h0)] >> $unsigned(reg2587)))};
                      reg2808 <= forvar2796[(4'hc):(3'h5)];
                      reg2809 <= (reg2636[(1'h0):(1'h0)] + reg2703[(1'h0):(1'h0)]);
                      reg2810 <= $unsigned($signed($unsigned($unsigned(reg2602))));
                    end
                  else
                    begin
                      reg2807 <= $unsigned($signed($signed((reg2738 ?
                          wire2670 : reg2828))));
                      reg2808 <= reg2855;
                      reg2809 <= $unsigned((reg2772[(3'h4):(3'h4)] ?
                          (reg2798 ?
                              wire2581[(1'h1):(1'h1)] : ((8'ha0) <<< reg2828)) : (^~$signed(wire2668))));
                    end
                  for (forvar2811 = (1'h0); (forvar2811 < (2'h2)); forvar2811 = (forvar2811 + (1'h1)))
                    begin
                      reg2812 <= {{(|(reg2845 && reg2695))}};
                    end
                end
              else
                begin
                  for (forvar2805 = (1'h0); (forvar2805 < (1'h1)); forvar2805 = (forvar2805 + (1'h1)))
                    begin
                      reg2806 <= (8'ha9);
                      reg2807 <= (-$signed(((reg2640 ?
                          reg2589 : reg2827) && {reg2857})));
                      reg2808 <= wire2583[(2'h2):(1'h0)];
                      reg2809 <= reg2736[(2'h3):(2'h3)];
                    end
                end
              if (reg2801)
                begin
                  for (forvar2813 = (1'h0); (forvar2813 < (2'h2)); forvar2813 = (forvar2813 + (1'h1)))
                    begin
                      reg2814 <= $unsigned(($unsigned(wire2672[(1'h0):(1'h0)]) ^ {(reg2805 ?
                              reg2603 : (8'hb7))}));
                      reg2815 <= $unsigned($unsigned(($signed(reg2705) >> {reg2653})));
                      reg2816 <= (^$signed($signed($signed(reg2702))));
                      reg2817 <= reg2806[(4'h8):(4'h8)];
                    end
                  for (forvar2818 = (1'h0); (forvar2818 < (1'h1)); forvar2818 = (forvar2818 + (1'h1)))
                    begin
                      reg2819 <= ($unsigned(forvar2847) ?
                          ((|(!reg2742)) ^ (reg2793 ?
                              (~&forvar2827) : $unsigned(reg2663))) : {(~^(reg2611 ?
                                  reg2731 : reg2860))});
                      reg2820 <= {{(~reg2659)}};
                    end
                  for (forvar2821 = (1'h0); (forvar2821 < (2'h2)); forvar2821 = (forvar2821 + (1'h1)))
                    begin
                      reg2822 <= reg2840[(4'ha):(1'h1)];
                    end
                end
              else
                begin
                  if ((!reg2608))
                    begin
                      reg2813 <= ((!reg2642) ?
                          $unsigned($signed(((8'ha0) <= reg2739))) : ((wire2585[(1'h0):(1'h0)] >= $signed(reg2777)) ?
                              $signed($unsigned(reg2719)) : $unsigned((forvar2777 ~^ (8'hb9)))));
                      reg2814 <= (({reg2617} >> $signed((forvar2865 + reg2684))) ~^ (-$unsigned(((8'haa) ?
                          reg2719 : forvar2818))));
                      reg2815 <= ({$unsigned($unsigned(reg2725))} ~^ reg2591[(3'h7):(3'h4)]);
                    end
                  else
                    begin
                      reg2813 <= ($signed({$signed(reg2767)}) < $signed((+$unsigned(reg2774))));
                    end
                  for (forvar2816 = (1'h0); (forvar2816 < (2'h2)); forvar2816 = (forvar2816 + (1'h1)))
                    begin
                      reg2817 <= {$unsigned((reg2700 ?
                              $signed(reg2608) : $signed(reg2786)))};
                      reg2818 <= {((-forvar2782) - (reg2786[(4'ha):(3'h7)] ?
                              (reg2846 ? reg2868 : reg2715) : (8'hb5)))};
                      reg2819 <= $unsigned(($unsigned($signed(reg2629)) & (8'hb9)));
                      reg2820 <= ((~((wire2672 << reg2825) ?
                              reg2835[(2'h3):(1'h0)] : $signed(reg2655))) ?
                          $signed((~&$signed((8'ha6)))) : ($signed(reg2812) ?
                              ((reg2738 << forvar2857) << (^reg2837)) : (|((8'hba) ?
                                  reg2741 : reg2805))));
                    end
                end
            end
          for (forvar2833 = (1'h0); (forvar2833 < (1'h0)); forvar2833 = (forvar2833 + (1'h1)))
            begin
              if (reg2725[(3'h6):(1'h1)])
                begin
                  if ((((reg2693[(3'h4):(1'h0)] | reg2789) ?
                          forvar2865 : ((^reg2711) ?
                              (-reg2641) : ((8'hb3) <<< reg2768))) ?
                      $signed($unsigned((~&reg2662))) : ((^~(reg2809 * reg2855)) ?
                          $signed(wire2585[(1'h1):(1'h1)]) : reg2791)))
                    begin
                      reg2834 <= (((~$signed(forvar2858)) ?
                              ({wire2580} ?
                                  $signed((8'hb5)) : (~(8'ha8))) : reg2786) ?
                          reg2586 : (reg2828[(2'h2):(2'h2)] <= (reg2738[(3'h6):(2'h2)] ?
                              (|reg2838) : {reg2714})));
                      reg2835 <= $signed({reg2858[(3'h7):(1'h0)]});
                    end
                  else
                    begin
                      reg2834 <= ((|reg2738[(4'h9):(3'h4)]) ?
                          (forvar2782 * $unsigned(reg2586[(1'h0):(1'h0)])) : {reg2785[(3'h5):(1'h0)]});
                      reg2835 <= $unsigned(((((8'h9d) | reg2684) != $unsigned(reg2614)) < $signed((reg2725 ?
                          (8'ha8) : forvar2827))));
                      reg2836 <= (^(^reg2807[(3'h6):(1'h0)]));
                      reg2837 <= reg2779;
                    end
                end
              else
                begin
                  for (forvar2834 = (1'h0); (forvar2834 < (1'h1)); forvar2834 = (forvar2834 + (1'h1)))
                    begin
                      reg2835 <= ($signed((!(reg2705 >>> reg2630))) ?
                          ($unsigned($signed(reg2863)) ?
                              $signed($signed((8'hb5))) : ($unsigned(forvar2827) || (reg2777 ?
                                  reg2659 : reg2762))) : reg2845);
                      reg2836 <= forvar2805;
                      reg2837 <= ($signed($unsigned((reg2642 - reg2831))) ?
                          $unsigned(($signed(reg2727) - reg2763)) : ((&reg2650) ~^ ((8'ha8) <<< reg2621)));
                      reg2838 <= $unsigned(reg2821);
                    end
                  reg2839 <= $unsigned(reg2700);
                end
            end
          if ((^~$signed(((reg2786 ? reg2812 : (8'haa)) >> (~^reg2723)))))
            begin
              reg2840 <= {reg2871[(3'h6):(2'h3)]};
            end
          else
            begin
              for (forvar2840 = (1'h0); (forvar2840 < (2'h2)); forvar2840 = (forvar2840 + (1'h1)))
                begin
                  if (reg2661[(4'ha):(3'h7)])
                    begin
                      reg2841 <= $signed($unsigned(($signed(forvar2827) ?
                          $unsigned(reg2838) : (|(8'hb4)))));
                    end
                  else
                    begin
                      reg2841 <= $signed((8'hab));
                      reg2842 <= (!(forvar2790 | $signed($unsigned(reg2815))));
                    end
                  for (forvar2843 = (1'h0); (forvar2843 < (1'h1)); forvar2843 = (forvar2843 + (1'h1)))
                    begin
                      reg2844 <= ((8'hb2) - reg2649[(1'h1):(1'h1)]);
                      reg2845 <= ((|(reg2744 ?
                          wire2581[(1'h0):(1'h0)] : {reg2824})) >>> $signed($signed(reg2615[(3'h6):(1'h1)])));
                    end
                  if ((8'hb7))
                    begin
                      reg2846 <= forvar2827[(3'h5):(1'h1)];
                      reg2847 <= reg2586[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg2846 <= (-reg2694);
                      reg2847 <= reg2750;
                      reg2848 <= {(reg2682 && reg2773[(4'ha):(4'h9)])};
                    end
                  for (forvar2849 = (1'h0); (forvar2849 < (1'h1)); forvar2849 = (forvar2849 + (1'h1)))
                    begin
                      reg2850 <= {({(reg2657 * reg2620)} ?
                              $signed((+reg2597)) : (~^$unsigned(forvar2805)))};
                      reg2851 <= (!reg2593[(4'h8):(2'h3)]);
                      reg2852 <= reg2844[(1'h1):(1'h0)];
                    end
                end
              reg2853 <= $unsigned(forvar2833);
              for (forvar2854 = (1'h0); (forvar2854 < (1'h0)); forvar2854 = (forvar2854 + (1'h1)))
                begin
                  if (forvar2827[(4'ha):(3'h5)])
                    begin
                      reg2855 <= (~&(-$signed((reg2748 <<< reg2838))));
                      reg2856 <= reg2708;
                      reg2857 <= $unsigned($unsigned($unsigned($signed(reg2713))));
                      reg2858 <= {(8'hb9)};
                    end
                  else
                    begin
                      reg2855 <= reg2635[(2'h3):(1'h0)];
                      reg2856 <= ((~|$unsigned($signed((8'ha6)))) & ($unsigned((reg2780 < (8'h9c))) ?
                          reg2812[(1'h1):(1'h0)] : $unsigned(reg2694[(1'h1):(1'h1)])));
                    end
                  for (forvar2859 = (1'h0); (forvar2859 < (2'h3)); forvar2859 = (forvar2859 + (1'h1)))
                    begin
                      reg2860 <= ((~&(8'ha0)) << $signed($signed((reg2602 ?
                          forvar2822 : reg2697))));
                      reg2861 <= (~|forvar2796);
                      reg2862 <= forvar2803;
                      reg2863 <= {($signed($unsigned(wire2672)) >>> {(^~(8'ha1))})};
                    end
                  for (forvar2864 = (1'h0); (forvar2864 < (1'h0)); forvar2864 = (forvar2864 + (1'h1)))
                    begin
                      reg2865 <= (|reg2818[(3'h5):(2'h3)]);
                      reg2866 <= {forvar2852};
                      reg2867 <= $unsigned(reg2833[(4'h8):(3'h7)]);
                    end
                  reg2868 <= (-($signed(reg2827[(2'h2):(2'h2)]) * (^(~^forvar2840))));
                end
              reg2869 <= reg2704;
            end
        end
      for (forvar2880 = (1'h0); (forvar2880 < (1'h1)); forvar2880 = (forvar2880 + (1'h1)))
        begin
          reg2881 <= (^$signed(reg2722[(3'h4):(3'h4)]));
          for (forvar2882 = (1'h0); (forvar2882 < (2'h2)); forvar2882 = (forvar2882 + (1'h1)))
            begin
              for (forvar2883 = (1'h0); (forvar2883 < (1'h0)); forvar2883 = (forvar2883 + (1'h1)))
                begin
                  if (reg2696)
                    begin
                      reg2884 <= (~&($signed({reg2872}) ?
                          (|reg2855[(2'h2):(1'h0)]) : reg2766));
                      reg2885 <= (reg2856 || (^~((~^wire2585) ^~ {(8'ha1)})));
                    end
                  else
                    begin
                      reg2884 <= $unsigned($unsigned((&forvar2849[(2'h3):(2'h3)])));
                      reg2885 <= reg2838;
                      reg2886 <= (reg2660 <= (~^(8'hab)));
                      reg2887 <= (^~reg2695);
                    end
                end
              for (forvar2888 = (1'h0); (forvar2888 < (1'h1)); forvar2888 = (forvar2888 + (1'h1)))
                begin
                  for (forvar2889 = (1'h0); (forvar2889 < (2'h2)); forvar2889 = (forvar2889 + (1'h1)))
                    begin
                      reg2890 <= (reg2835 == (reg2874 ^~ wire2668));
                    end
                  if ($signed((((reg2693 >> reg2656) <<< (reg2805 ?
                          (8'hb1) : (8'had))) ?
                      (^{forvar2784}) : $signed((reg2842 - (8'ha2))))))
                    begin
                      reg2891 <= (forvar2796[(3'h5):(3'h4)] ?
                          (&$signed(reg2850[(1'h0):(1'h0)])) : ($signed((^~reg2807)) <<< reg2652[(4'h8):(2'h3)]));
                    end
                  else
                    begin
                      reg2891 <= {$unsigned(((reg2650 ?
                              reg2820 : reg2719) >> ((8'hb3) ?
                              reg2723 : reg2766)))};
                      reg2892 <= (8'hac);
                      reg2893 <= (reg2816 >> (($unsigned(reg2666) ^~ reg2831) ?
                          ((reg2862 ? reg2887 : reg2768) ?
                              (reg2702 >> reg2730) : $unsigned((8'hab))) : reg2849[(2'h2):(1'h1)]));
                    end
                  for (forvar2894 = (1'h0); (forvar2894 < (1'h1)); forvar2894 = (forvar2894 + (1'h1)))
                    begin
                      reg2895 <= $unsigned(reg2754);
                      reg2896 <= ((~(reg2865[(1'h1):(1'h1)] ?
                              {reg2664} : ((8'hb7) ? reg2799 : reg2874))) ?
                          reg2833[(3'h7):(2'h2)] : $unsigned(reg2618));
                      reg2897 <= $signed(reg2853);
                    end
                  if ($signed((reg2596[(2'h2):(2'h2)] * (reg2839 ?
                      {reg2830} : reg2785[(2'h3):(1'h1)]))))
                    begin
                      reg2898 <= forvar2862[(3'h6):(2'h3)];
                      reg2899 <= $unsigned((reg2627 >> $signed((|reg2644))));
                    end
                  else
                    begin
                      reg2898 <= $signed({(~(~&reg2696))});
                      reg2899 <= $signed($signed((|(8'ha8))));
                    end
                end
              for (forvar2900 = (1'h0); (forvar2900 < (1'h0)); forvar2900 = (forvar2900 + (1'h1)))
                begin
                  if ($unsigned(((|reg2615[(1'h1):(1'h1)]) && ((forvar2773 > forvar2870) ?
                      (reg2659 ^ reg2876) : (~^reg2840)))))
                    begin
                      reg2901 <= (reg2802[(4'h9):(1'h0)] ?
                          ($unsigned((~reg2701)) * $unsigned(reg2852[(3'h5):(1'h1)])) : $signed((8'ha6)));
                      reg2902 <= {($signed((|reg2857)) ?
                              $signed((reg2866 ?
                                  reg2726 : reg2678)) : reg2705[(1'h1):(1'h0)])};
                    end
                  else
                    begin
                      reg2901 <= $unsigned((~&($unsigned(reg2804) ?
                          $signed(forvar2854) : (+reg2857))));
                    end
                  for (forvar2903 = (1'h0); (forvar2903 < (2'h3)); forvar2903 = (forvar2903 + (1'h1)))
                    begin
                      reg2904 <= $signed($unsigned(($unsigned(reg2805) == $signed((8'hac)))));
                    end
                  for (forvar2905 = (1'h0); (forvar2905 < (1'h1)); forvar2905 = (forvar2905 + (1'h1)))
                    begin
                      reg2906 <= reg2722[(1'h0):(1'h0)];
                      reg2907 <= {forvar2803[(3'h4):(3'h4)]};
                      reg2908 <= reg2603[(2'h3):(2'h3)];
                      reg2909 <= (({(forvar2821 <<< reg2752)} || (((8'hb9) >>> reg2836) | forvar2865)) ?
                          reg2700 : ({(reg2658 < reg2613)} == ((!reg2790) ?
                              reg2598[(3'h6):(2'h2)] : (reg2845 * reg2739))));
                    end
                end
            end
          reg2910 <= $unsigned($unsigned($signed(((8'h9c) || reg2819))));
        end
      if ($unsigned((&(reg2606 ?
          (reg2659 ? reg2868 : reg2737) : reg2789[(3'h5):(1'h1)]))))
        begin
          if ((~&reg2717))
            begin
              reg2911 <= reg2609[(4'hc):(3'h5)];
            end
          else
            begin
              if (($unsigned(reg2615[(3'h6):(2'h3)]) >> $signed($signed((reg2712 ?
                  reg2886 : (8'had))))))
                begin
                  if (reg2718[(1'h1):(1'h0)])
                    begin
                      reg2911 <= (8'ha2);
                      reg2912 <= $unsigned({(~|(~|reg2632))});
                    end
                  else
                    begin
                      reg2911 <= reg2781[(1'h0):(1'h0)];
                    end
                  reg2913 <= forvar2837[(1'h1):(1'h0)];
                  if (({(~$unsigned(forvar2799))} ?
                      reg2586[(2'h3):(1'h1)] : (~^reg2838)))
                    begin
                      reg2914 <= $unsigned((({reg2737} ?
                              $unsigned(reg2818) : (~^reg2635)) ?
                          $unsigned(forvar2774) : (8'haa)));
                    end
                  else
                    begin
                      reg2914 <= $signed(reg2908);
                    end
                end
              else
                begin
                  if ((reg2724[(2'h2):(1'h0)] ?
                      $signed(reg2786[(2'h2):(1'h0)]) : ($unsigned($unsigned(reg2736)) ?
                          {reg2765[(3'h5):(2'h2)]} : (reg2623[(1'h0):(1'h0)] ^~ $unsigned(reg2600)))))
                    begin
                      reg2911 <= reg2849;
                      reg2912 <= (^(((reg2890 == reg2850) ?
                          {(8'h9c)} : reg2755[(4'hf):(4'h8)]) & reg2832[(4'hb):(3'h6)]));
                      reg2913 <= ($unsigned(reg2682[(2'h2):(1'h1)]) ?
                          $signed(((reg2808 ? reg2842 : reg2734) ?
                              forvar2820 : reg2757)) : {(&forvar2792)});
                      reg2914 <= {($signed($unsigned(reg2911)) ?
                              ((reg2852 ?
                                  forvar2889 : reg2861) >> forvar2777[(3'h7):(1'h1)]) : (-(reg2913 ?
                                  reg2819 : reg2762)))};
                    end
                  else
                    begin
                      reg2911 <= (forvar2903[(1'h1):(1'h0)] ?
                          (({reg2588} ?
                              (wire2673 ^~ forvar2782) : $unsigned((8'ha3))) ~^ ((forvar2782 != reg2907) || $unsigned(reg2715))) : {(~reg2807)});
                      reg2912 <= $signed(((~&(reg2904 ?
                          reg2594 : reg2808)) && {(&reg2704)}));
                    end
                end
              if (reg2737[(3'h4):(2'h3)])
                begin
                  reg2915 <= $unsigned((8'hab));
                end
              else
                begin
                  for (forvar2915 = (1'h0); (forvar2915 < (1'h1)); forvar2915 = (forvar2915 + (1'h1)))
                    begin
                      reg2916 <= ({$signed((reg2756 ?
                              reg2791 : reg2591))} & $unsigned(reg2813[(3'h4):(2'h3)]));
                      reg2917 <= (reg2625 ?
                          (8'h9f) : ($unsigned(reg2595[(4'ha):(1'h1)]) | $unsigned($unsigned(reg2765))));
                      reg2918 <= (~&(reg2771 ?
                          (^(forvar2807 == reg2901)) : ((!reg2658) <= {reg2639})));
                      reg2919 <= forvar2853[(1'h0):(1'h0)];
                    end
                  reg2920 <= $unsigned($signed(({reg2906} ?
                      (reg2798 << reg2800) : reg2692[(1'h1):(1'h1)])));
                  reg2921 <= reg2838;
                end
            end
          if (((~^(8'ha7)) ?
              (forvar2807[(1'h1):(1'h0)] <<< $unsigned($unsigned(wire2585))) : {$signed(((8'hb3) ?
                      reg2653 : reg2837))}))
            begin
              for (forvar2922 = (1'h0); (forvar2922 < (1'h1)); forvar2922 = (forvar2922 + (1'h1)))
                begin
                  for (forvar2923 = (1'h0); (forvar2923 < (2'h3)); forvar2923 = (forvar2923 + (1'h1)))
                    begin
                      reg2924 <= $signed(reg2617);
                      reg2925 <= reg2725;
                      reg2926 <= {{$signed(reg2759[(3'h5):(3'h5)])}};
                      reg2927 <= reg2692;
                    end
                  for (forvar2928 = (1'h0); (forvar2928 < (2'h3)); forvar2928 = (forvar2928 + (1'h1)))
                    begin
                      reg2929 <= ($unsigned({(reg2702 >>> (8'h9f))}) ?
                          $unsigned(reg2911[(2'h3):(2'h2)]) : (({reg2659} ?
                              reg2710 : {reg2843}) * reg2659[(3'h5):(2'h3)]));
                      reg2930 <= ((|$signed(reg2702)) ?
                          $signed($signed((reg2612 ?
                              reg2746 : reg2693))) : (~^({reg2588} ?
                              (reg2686 ?
                                  reg2778 : wire2585) : reg2821[(4'h8):(1'h0)])));
                      reg2931 <= (({$signed(reg2781)} && $signed(forvar2864)) ^ $signed(((reg2621 ?
                          reg2605 : reg2777) | reg2608)));
                    end
                  for (forvar2932 = (1'h0); (forvar2932 < (2'h3)); forvar2932 = (forvar2932 + (1'h1)))
                    begin
                      reg2933 <= ($unsigned(forvar2870) ?
                          (({reg2853} <= ((8'had) ?
                              reg2924 : reg2786)) >= (reg2730 ?
                              $signed(reg2639) : (reg2789 >> reg2843))) : $unsigned($unsigned(reg2859)));
                      reg2934 <= reg2655;
                      reg2935 <= ($unsigned($signed((^reg2893))) ?
                          $unsigned($signed({(8'had)})) : {((8'ha9) ?
                                  forvar2779 : $signed(forvar2787))});
                      reg2936 <= ($unsigned(reg2817) ?
                          $unsigned((forvar2803[(1'h0):(1'h0)] ?
                              (-(8'ha1)) : $unsigned(reg2712))) : ($signed(reg2705[(4'hd):(3'h7)]) ?
                              ((wire2668 && reg2589) < ((8'hb7) + reg2721)) : ((reg2877 ?
                                      forvar2779 : forvar2882) ?
                                  $unsigned((8'ha5)) : (reg2744 ?
                                      reg2660 : forvar2774))));
                    end
                end
              reg2937 <= $signed($unsigned(((forvar2840 ?
                  (8'hab) : forvar2812) > reg2593)));
            end
          else
            begin
              for (forvar2922 = (1'h0); (forvar2922 < (1'h1)); forvar2922 = (forvar2922 + (1'h1)))
                begin
                  for (forvar2923 = (1'h0); (forvar2923 < (1'h1)); forvar2923 = (forvar2923 + (1'h1)))
                    begin
                      reg2924 <= forvar2833[(3'h6):(3'h4)];
                      reg2925 <= reg2823[(1'h0):(1'h0)];
                      reg2926 <= (reg2805[(4'hb):(3'h6)] <<< reg2746[(2'h2):(1'h0)]);
                    end
                  for (forvar2927 = (1'h0); (forvar2927 < (2'h3)); forvar2927 = (forvar2927 + (1'h1)))
                    begin
                      reg2928 <= (8'hb0);
                      reg2929 <= (reg2837[(4'h9):(3'h4)] - (!((8'ha1) ?
                          (reg2871 | reg2935) : forvar2862)));
                      reg2930 <= $unsigned(wire2584);
                      reg2931 <= {((wire2672[(2'h3):(2'h3)] ^ (wire2585 ?
                              reg2813 : reg2866)) != (~|((8'hb3) != reg2667)))};
                    end
                  for (forvar2932 = (1'h0); (forvar2932 < (2'h3)); forvar2932 = (forvar2932 + (1'h1)))
                    begin
                      reg2933 <= (~|reg2698[(4'ha):(3'h4)]);
                    end
                  for (forvar2934 = (1'h0); (forvar2934 < (2'h3)); forvar2934 = (forvar2934 + (1'h1)))
                    begin
                      reg2935 <= forvar2915;
                    end
                end
              for (forvar2936 = (1'h0); (forvar2936 < (2'h2)); forvar2936 = (forvar2936 + (1'h1)))
                begin
                  if ($unsigned((~|(((8'haa) ? (8'h9f) : reg2935) ?
                      $signed(reg2652) : reg2840[(4'hc):(4'ha)]))))
                    begin
                      reg2937 <= $signed(($unsigned((8'hb9)) || (^{reg2849})));
                      reg2938 <= (8'ha8);
                    end
                  else
                    begin
                      reg2937 <= reg2833;
                    end
                  if (reg2805)
                    begin
                      reg2939 <= $signed((~|($unsigned(reg2592) ?
                          $signed(reg2746) : $unsigned((8'ha6)))));
                      reg2940 <= (($unsigned((+reg2629)) > reg2833) ?
                          $unsigned($unsigned(forvar2799)) : (^(reg2700 | forvar2936[(4'hb):(2'h2)])));
                    end
                  else
                    begin
                      reg2939 <= ((8'hba) ? {$signed((|reg2795))} : wire2669);
                      reg2940 <= $signed(reg2807);
                      reg2941 <= ((-(reg2738 ?
                              $unsigned(reg2818) : (^~reg2766))) ?
                          (($signed(reg2743) ? $signed(reg2656) : {reg2924}) ?
                              reg2627[(1'h1):(1'h1)] : $signed($signed(reg2748))) : $signed(forvar2807[(2'h2):(1'h1)]));
                      reg2942 <= (reg2734[(3'h7):(3'h7)] ?
                          (^~(forvar2800 ^~ (forvar2774 ?
                              reg2620 : reg2892))) : (reg2788 ?
                              reg2855 : $unsigned((~&forvar2894))));
                    end
                  for (forvar2943 = (1'h0); (forvar2943 < (2'h2)); forvar2943 = (forvar2943 + (1'h1)))
                    begin
                      reg2944 <= reg2619;
                      reg2945 <= (+(8'ha4));
                    end
                end
            end
          for (forvar2946 = (1'h0); (forvar2946 < (1'h0)); forvar2946 = (forvar2946 + (1'h1)))
            begin
              reg2947 <= (!(forvar2865[(2'h2):(1'h1)] != $signed((reg2848 ?
                  reg2765 : forvar2859))));
            end
        end
      else
        begin
          for (forvar2911 = (1'h0); (forvar2911 < (1'h1)); forvar2911 = (forvar2911 + (1'h1)))
            begin
              if (reg2702)
                begin
                  reg2912 <= $signed({$unsigned($signed(forvar2822))});
                  if (reg2830[(3'h6):(3'h4)])
                    begin
                      reg2913 <= reg2780;
                      reg2914 <= $signed($signed($signed(reg2916[(3'h5):(3'h4)])));
                      reg2915 <= reg2686;
                      reg2916 <= $signed(reg2691);
                    end
                  else
                    begin
                      reg2913 <= (|{reg2719});
                      reg2914 <= (!$signed(((reg2740 == (8'ha5)) <<< (8'hb7))));
                      reg2915 <= (reg2859[(1'h1):(1'h1)] ?
                          (|forvar2814[(3'h6):(3'h5)]) : (((^reg2858) == $unsigned(reg2824)) ^~ $unsigned($signed(forvar2800))));
                      reg2916 <= $unsigned(reg2642);
                    end
                  for (forvar2917 = (1'h0); (forvar2917 < (2'h2)); forvar2917 = (forvar2917 + (1'h1)))
                    begin
                      reg2918 <= {forvar2867};
                    end
                end
              else
                begin
                  if (({$signed($unsigned(reg2628))} ?
                      forvar2894 : ({reg2639[(1'h1):(1'h1)]} * $unsigned($signed((8'hb9))))))
                    begin
                      reg2912 <= reg2789[(3'h4):(3'h4)];
                      reg2913 <= (forvar2857[(2'h2):(1'h0)] ?
                          {(!(reg2716 - reg2639))} : $unsigned(((~|reg2625) ?
                              $signed(forvar2936) : $unsigned(reg2871))));
                      reg2914 <= (reg2631[(3'h5):(3'h5)] <<< $unsigned($signed(((8'ha4) == reg2815))));
                    end
                  else
                    begin
                      reg2912 <= (^{$unsigned((|reg2757))});
                      reg2913 <= reg2897;
                      reg2914 <= $signed((|$unsigned({forvar2905})));
                    end
                  if ((8'ha2))
                    begin
                      reg2915 <= $unsigned(forvar2799[(3'h5):(1'h1)]);
                      reg2916 <= reg2759[(4'hd):(4'ha)];
                      reg2917 <= (forvar2812 ?
                          (reg2700 ?
                              ($unsigned(reg2936) ?
                                  reg2645 : (reg2812 ?
                                      reg2928 : reg2878)) : reg2800[(1'h0):(1'h0)]) : forvar2936);
                    end
                  else
                    begin
                      reg2915 <= {{($unsigned((8'hb9)) ^ $unsigned(reg2651))}};
                      reg2916 <= {reg2934[(3'h4):(1'h0)]};
                      reg2917 <= (reg2749 ?
                          reg2819 : $unsigned({(forvar2903 ?
                                  reg2696 : reg2790)}));
                    end
                  for (forvar2918 = (1'h0); (forvar2918 < (1'h1)); forvar2918 = (forvar2918 + (1'h1)))
                    begin
                      reg2919 <= $signed(reg2646[(1'h0):(1'h0)]);
                      reg2920 <= wire2582;
                      reg2921 <= $signed(((8'hb9) ?
                          $unsigned($unsigned(reg2663)) : (~reg2745)));
                    end
                  if (((({reg2841} | reg2606[(2'h2):(1'h1)]) == ($signed(reg2606) - ((8'ha5) * reg2736))) ~^ $unsigned($unsigned($unsigned(reg2658)))))
                    begin
                      reg2922 <= {(~$unsigned((8'had)))};
                      reg2923 <= $signed((~^(+$signed(reg2871))));
                    end
                  else
                    begin
                      reg2922 <= $unsigned($unsigned(($unsigned(forvar2840) & $signed(reg2589))));
                      reg2923 <= {wire2581};
                    end
                end
              reg2924 <= (reg2719 || $unsigned($signed($signed(reg2818))));
              if ((-$unsigned($unsigned(reg2588[(3'h6):(1'h0)]))))
                begin
                  if (((&forvar2809[(3'h6):(1'h1)]) <= {reg2659[(3'h5):(1'h0)]}))
                    begin
                      reg2925 <= (reg2772[(1'h1):(1'h1)] ?
                          reg2915[(3'h7):(1'h0)] : $signed((~|(&wire2671))));
                      reg2926 <= (reg2666 <= {($unsigned(forvar2857) & reg2763)});
                      reg2927 <= {((forvar2779[(3'h7):(3'h4)] < {(8'h9d)}) ?
                              (~&$unsigned(reg2615)) : {(reg2920 + (8'ha1))})};
                      reg2928 <= $signed(reg2766[(3'h7):(2'h3)]);
                    end
                  else
                    begin
                      reg2925 <= $signed($signed((^(8'hae))));
                      reg2926 <= (~|$signed(reg2729[(3'h6):(3'h4)]));
                      reg2927 <= ($unsigned($unsigned(((8'hb9) ~^ forvar2922))) ?
                          {reg2858[(2'h3):(1'h0)]} : (wire2583[(2'h2):(2'h2)] + $signed((|forvar2787))));
                      reg2928 <= (forvar2792[(3'h4):(2'h2)] ?
                          $unsigned($unsigned($unsigned(reg2765))) : $signed($unsigned((forvar2946 >>> reg2659))));
                    end
                  for (forvar2929 = (1'h0); (forvar2929 < (1'h0)); forvar2929 = (forvar2929 + (1'h1)))
                    begin
                      reg2930 <= {reg2914};
                      reg2931 <= ({(~&{(8'h9f)})} <<< (({reg2754} ?
                          (forvar2818 ?
                              forvar2934 : forvar2813) : $unsigned(forvar2867)) == reg2650[(3'h5):(1'h1)]));
                      reg2932 <= reg2935[(2'h3):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar2925 = (1'h0); (forvar2925 < (1'h1)); forvar2925 = (forvar2925 + (1'h1)))
                    begin
                      reg2926 <= (&(wire2672 >>> reg2891[(2'h3):(1'h0)]));
                    end
                end
            end
          reg2933 <= (8'ha3);
          if ((forvar2888[(2'h3):(2'h2)] * $unsigned(((+wire2583) ?
              reg2861 : $unsigned(reg2907)))))
            begin
              for (forvar2934 = (1'h0); (forvar2934 < (2'h3)); forvar2934 = (forvar2934 + (1'h1)))
                begin
                  for (forvar2935 = (1'h0); (forvar2935 < (1'h0)); forvar2935 = (forvar2935 + (1'h1)))
                    begin
                      reg2936 <= (reg2937[(2'h2):(1'h0)] ?
                          {forvar2813} : (reg2594 ?
                              $unsigned($signed((8'h9e))) : ((reg2806 >> wire2580) ?
                                  (forvar2889 ?
                                      reg2742 : reg2629) : forvar2854)));
                      reg2937 <= (+reg2734[(1'h0):(1'h0)]);
                    end
                  if ((~|reg2722[(1'h0):(1'h0)]))
                    begin
                      reg2938 <= ($unsigned($signed((reg2654 >>> reg2721))) ?
                          ((reg2719[(2'h2):(2'h2)] ~^ (forvar2803 >> forvar2813)) ^ (8'ha2)) : $signed(reg2611));
                      reg2939 <= reg2761;
                    end
                  else
                    begin
                      reg2938 <= $signed(forvar2883);
                      reg2939 <= ((+((!forvar2946) >= $signed(reg2715))) ?
                          $unsigned($signed(forvar2864)) : reg2926[(3'h5):(1'h1)]);
                      reg2940 <= reg2627[(1'h0):(1'h0)];
                    end
                  for (forvar2941 = (1'h0); (forvar2941 < (2'h3)); forvar2941 = (forvar2941 + (1'h1)))
                    begin
                      reg2942 <= (~&$signed(forvar2905));
                      reg2943 <= reg2706[(1'h1):(1'h1)];
                      reg2944 <= reg2758[(3'h4):(2'h2)];
                    end
                  for (forvar2945 = (1'h0); (forvar2945 < (1'h0)); forvar2945 = (forvar2945 + (1'h1)))
                    begin
                      reg2946 <= (~^(~|(8'ha7)));
                    end
                end
            end
          else
            begin
              reg2934 <= (-(reg2770[(1'h1):(1'h0)] != (^$unsigned(reg2831))));
              for (forvar2935 = (1'h0); (forvar2935 < (1'h1)); forvar2935 = (forvar2935 + (1'h1)))
                begin
                  if (reg2798[(3'h7):(2'h2)])
                    begin
                      reg2936 <= $signed(reg2629[(1'h0):(1'h0)]);
                      reg2937 <= $signed((~$signed((~^reg2921))));
                    end
                  else
                    begin
                      reg2936 <= (8'haf);
                      reg2937 <= $signed(((~reg2662) ?
                          $signed($unsigned(reg2939)) : $signed($unsigned(reg2931))));
                    end
                  for (forvar2938 = (1'h0); (forvar2938 < (2'h2)); forvar2938 = (forvar2938 + (1'h1)))
                    begin
                      reg2939 <= reg2731;
                      reg2940 <= reg2838[(4'h8):(2'h2)];
                      reg2941 <= $signed(reg2639);
                    end
                end
              for (forvar2942 = (1'h0); (forvar2942 < (2'h2)); forvar2942 = (forvar2942 + (1'h1)))
                begin
                  if ((+{reg2742[(1'h1):(1'h1)]}))
                    begin
                      reg2943 <= reg2874[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg2943 <= reg2656;
                    end
                end
              if ((&((8'hac) > $signed(reg2822[(1'h1):(1'h0)]))))
                begin
                  for (forvar2944 = (1'h0); (forvar2944 < (1'h0)); forvar2944 = (forvar2944 + (1'h1)))
                    begin
                      reg2945 <= $unsigned({reg2652[(3'h7):(2'h2)]});
                      reg2946 <= reg2918;
                      reg2947 <= $signed(reg2890[(2'h3):(1'h1)]);
                    end
                  for (forvar2948 = (1'h0); (forvar2948 < (2'h3)); forvar2948 = (forvar2948 + (1'h1)))
                    begin
                      reg2949 <= reg2907;
                      reg2950 <= $signed((|$signed((^(8'h9f)))));
                      reg2951 <= (reg2818[(4'ha):(3'h6)] || wire2668);
                      reg2952 <= (8'ha1);
                    end
                end
              else
                begin
                  for (forvar2944 = (1'h0); (forvar2944 < (1'h0)); forvar2944 = (forvar2944 + (1'h1)))
                    begin
                      reg2945 <= $signed((reg2791[(4'ha):(4'ha)] ?
                          reg2858 : ({wire2673} ? reg2869 : (+reg2587))));
                      reg2946 <= $signed(reg2683);
                      reg2947 <= ({(reg2904[(1'h1):(1'h0)] ?
                              (reg2652 ?
                                  (8'ha3) : reg2826) : reg2630)} >>> $unsigned($unsigned((~|reg2751))));
                      reg2948 <= reg2779[(1'h0):(1'h0)];
                    end
                end
            end
          for (forvar2953 = (1'h0); (forvar2953 < (2'h3)); forvar2953 = (forvar2953 + (1'h1)))
            begin
              reg2954 <= reg2911[(3'h4):(2'h3)];
              if ($unsigned((&forvar2943[(1'h0):(1'h0)])))
                begin
                  reg2955 <= $unsigned((!reg2811[(4'ha):(1'h0)]));
                  reg2956 <= $unsigned((($unsigned(reg2854) ?
                      ((8'hb8) <= reg2831) : (reg2775 || wire2580)) == $unsigned((8'ha6))));
                  if ($unsigned(($signed((reg2708 ? forvar2857 : (8'hab))) ?
                      reg2805 : ((forvar2932 - reg2779) | $unsigned(wire2668)))))
                    begin
                      reg2957 <= $unsigned(((forvar2877 ?
                          $signed(reg2684) : (reg2909 ?
                              reg2777 : reg2616)) == reg2709));
                    end
                  else
                    begin
                      reg2957 <= (wire2672[(1'h0):(1'h0)] >> $unsigned(forvar2833));
                      reg2958 <= (reg2897[(4'h9):(1'h1)] ?
                          $signed(((forvar2932 << (8'hba)) & wire2583)) : ($signed((^~reg2922)) ?
                              reg2682 : ((reg2636 ? reg2857 : (8'ha6)) ?
                                  (~^reg2631) : (~|reg2737))));
                      reg2959 <= wire2671[(2'h2):(2'h2)];
                      reg2960 <= (|$signed($unsigned(reg2708)));
                    end
                  if ($signed(reg2929[(2'h3):(2'h3)]))
                    begin
                      reg2961 <= $unsigned((~^reg2726));
                      reg2962 <= ($unsigned({(reg2722 - (8'hb4))}) ?
                          ($signed((reg2605 ?
                              forvar2793 : (8'hac))) <<< reg2956) : reg2854[(4'h9):(3'h6)]);
                    end
                  else
                    begin
                      reg2961 <= ($signed(reg2756) ?
                          reg2588 : $unsigned((|$signed(forvar2834))));
                      reg2962 <= $signed(forvar2905[(1'h0):(1'h0)]);
                      reg2963 <= ($unsigned($signed(((8'ha4) ?
                          reg2911 : (8'ha1)))) * $unsigned((|(reg2842 ?
                          forvar2799 : reg2619))));
                    end
                end
              else
                begin
                  if ($signed($unsigned(({forvar2888} ?
                      $signed(reg2621) : reg2696[(1'h0):(1'h0)]))))
                    begin
                      reg2955 <= ((^~$unsigned((reg2820 >= reg2731))) + $unsigned($unsigned($signed(reg2886))));
                      reg2956 <= $signed((reg2738 && $signed({reg2657})));
                      reg2957 <= (($signed(reg2621) ?
                          ($unsigned(reg2850) ?
                              reg2850 : reg2695[(1'h0):(1'h0)]) : ($signed(reg2731) ?
                              $unsigned(forvar2944) : $signed(reg2774))) >> $signed(reg2722[(2'h2):(1'h0)]));
                      reg2958 <= $unsigned(reg2956);
                    end
                  else
                    begin
                      reg2955 <= ($signed($unsigned(reg2737)) ?
                          (((reg2815 >>> reg2699) ?
                                  (reg2814 <<< reg2777) : (|reg2963)) ?
                              $unsigned((forvar2864 ?
                                  reg2712 : forvar2867)) : reg2921) : ($signed($unsigned(forvar2945)) ?
                              (|((8'hb6) > reg2635)) : (~(reg2841 ?
                                  reg2871 : forvar2790))));
                      reg2956 <= reg2599;
                      reg2957 <= (8'hb7);
                      reg2958 <= {($signed($unsigned(reg2659)) ?
                              ((reg2684 ? forvar2857 : (8'h9c)) ?
                                  reg2886[(4'he):(4'hb)] : $unsigned(wire2580)) : forvar2859)};
                    end
                end
            end
        end
      for (forvar2964 = (1'h0); (forvar2964 < (1'h1)); forvar2964 = (forvar2964 + (1'h1)))
        begin
          if (reg2797)
            begin
              if ($signed(reg2621[(2'h2):(1'h1)]))
                begin
                  for (forvar2965 = (1'h0); (forvar2965 < (2'h3)); forvar2965 = (forvar2965 + (1'h1)))
                    begin
                      reg2966 <= reg2752;
                      reg2967 <= $signed((^(reg2650 ? {(8'ha9)} : reg2742)));
                    end
                  if (($signed($unsigned((~&reg2912))) ?
                      $signed($unsigned((wire2671 <<< reg2823))) : (~|($unsigned((8'hb7)) >> (reg2748 || reg2633)))))
                    begin
                      reg2968 <= (($unsigned($signed(reg2828)) ?
                              (8'hb0) : (reg2924 && (forvar2818 ?
                                  reg2768 : reg2588))) ?
                          reg2926[(2'h3):(2'h2)] : (((reg2785 ?
                                  forvar2809 : reg2780) + reg2943) ?
                              reg2930 : (~((8'hb3) ^~ reg2885))));
                    end
                  else
                    begin
                      reg2968 <= (^~{(~^(~^forvar2774))});
                      reg2969 <= ($signed(reg2641[(3'h5):(2'h3)]) ?
                          ((~|(~&reg2615)) ?
                              $signed((8'haa)) : $unsigned(reg2931)) : $unsigned(reg2590));
                    end
                end
              else
                begin
                  for (forvar2965 = (1'h0); (forvar2965 < (2'h2)); forvar2965 = (forvar2965 + (1'h1)))
                    begin
                      reg2966 <= reg2702;
                      reg2967 <= ((((reg2837 ? forvar2932 : wire2668) ?
                              $unsigned(reg2918) : (~(8'had))) >>> $signed(reg2863)) ?
                          (|(^(-reg2736))) : {$signed((reg2713 >> reg2890))});
                      reg2968 <= reg2969[(2'h2):(2'h2)];
                      reg2969 <= $signed(reg2837[(1'h0):(1'h0)]);
                    end
                end
              reg2970 <= (((&reg2955) ^ $unsigned(reg2873)) ?
                  reg2901 : (wire2583 ?
                      $unsigned($unsigned(reg2761)) : reg2879[(1'h1):(1'h0)]));
            end
          else
            begin
              reg2965 <= $unsigned(reg2855);
              if ((reg2893 ^~ {{(reg2605 >> reg2963)}}))
                begin
                  reg2966 <= (~^{reg2759[(2'h2):(2'h2)]});
                  reg2967 <= ($unsigned(((forvar2840 ? reg2733 : reg2706) ?
                      (+reg2836) : reg2627)) && (~^(&$unsigned((8'ha2)))));
                  for (forvar2968 = (1'h0); (forvar2968 < (1'h1)); forvar2968 = (forvar2968 + (1'h1)))
                    begin
                      reg2969 <= reg2797[(3'h6):(3'h6)];
                      reg2970 <= (+$signed((!reg2801[(4'hb):(3'h6)])));
                      reg2971 <= (((|reg2658) ^~ forvar2945) || reg2609[(4'he):(1'h1)]);
                      reg2972 <= $signed(($signed(reg2815[(3'h6):(3'h5)]) >> {((8'h9c) ?
                              forvar2782 : (8'hba))}));
                    end
                end
              else
                begin
                  for (forvar2966 = (1'h0); (forvar2966 < (1'h1)); forvar2966 = (forvar2966 + (1'h1)))
                    begin
                      reg2967 <= forvar2900;
                      reg2968 <= reg2762[(3'h5):(1'h0)];
                    end
                  reg2969 <= {(!(^~$signed(forvar2800)))};
                end
              reg2973 <= ($unsigned($unsigned(reg2614[(4'hd):(2'h3)])) ?
                  reg2784 : $signed((~&$signed(wire2669))));
            end
          if ($signed($unsigned((~|(^~reg2747)))))
            begin
              for (forvar2974 = (1'h0); (forvar2974 < (2'h3)); forvar2974 = (forvar2974 + (1'h1)))
                begin
                  reg2975 <= (^~(-(~&(reg2607 ? reg2648 : reg2942))));
                  for (forvar2976 = (1'h0); (forvar2976 < (2'h3)); forvar2976 = (forvar2976 + (1'h1)))
                    begin
                      reg2977 <= (|({$unsigned((8'hb1))} ?
                          ($unsigned(reg2733) * $unsigned(reg2929)) : $unsigned($signed((8'hb2)))));
                      reg2978 <= reg2608[(4'he):(2'h3)];
                    end
                  for (forvar2979 = (1'h0); (forvar2979 < (2'h2)); forvar2979 = (forvar2979 + (1'h1)))
                    begin
                      reg2980 <= (8'ha5);
                      reg2981 <= reg2598;
                      reg2982 <= $signed(forvar2803[(1'h1):(1'h0)]);
                    end
                  if ($unsigned((reg2850 ?
                      reg2943[(3'h5):(2'h2)] : reg2966[(1'h1):(1'h1)])))
                    begin
                      reg2983 <= $unsigned((!reg2921[(3'h6):(3'h5)]));
                      reg2984 <= (!(((reg2887 ?
                              reg2906 : reg2708) >> (~&forvar2782)) ?
                          $unsigned($signed(reg2726)) : (|reg2634)));
                      reg2985 <= (reg2934[(2'h3):(1'h0)] > $unsigned(($unsigned(reg2817) ?
                          $signed(reg2733) : (reg2805 ? reg2867 : reg2977))));
                      reg2986 <= (-reg2620[(4'h9):(1'h0)]);
                    end
                  else
                    begin
                      reg2983 <= $unsigned(forvar2782);
                    end
                end
              if (reg2755[(5'h10):(4'ha)])
                begin
                  for (forvar2987 = (1'h0); (forvar2987 < (1'h0)); forvar2987 = (forvar2987 + (1'h1)))
                    begin
                      reg2988 <= reg2980;
                      reg2989 <= (reg2683 ?
                          (^~($unsigned((8'hb5)) ?
                              forvar2807[(1'h0):(1'h0)] : $unsigned((8'ha0)))) : (^~reg2686));
                      reg2990 <= $unsigned(reg2733);
                    end
                  if (((!$unsigned(forvar2862)) >> $unsigned(($unsigned(reg2984) | reg2588))))
                    begin
                      reg2991 <= {$signed(reg2852[(4'ha):(1'h1)])};
                      reg2992 <= $unsigned((({reg2701} ~^ (reg2968 ?
                          reg2968 : forvar2774)) ~^ (!$signed((8'ha8)))));
                    end
                  else
                    begin
                      reg2991 <= $signed($signed({$unsigned(reg2783)}));
                    end
                end
              else
                begin
                  for (forvar2987 = (1'h0); (forvar2987 < (1'h0)); forvar2987 = (forvar2987 + (1'h1)))
                    begin
                      reg2988 <= $unsigned($signed($signed((reg2857 && reg2630))));
                      reg2989 <= ($signed($unsigned((~|forvar2905))) ?
                          $unsigned(reg2983) : {(~&{(8'ha3)})});
                      reg2990 <= $unsigned((((reg2724 >= forvar2905) ?
                          reg2715[(4'hd):(3'h6)] : reg2628) < ($unsigned(reg2896) ?
                          reg2963[(4'h8):(3'h6)] : reg2919[(2'h3):(1'h1)])));
                    end
                  if ($unsigned(({reg2860} ?
                      ((^~reg2817) ~^ reg2781[(2'h3):(1'h1)]) : $unsigned((forvar2847 ?
                          forvar2834 : reg2943)))))
                    begin
                      reg2991 <= {$unsigned({(|reg2738)})};
                      reg2992 <= reg2699;
                    end
                  else
                    begin
                      reg2991 <= (reg2590 >> ($unsigned((-reg2985)) - {(forvar2900 == reg2713)}));
                      reg2992 <= (^(((reg2710 - forvar2944) || (~&(8'hb7))) ?
                          ({reg2909} ?
                              reg2615 : (forvar2818 ?
                                  (8'hb1) : reg2613)) : (reg2828 ?
                              (~^reg2781) : (reg2618 <= reg2825))));
                      reg2993 <= ((&$signed((8'ha6))) == $unsigned({(reg2873 > reg2824)}));
                      reg2994 <= (reg2629 || $signed((^(forvar2803 || reg2924))));
                    end
                end
              for (forvar2995 = (1'h0); (forvar2995 < (1'h1)); forvar2995 = (forvar2995 + (1'h1)))
                begin
                  for (forvar2996 = (1'h0); (forvar2996 < (1'h1)); forvar2996 = (forvar2996 + (1'h1)))
                    begin
                      reg2997 <= ({reg2738[(3'h6):(2'h3)]} && (^~forvar2936));
                      reg2998 <= ($unsigned(reg2620) | ($signed((reg2924 ?
                          reg2925 : reg2743)) >>> reg2839));
                      reg2999 <= $signed({(!(~reg2845))});
                    end
                  for (forvar3000 = (1'h0); (forvar3000 < (2'h3)); forvar3000 = (forvar3000 + (1'h1)))
                    begin
                      reg3001 <= ({(((8'hb7) * (8'hb6)) * {reg2951})} ?
                          reg2724[(4'ha):(1'h0)] : reg2712[(3'h5):(2'h2)]);
                    end
                  if ((-({$unsigned(reg2607)} * forvar2820[(4'hb):(2'h2)])))
                    begin
                      reg3002 <= $signed(reg2998);
                      reg3003 <= {$signed((~|{reg2918}))};
                      reg3004 <= $unsigned((^~$unsigned((reg2715 <<< reg2835))));
                    end
                  else
                    begin
                      reg3002 <= reg2950[(4'ha):(2'h3)];
                      reg3003 <= reg2879;
                      reg3004 <= (!forvar2925[(1'h0):(1'h0)]);
                      reg3005 <= $unsigned($signed($signed((|forvar2889))));
                    end
                end
              for (forvar3006 = (1'h0); (forvar3006 < (1'h1)); forvar3006 = (forvar3006 + (1'h1)))
                begin
                  reg3007 <= $signed($unsigned(((reg2718 ? reg2642 : (8'hb2)) ?
                      reg2809 : (reg2983 - reg2745))));
                  if (forvar2888)
                    begin
                      reg3008 <= (^($unsigned(reg2633[(3'h5):(3'h4)]) ?
                          (^$signed(reg2614)) : forvar2821[(2'h3):(2'h3)]));
                    end
                  else
                    begin
                      reg3008 <= ((($unsigned(reg2653) << reg2881) ^~ (reg2715[(1'h1):(1'h1)] ?
                              reg2799[(1'h0):(1'h0)] : (^~forvar2809))) ?
                          reg2636[(3'h5):(2'h2)] : reg2778);
                      reg3009 <= (~|{(reg2765 - (~(8'ha9)))});
                      reg3010 <= (^~reg2826[(3'h6):(1'h1)]);
                    end
                end
            end
          else
            begin
              for (forvar2974 = (1'h0); (forvar2974 < (2'h3)); forvar2974 = (forvar2974 + (1'h1)))
                begin
                  for (forvar2975 = (1'h0); (forvar2975 < (1'h0)); forvar2975 = (forvar2975 + (1'h1)))
                    begin
                      reg2976 <= (reg2625 != forvar2857);
                      reg2977 <= $signed(reg2746);
                      reg2978 <= forvar2816;
                    end
                  for (forvar2979 = (1'h0); (forvar2979 < (2'h3)); forvar2979 = (forvar2979 + (1'h1)))
                    begin
                      reg2980 <= {($unsigned({reg2704}) ?
                              ((reg2753 > reg2775) & {reg2860}) : $unsigned($unsigned(reg2839)))};
                      reg2981 <= reg2738;
                      reg2982 <= $unsigned(($signed({reg2786}) ?
                          reg2809[(2'h3):(1'h0)] : reg2983));
                    end
                  if ($signed($unsigned({$unsigned(reg2969)})))
                    begin
                      reg2983 <= (({(forvar2790 ?
                                  reg2927 : forvar2816)} <= reg2988) ?
                          $signed({(reg2965 * reg2908)}) : $signed(forvar2800[(3'h7):(2'h3)]));
                      reg2984 <= ((reg2788[(1'h0):(1'h0)] > {{reg2841}}) ^ $unsigned(($signed(reg2716) ?
                          (wire2584 | reg2921) : $signed(reg2634))));
                    end
                  else
                    begin
                      reg2983 <= $unsigned(forvar2822);
                      reg2984 <= ((reg2641[(2'h3):(1'h0)] ?
                              forvar2905[(1'h0):(1'h0)] : (^(forvar2875 - reg2786))) ?
                          reg2899 : {$signed(reg2930[(3'h7):(3'h4)])});
                    end
                  if ((~^(!$signed((+(8'hb8))))))
                    begin
                      reg2985 <= $signed(((forvar2816 ?
                              (^~reg2813) : (reg2733 ? reg2984 : reg2975)) ?
                          $unsigned(forvar2800[(3'h7):(1'h1)]) : {(reg2621 > reg2982)}));
                      reg2986 <= ($unsigned((((8'ha7) && (8'hb6)) <<< ((8'hac) ?
                          (8'hb6) : reg2898))) * {$signed((reg2830 > (8'hb0)))});
                      reg2987 <= $unsigned(reg2617[(4'h8):(3'h5)]);
                    end
                  else
                    begin
                      reg2985 <= reg2663;
                    end
                end
              for (forvar2988 = (1'h0); (forvar2988 < (2'h3)); forvar2988 = (forvar2988 + (1'h1)))
                begin
                  for (forvar2989 = (1'h0); (forvar2989 < (2'h3)); forvar2989 = (forvar2989 + (1'h1)))
                    begin
                      reg2990 <= forvar2857[(2'h2):(1'h0)];
                    end
                  if ((+reg2926[(1'h1):(1'h1)]))
                    begin
                      reg2991 <= reg2879[(1'h0):(1'h0)];
                      reg2992 <= (^~$signed($signed($signed(reg2602))));
                    end
                  else
                    begin
                      reg2991 <= $signed($signed(($unsigned(reg2596) + reg2713[(2'h3):(2'h2)])));
                      reg2992 <= $signed((8'hab));
                      reg2993 <= $unsigned((($unsigned(forvar2792) ?
                          {reg2615} : {(8'hb5)}) == forvar2966));
                    end
                  for (forvar2994 = (1'h0); (forvar2994 < (2'h2)); forvar2994 = (forvar2994 + (1'h1)))
                    begin
                      reg2995 <= (~|forvar2925);
                      reg2996 <= (reg2754[(4'hd):(2'h3)] > ($signed((reg2757 ?
                              reg2711 : forvar2929)) ?
                          (forvar2953 != (reg2815 << reg3009)) : $signed($unsigned(reg2815))));
                      reg2997 <= (8'hb1);
                    end
                end
            end
          if (reg2806)
            begin
              for (forvar3011 = (1'h0); (forvar3011 < (2'h2)); forvar3011 = (forvar3011 + (1'h1)))
                begin
                  for (forvar3012 = (1'h0); (forvar3012 < (1'h1)); forvar3012 = (forvar3012 + (1'h1)))
                    begin
                      reg3013 <= (((8'hb4) ?
                          (~reg2927) : $unsigned(reg2644)) << forvar2946);
                    end
                  reg3014 <= (^~$unsigned(reg2790));
                  reg3015 <= forvar2807[(2'h2):(1'h0)];
                  reg3016 <= ((^$signed((reg2975 ? (8'hb9) : forvar3006))) ?
                      ((&$signed(forvar2814)) - forvar2935) : reg2768);
                end
              for (forvar3017 = (1'h0); (forvar3017 < (2'h2)); forvar3017 = (forvar3017 + (1'h1)))
                begin
                  if ($unsigned(((&(reg2611 ?
                      reg2597 : forvar2782)) && (+(reg2980 ?
                      reg2745 : reg2738)))))
                    begin
                      reg3018 <= $unsigned((-reg2703[(3'h5):(3'h5)]));
                      reg3019 <= reg2752;
                    end
                  else
                    begin
                      reg3018 <= (8'ha2);
                    end
                  if ({(reg2627 * (8'h9c))})
                    begin
                      reg3020 <= ($unsigned($signed(reg3003[(1'h0):(1'h0)])) - (~|(forvar2789 ?
                          (|reg2973) : $signed(reg2779))));
                      reg3021 <= $unsigned(($unsigned(reg2682[(3'h6):(2'h3)]) ~^ (&(reg2792 >= reg2839))));
                      reg3022 <= (reg2909[(1'h1):(1'h1)] ?
                          (8'h9c) : (~|reg2981));
                      reg3023 <= $signed(($unsigned(reg2747) * $signed(reg2654)));
                    end
                  else
                    begin
                      reg3020 <= {(((reg3022 ~^ wire2670) <= $unsigned(reg2708)) >= $signed((~&reg2684)))};
                      reg3021 <= {(8'hb0)};
                      reg3022 <= $unsigned(reg2992);
                    end
                  reg3024 <= (+({{forvar2883}} ? (+reg3005) : {(~reg2682)}));
                  for (forvar3025 = (1'h0); (forvar3025 < (1'h0)); forvar3025 = (forvar3025 + (1'h1)))
                    begin
                      reg3026 <= (+(8'hb4));
                      reg3027 <= ($unsigned($signed(forvar2814)) ^~ (((|reg2876) ^ (reg2943 > reg2982)) ?
                          reg2972[(3'h4):(2'h3)] : (|reg2899[(4'ha):(3'h7)])));
                      reg3028 <= (~|$unsigned((^(reg2923 == reg2801))));
                      reg3029 <= $signed(wire2672);
                    end
                end
              if (reg2831)
                begin
                  for (forvar3030 = (1'h0); (forvar3030 < (2'h2)); forvar3030 = (forvar3030 + (1'h1)))
                    begin
                      reg3031 <= $signed(reg2597[(3'h5):(1'h1)]);
                      reg3032 <= $unsigned({reg2798});
                      reg3033 <= reg2599;
                      reg3034 <= forvar2923[(4'ha):(3'h6)];
                    end
                end
              else
                begin
                  if (reg2791)
                    begin
                      reg3030 <= reg2621;
                      reg3031 <= reg2791;
                      reg3032 <= $signed((~|forvar2867));
                      reg3033 <= $unsigned({$unsigned((~^(8'hb3)))});
                    end
                  else
                    begin
                      reg3030 <= forvar2968[(2'h3):(2'h3)];
                      reg3031 <= reg2725[(4'ha):(4'ha)];
                    end
                  for (forvar3034 = (1'h0); (forvar3034 < (2'h3)); forvar3034 = (forvar3034 + (1'h1)))
                    begin
                      reg3035 <= $signed(($signed(reg2730) & {(reg2904 >= reg2794)}));
                      reg3036 <= $unsigned(reg2973[(3'h5):(2'h2)]);
                      reg3037 <= reg2803[(4'hc):(2'h2)];
                    end
                end
            end
          else
            begin
              for (forvar3011 = (1'h0); (forvar3011 < (2'h3)); forvar3011 = (forvar3011 + (1'h1)))
                begin
                  for (forvar3012 = (1'h0); (forvar3012 < (2'h3)); forvar3012 = (forvar3012 + (1'h1)))
                    begin
                      reg3013 <= (reg2620 | reg2707[(4'hd):(2'h2)]);
                    end
                  reg3014 <= $signed($signed((-forvar2942)));
                end
              for (forvar3015 = (1'h0); (forvar3015 < (1'h0)); forvar3015 = (forvar3015 + (1'h1)))
                begin
                  for (forvar3016 = (1'h0); (forvar3016 < (2'h3)); forvar3016 = (forvar3016 + (1'h1)))
                    begin
                      reg3017 <= ((+(!reg2892[(3'h5):(3'h5)])) ?
                          (8'hab) : forvar2841[(3'h5):(2'h3)]);
                      reg3018 <= reg2691[(4'h8):(3'h7)];
                      reg3019 <= forvar2852[(1'h1):(1'h0)];
                      reg3020 <= (|(8'ha5));
                    end
                end
              for (forvar3021 = (1'h0); (forvar3021 < (1'h1)); forvar3021 = (forvar3021 + (1'h1)))
                begin
                  if ($unsigned($signed((reg2839 == {reg2830}))))
                    begin
                      reg3022 <= (^reg2586[(1'h0):(1'h0)]);
                      reg3023 <= $signed($signed(((reg2907 >>> reg2994) ?
                          {forvar2974} : (reg2935 ^ reg2872))));
                      reg3024 <= forvar2974[(3'h7):(3'h5)];
                      reg3025 <= ($signed($signed(forvar2948)) ?
                          reg2824[(2'h3):(2'h2)] : ($signed((reg2914 ~^ reg2720)) ?
                              ($signed(reg2743) ?
                                  $signed(reg2708) : (reg2881 ?
                                      (8'hae) : forvar2841)) : reg2937[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg3022 <= $unsigned(($unsigned((reg2784 ~^ reg2759)) <= ($signed(forvar2966) ?
                          $signed(reg2990) : forvar2870)));
                      reg3023 <= (&reg2851);
                      reg3024 <= reg2661;
                    end
                  for (forvar3026 = (1'h0); (forvar3026 < (1'h0)); forvar3026 = (forvar3026 + (1'h1)))
                    begin
                      reg3027 <= reg2586[(1'h0):(1'h0)];
                      reg3028 <= (($unsigned($signed(reg2622)) <= {$signed(reg2908)}) ^~ forvar2833);
                      reg3029 <= reg2837;
                    end
                  for (forvar3030 = (1'h0); (forvar3030 < (2'h3)); forvar3030 = (forvar3030 + (1'h1)))
                    begin
                      reg3031 <= (((&(-reg2944)) ?
                              reg2967 : (^~(reg2971 ? reg2663 : reg2763))) ?
                          (|((~^(8'ha1)) ?
                              {reg2629} : $unsigned(reg2621))) : $signed(reg2871));
                      reg3032 <= ((~$signed($signed(reg2885))) ?
                          (8'ha9) : (8'ha8));
                      reg3033 <= {($signed(reg2869[(3'h6):(1'h0)]) ?
                              $unsigned(reg2654) : ({reg2851} ?
                                  (reg2782 ?
                                      forvar3034 : forvar2840) : $unsigned(reg2833)))};
                      reg3034 <= $signed(forvar2820);
                    end
                end
              reg3035 <= $unsigned((reg2965 ? (8'ha3) : $signed(forvar2923)));
            end
        end
    end
  assign wire3038 = (((^~$signed(reg2798)) ?
                            {(~reg2930)} : $signed(reg2830[(3'h7):(3'h5)])) ?
                        $signed(reg2762) : reg2749);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2393
#(parameter param2501 = (({((8'hae) ? (8'haf) : (8'hb8))} | (8'h9c)) ? (~&(!((8'ha9) ? (8'ha3) : (8'ha6)))) : ({((8'ha2) ~^ (8'h9d))} ? (^((8'ha1) & (8'hb3))) : (((8'hb1) ? (8'haf) : (8'hb6)) >>> ((8'ha3) <<< (8'ha2))))))
(y, clk, wire2398, wire2397, wire2396, wire2395, wire2394);
  output wire [(32'h48d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire2398;
  input wire signed [(4'hb):(1'h0)] wire2397;
  input wire signed [(4'ha):(1'h0)] wire2396;
  input wire [(5'h10):(1'h0)] wire2395;
  input wire signed [(4'h9):(1'h0)] wire2394;
  wire signed [(3'h7):(1'h0)] wire2500;
  wire signed [(3'h7):(1'h0)] wire2499;
  wire [(2'h2):(1'h0)] wire2498;
  wire signed [(5'h10):(1'h0)] wire2497;
  wire [(3'h6):(1'h0)] wire2496;
  reg [(3'h7):(1'h0)] reg2495 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2494 = (1'h0);
  reg [(3'h7):(1'h0)] reg2493 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2492 = (1'h0);
  reg [(4'hb):(1'h0)] reg2487 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2491 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2490 = (1'h0);
  reg [(4'ha):(1'h0)] reg2489 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2488 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2477 = (1'h0);
  reg [(4'ha):(1'h0)] reg2485 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2484 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2483 = (1'h0);
  reg [(4'hc):(1'h0)] reg2482 = (1'h0);
  reg [(4'hb):(1'h0)] reg2481 = (1'h0);
  reg [(4'he):(1'h0)] reg2480 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2479 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2478 = (1'h0);
  reg [(2'h3):(1'h0)] reg2476 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2475 = (1'h0);
  reg [(4'hb):(1'h0)] reg2473 = (1'h0);
  reg [(5'h10):(1'h0)] reg2472 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2471 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2470 = (1'h0);
  reg [(4'h9):(1'h0)] reg2467 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2465 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2464 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2463 = (1'h0);
  reg [(4'h9):(1'h0)] reg2458 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2456 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2455 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2453 = (1'h0);
  reg [(4'he):(1'h0)] reg2452 = (1'h0);
  reg [(2'h2):(1'h0)] reg2450 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2449 = (1'h0);
  reg [(4'ha):(1'h0)] reg2448 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2446 = (1'h0);
  reg [(4'ha):(1'h0)] reg2443 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2427 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2424 = (1'h0);
  reg [(5'h10):(1'h0)] reg2416 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2445 = (1'h0);
  reg [(4'h8):(1'h0)] reg2444 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2442 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2441 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2439 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2437 = (1'h0);
  reg [(5'h10):(1'h0)] reg2440 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2438 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2436 = (1'h0);
  reg [(4'hc):(1'h0)] reg2434 = (1'h0);
  reg [(4'hf):(1'h0)] reg2433 = (1'h0);
  reg [(3'h7):(1'h0)] reg2432 = (1'h0);
  reg [(4'hf):(1'h0)] reg2431 = (1'h0);
  reg [(4'hf):(1'h0)] reg2430 = (1'h0);
  reg [(3'h5):(1'h0)] reg2429 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2428 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2425 = (1'h0);
  reg [(3'h4):(1'h0)] reg2419 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2423 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2422 = (1'h0);
  reg [(4'hf):(1'h0)] reg2421 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2420 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2418 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2417 = (1'h0);
  reg [(2'h3):(1'h0)] reg2406 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2411 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2415 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2414 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2412 = (1'h0);
  reg [(4'hc):(1'h0)] reg2410 = (1'h0);
  reg [(4'hb):(1'h0)] reg2409 = (1'h0);
  reg [(2'h2):(1'h0)] reg2408 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2407 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2405 = (1'h0);
  reg [(2'h2):(1'h0)] reg2404 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2403 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2400 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2492 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2490 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2488 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2487 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2486 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2478 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2477 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2474 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2469 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2468 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2466 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2462 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2461 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2460 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2459 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2457 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2454 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2451 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2447 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2441 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2444 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2440 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2434 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2430 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2421 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2418 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2443 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2439 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2437 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2435 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2427 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2426 = (1'h0);
  reg [(4'he):(1'h0)] forvar2424 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2419 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2416 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2405 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2413 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2411 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2406 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2402 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2401 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2399 = (1'h0);
  assign y = {wire2500,
                 wire2499,
                 wire2498,
                 wire2497,
                 wire2496,
                 reg2495,
                 reg2494,
                 reg2493,
                 reg2492,
                 reg2487,
                 reg2491,
                 reg2490,
                 reg2489,
                 reg2488,
                 reg2477,
                 reg2485,
                 reg2484,
                 reg2483,
                 reg2482,
                 reg2481,
                 reg2480,
                 reg2479,
                 reg2478,
                 reg2476,
                 reg2475,
                 reg2473,
                 reg2472,
                 reg2471,
                 reg2470,
                 reg2467,
                 reg2465,
                 reg2464,
                 reg2463,
                 reg2458,
                 reg2456,
                 reg2455,
                 reg2453,
                 reg2452,
                 reg2450,
                 reg2449,
                 reg2448,
                 reg2446,
                 reg2443,
                 reg2427,
                 reg2424,
                 reg2416,
                 reg2445,
                 reg2444,
                 reg2442,
                 reg2441,
                 reg2439,
                 reg2437,
                 reg2440,
                 reg2438,
                 reg2436,
                 reg2434,
                 reg2433,
                 reg2432,
                 reg2431,
                 reg2430,
                 reg2429,
                 reg2428,
                 reg2425,
                 reg2419,
                 reg2423,
                 reg2422,
                 reg2421,
                 reg2420,
                 reg2418,
                 reg2417,
                 reg2406,
                 reg2411,
                 reg2415,
                 reg2414,
                 reg2412,
                 reg2410,
                 reg2409,
                 reg2408,
                 reg2407,
                 reg2405,
                 reg2404,
                 reg2403,
                 reg2400,
                 forvar2492,
                 forvar2490,
                 forvar2488,
                 forvar2487,
                 forvar2486,
                 forvar2478,
                 forvar2477,
                 forvar2474,
                 forvar2469,
                 forvar2468,
                 forvar2466,
                 forvar2462,
                 forvar2461,
                 forvar2460,
                 forvar2459,
                 forvar2457,
                 forvar2454,
                 forvar2451,
                 forvar2447,
                 forvar2441,
                 forvar2444,
                 forvar2440,
                 forvar2434,
                 forvar2430,
                 forvar2421,
                 forvar2418,
                 forvar2443,
                 forvar2439,
                 forvar2437,
                 forvar2435,
                 forvar2427,
                 forvar2426,
                 forvar2424,
                 forvar2419,
                 forvar2416,
                 forvar2405,
                 forvar2413,
                 forvar2411,
                 forvar2406,
                 forvar2402,
                 forvar2401,
                 forvar2399,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar2399 = (1'h0); (forvar2399 < (2'h2)); forvar2399 = (forvar2399 + (1'h1)))
        begin
          reg2400 <= $signed(wire2396[(4'ha):(1'h0)]);
          if (wire2394[(4'h8):(2'h3)])
            begin
              for (forvar2401 = (1'h0); (forvar2401 < (1'h1)); forvar2401 = (forvar2401 + (1'h1)))
                begin
                  for (forvar2402 = (1'h0); (forvar2402 < (1'h1)); forvar2402 = (forvar2402 + (1'h1)))
                    begin
                      reg2403 <= forvar2399[(3'h6):(3'h4)];
                      reg2404 <= (^~((+$signed(wire2397)) ?
                          reg2400[(2'h2):(1'h0)] : (^~wire2396[(2'h3):(2'h2)])));
                      reg2405 <= forvar2399[(3'h6):(1'h0)];
                    end
                  for (forvar2406 = (1'h0); (forvar2406 < (2'h3)); forvar2406 = (forvar2406 + (1'h1)))
                    begin
                      reg2407 <= $unsigned(($signed((reg2404 - wire2397)) ?
                          (-$unsigned(reg2400)) : ((reg2405 == wire2397) ?
                              forvar2406[(3'h7):(3'h4)] : $unsigned(forvar2402))));
                      reg2408 <= wire2394;
                    end
                end
              reg2409 <= wire2397[(4'hb):(1'h1)];
              reg2410 <= (~((-$signed(reg2404)) ? reg2408 : wire2398));
              if (({wire2394} + reg2409))
                begin
                  for (forvar2411 = (1'h0); (forvar2411 < (2'h3)); forvar2411 = (forvar2411 + (1'h1)))
                    begin
                      reg2412 <= $signed($signed(((reg2403 && reg2400) ?
                          $unsigned(reg2408) : reg2409)));
                    end
                  for (forvar2413 = (1'h0); (forvar2413 < (2'h2)); forvar2413 = (forvar2413 + (1'h1)))
                    begin
                      reg2414 <= $signed(($signed($unsigned(reg2409)) ?
                          (wire2397 ?
                              forvar2406 : (reg2405 ?
                                  reg2403 : wire2395)) : $unsigned(forvar2401)));
                      reg2415 <= (+(($unsigned(forvar2406) ~^ (reg2408 >>> forvar2413)) ^~ (+(wire2397 && wire2398))));
                    end
                end
              else
                begin
                  if (forvar2402)
                    begin
                      reg2411 <= $signed(reg2405);
                    end
                  else
                    begin
                      reg2411 <= wire2397;
                      reg2412 <= $unsigned($signed(reg2405));
                    end
                end
            end
          else
            begin
              for (forvar2401 = (1'h0); (forvar2401 < (2'h3)); forvar2401 = (forvar2401 + (1'h1)))
                begin
                  for (forvar2402 = (1'h0); (forvar2402 < (2'h3)); forvar2402 = (forvar2402 + (1'h1)))
                    begin
                      reg2403 <= $unsigned(reg2400);
                    end
                  reg2404 <= $signed($signed((~&reg2405[(3'h6):(2'h3)])));
                  for (forvar2405 = (1'h0); (forvar2405 < (2'h2)); forvar2405 = (forvar2405 + (1'h1)))
                    begin
                      reg2406 <= forvar2413[(1'h1):(1'h1)];
                    end
                  if ($unsigned(forvar2402))
                    begin
                      reg2407 <= (($unsigned($signed(wire2395)) << $unsigned(reg2404)) ?
                          (^~{{wire2395}}) : ((8'hb4) | ($signed(forvar2401) || reg2412)));
                      reg2408 <= $unsigned(forvar2401[(1'h1):(1'h0)]);
                      reg2409 <= ($signed(((~&reg2407) ?
                              reg2409[(3'h6):(2'h2)] : {(8'h9e)})) ?
                          reg2414[(1'h0):(1'h0)] : (~^$unsigned(reg2412[(4'hb):(3'h7)])));
                    end
                  else
                    begin
                      reg2407 <= $unsigned((|{{wire2396}}));
                      reg2408 <= (~|$signed((!$unsigned(wire2395))));
                    end
                end
            end
        end
      if ($unsigned((((~|forvar2406) * {forvar2401}) == $signed(((8'h9f) ?
          reg2405 : reg2406)))))
        begin
          for (forvar2416 = (1'h0); (forvar2416 < (1'h1)); forvar2416 = (forvar2416 + (1'h1)))
            begin
              if ($signed((~$unsigned(forvar2406[(3'h4):(1'h1)]))))
                begin
                  if ((~^wire2395[(3'h7):(3'h6)]))
                    begin
                      reg2417 <= (8'haa);
                      reg2418 <= $unsigned(reg2407[(3'h5):(3'h5)]);
                    end
                  else
                    begin
                      reg2417 <= ((($unsigned((8'hb2)) <<< (8'had)) == (forvar2401 ?
                          $unsigned(forvar2411) : {forvar2406})) ^ $signed(reg2412[(4'hb):(3'h5)]));
                    end
                  for (forvar2419 = (1'h0); (forvar2419 < (1'h1)); forvar2419 = (forvar2419 + (1'h1)))
                    begin
                      reg2420 <= $unsigned($signed((-forvar2405[(1'h1):(1'h0)])));
                      reg2421 <= (&wire2395[(1'h0):(1'h0)]);
                      reg2422 <= reg2400[(1'h1):(1'h1)];
                    end
                  reg2423 <= $unsigned({(((8'h9d) ?
                          reg2421 : reg2422) * $unsigned((8'hb8)))});
                end
              else
                begin
                  if (forvar2402)
                    begin
                      reg2417 <= (-reg2406[(1'h1):(1'h0)]);
                      reg2418 <= ((~((~^wire2395) ?
                          $unsigned((8'hb9)) : forvar2405[(2'h3):(1'h1)])) >>> (+forvar2399[(4'h9):(4'h9)]));
                      reg2419 <= wire2397;
                    end
                  else
                    begin
                      reg2417 <= (~|reg2422[(3'h4):(2'h3)]);
                      reg2418 <= reg2415[(3'h7):(3'h5)];
                      reg2419 <= reg2409;
                      reg2420 <= $unsigned(reg2421);
                    end
                  if ($unsigned({($signed(forvar2402) ?
                          reg2411 : $signed((8'hba)))}))
                    begin
                      reg2421 <= reg2403[(1'h1):(1'h1)];
                      reg2422 <= (8'hac);
                      reg2423 <= ((-$unsigned(forvar2405)) ?
                          $signed(reg2403[(2'h3):(2'h3)]) : (!((reg2423 ?
                              reg2414 : reg2415) && (forvar2399 >= wire2394))));
                    end
                  else
                    begin
                      reg2421 <= $signed($unsigned($signed($unsigned((8'hb3)))));
                      reg2422 <= wire2395;
                      reg2423 <= (8'hac);
                    end
                  for (forvar2424 = (1'h0); (forvar2424 < (1'h0)); forvar2424 = (forvar2424 + (1'h1)))
                    begin
                      reg2425 <= $unsigned($signed((reg2400[(1'h0):(1'h0)] ?
                          $signed(reg2415) : reg2422)));
                    end
                end
              for (forvar2426 = (1'h0); (forvar2426 < (1'h0)); forvar2426 = (forvar2426 + (1'h1)))
                begin
                  for (forvar2427 = (1'h0); (forvar2427 < (1'h1)); forvar2427 = (forvar2427 + (1'h1)))
                    begin
                      reg2428 <= forvar2424[(4'h9):(4'h9)];
                      reg2429 <= (|forvar2427[(3'h6):(1'h0)]);
                      reg2430 <= ($signed($unsigned((8'ha1))) + reg2410[(3'h5):(3'h5)]);
                      reg2431 <= forvar2419[(3'h6):(2'h2)];
                    end
                  if ((!$unsigned(($unsigned(reg2431) ?
                      wire2394[(2'h2):(1'h1)] : $signed(reg2400)))))
                    begin
                      reg2432 <= forvar2419[(3'h7):(1'h0)];
                      reg2433 <= $signed($signed(((~^reg2420) << (forvar2399 ?
                          reg2431 : reg2429))));
                      reg2434 <= forvar2405[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2432 <= reg2421;
                    end
                  for (forvar2435 = (1'h0); (forvar2435 < (2'h2)); forvar2435 = (forvar2435 + (1'h1)))
                    begin
                      reg2436 <= (^~({(reg2420 ?
                              (8'hae) : reg2405)} != ($unsigned((8'hb5)) >>> wire2394[(4'h8):(4'h8)])));
                    end
                end
            end
          if (reg2405)
            begin
              for (forvar2437 = (1'h0); (forvar2437 < (1'h0)); forvar2437 = (forvar2437 + (1'h1)))
                begin
                  reg2438 <= reg2415;
                  for (forvar2439 = (1'h0); (forvar2439 < (2'h2)); forvar2439 = (forvar2439 + (1'h1)))
                    begin
                      reg2440 <= ((8'ha5) ?
                          $signed($unsigned((8'ha1))) : $unsigned((~|reg2430)));
                    end
                end
            end
          else
            begin
              if ($unsigned(reg2422[(2'h2):(1'h0)]))
                begin
                  if ($unsigned((^~reg2412[(1'h1):(1'h0)])))
                    begin
                      reg2437 <= reg2410[(2'h3):(1'h0)];
                      reg2438 <= $unsigned(((8'hb0) + reg2409));
                      reg2439 <= reg2400[(2'h2):(2'h2)];
                      reg2440 <= {reg2410};
                    end
                  else
                    begin
                      reg2437 <= reg2429;
                      reg2438 <= (~^$unsigned(reg2410));
                      reg2439 <= reg2431[(1'h0):(1'h0)];
                    end
                  reg2441 <= reg2400;
                  reg2442 <= forvar2411;
                end
              else
                begin
                  reg2437 <= $signed($unsigned($signed(((8'ha6) ?
                      reg2403 : reg2406))));
                  reg2438 <= ($unsigned((~&(forvar2419 ^~ (8'h9e)))) + $signed(((reg2431 >>> reg2440) ?
                      (reg2433 >= forvar2427) : (~reg2404))));
                  for (forvar2439 = (1'h0); (forvar2439 < (2'h2)); forvar2439 = (forvar2439 + (1'h1)))
                    begin
                      reg2440 <= (^(reg2414[(2'h2):(2'h2)] >= forvar2402));
                      reg2441 <= (forvar2413 >= {((forvar2435 ?
                                  reg2415 : reg2405) ?
                              (reg2412 ? (8'ha8) : reg2437) : reg2436)});
                      reg2442 <= $unsigned(forvar2435);
                    end
                  for (forvar2443 = (1'h0); (forvar2443 < (2'h2)); forvar2443 = (forvar2443 + (1'h1)))
                    begin
                      reg2444 <= reg2403[(1'h0):(1'h0)];
                      reg2445 <= wire2396[(3'h4):(2'h2)];
                    end
                end
            end
        end
      else
        begin
          if (reg2406[(1'h0):(1'h0)])
            begin
              if ((~^$signed($signed(reg2417))))
                begin
                  reg2416 <= {reg2409};
                  if ($signed((8'ha5)))
                    begin
                      reg2417 <= (reg2406[(2'h3):(2'h2)] ~^ wire2398[(1'h1):(1'h0)]);
                      reg2418 <= ($unsigned(((|reg2442) & ((8'hb0) ?
                          reg2438 : reg2442))) > ((~&reg2406) ?
                          reg2438[(1'h0):(1'h0)] : (((8'ha4) ^ reg2437) ?
                              $signed(reg2431) : (wire2398 ^~ forvar2402))));
                      reg2419 <= $unsigned(forvar2435[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg2417 <= (~^reg2434[(3'h6):(2'h2)]);
                    end
                end
              else
                begin
                  for (forvar2416 = (1'h0); (forvar2416 < (1'h1)); forvar2416 = (forvar2416 + (1'h1)))
                    begin
                      reg2417 <= ($signed((reg2420 ?
                          (wire2396 == forvar2437) : $signed(reg2431))) ~^ ((8'hba) ?
                          (wire2397[(3'h5):(2'h3)] < $signed(reg2441)) : (~(+reg2404))));
                    end
                  for (forvar2418 = (1'h0); (forvar2418 < (1'h0)); forvar2418 = (forvar2418 + (1'h1)))
                    begin
                      reg2419 <= $unsigned($signed((reg2421[(3'h6):(3'h4)] >>> $signed(forvar2416))));
                      reg2420 <= (({reg2420[(1'h0):(1'h0)]} <= forvar2416) ?
                          $signed($unsigned(forvar2413)) : reg2404);
                      reg2421 <= reg2420[(2'h3):(2'h2)];
                      reg2422 <= $unsigned(($signed((reg2415 * reg2437)) ?
                          (-reg2404) : $signed((reg2433 ?
                              reg2440 : forvar2411))));
                    end
                  reg2423 <= {({(reg2445 ? reg2432 : reg2438)} ?
                          (reg2407 ?
                              (wire2397 || (8'hab)) : reg2444) : ((reg2429 ?
                              reg2400 : reg2429) > (8'ha4)))};
                end
            end
          else
            begin
              if ($signed(reg2438))
                begin
                  for (forvar2416 = (1'h0); (forvar2416 < (1'h0)); forvar2416 = (forvar2416 + (1'h1)))
                    begin
                      reg2417 <= (^~$signed(forvar2419[(1'h1):(1'h0)]));
                      reg2418 <= (~|reg2405);
                      reg2419 <= reg2432[(1'h1):(1'h0)];
                      reg2420 <= forvar2401;
                    end
                end
              else
                begin
                  for (forvar2416 = (1'h0); (forvar2416 < (1'h1)); forvar2416 = (forvar2416 + (1'h1)))
                    begin
                      reg2417 <= reg2438;
                      reg2418 <= reg2407[(2'h2):(2'h2)];
                    end
                  for (forvar2419 = (1'h0); (forvar2419 < (1'h1)); forvar2419 = (forvar2419 + (1'h1)))
                    begin
                      reg2420 <= (8'ha3);
                    end
                end
              if ((!$unsigned($unsigned((-(8'haf))))))
                begin
                  if ($unsigned({reg2409}))
                    begin
                      reg2421 <= reg2414[(2'h2):(2'h2)];
                      reg2422 <= $signed((((reg2420 >>> (8'h9d)) ?
                              $unsigned(reg2406) : (~forvar2435)) ?
                          ($signed(reg2438) ?
                              {reg2440} : (8'ha3)) : {reg2414}));
                      reg2423 <= {(reg2440 - ($unsigned(reg2441) == (reg2432 ?
                              reg2415 : reg2437)))};
                      reg2424 <= reg2439;
                    end
                  else
                    begin
                      reg2421 <= ((forvar2406[(3'h5):(3'h4)] ?
                              {(|reg2442)} : ($signed(forvar2413) ?
                                  (+reg2417) : $unsigned((8'hb2)))) ?
                          $unsigned($unsigned(forvar2406)) : (8'hb3));
                      reg2422 <= $unsigned($unsigned(reg2439[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar2421 = (1'h0); (forvar2421 < (2'h3)); forvar2421 = (forvar2421 + (1'h1)))
                    begin
                      reg2422 <= ($unsigned(reg2434[(2'h2):(2'h2)]) ?
                          {reg2434} : (forvar2418[(3'h4):(1'h0)] ?
                              (&(forvar2402 ? reg2410 : reg2440)) : reg2430));
                      reg2423 <= ($unsigned(((^~wire2398) << $unsigned(reg2415))) ?
                          {($unsigned(reg2400) ?
                                  reg2441 : (8'hb1))} : (&reg2419));
                      reg2424 <= $unsigned($unsigned(((forvar2439 < reg2438) ?
                          (^~reg2418) : reg2429[(1'h1):(1'h1)])));
                      reg2425 <= ((-reg2411) | {(reg2414[(1'h0):(1'h0)] >> (reg2419 != forvar2426))});
                    end
                end
              for (forvar2426 = (1'h0); (forvar2426 < (2'h2)); forvar2426 = (forvar2426 + (1'h1)))
                begin
                  if (reg2414)
                    begin
                      reg2427 <= reg2407;
                      reg2428 <= $signed(forvar2411);
                      reg2429 <= (|reg2434);
                    end
                  else
                    begin
                      reg2427 <= $signed((8'haa));
                    end
                  for (forvar2430 = (1'h0); (forvar2430 < (1'h1)); forvar2430 = (forvar2430 + (1'h1)))
                    begin
                      reg2431 <= {$signed((reg2404[(1'h0):(1'h0)] & (forvar2419 < forvar2416)))};
                      reg2432 <= {((((8'h9f) ? reg2404 : wire2394) ?
                                  (&forvar2430) : {forvar2443}) ?
                              $unsigned(reg2432[(1'h1):(1'h0)]) : {{reg2437}})};
                    end
                  reg2433 <= ($signed({$signed(reg2417)}) > forvar2437);
                end
              for (forvar2434 = (1'h0); (forvar2434 < (1'h1)); forvar2434 = (forvar2434 + (1'h1)))
                begin
                  for (forvar2435 = (1'h0); (forvar2435 < (1'h0)); forvar2435 = (forvar2435 + (1'h1)))
                    begin
                      reg2436 <= $unsigned(((^~((8'hb4) ?
                          forvar2399 : reg2436)) - (~&(reg2414 ?
                          reg2412 : reg2414))));
                      reg2437 <= ((~$unsigned($signed(reg2412))) ?
                          $signed((&(+wire2397))) : {(wire2397[(4'h8):(2'h3)] <<< (forvar2399 ?
                                  wire2398 : wire2395))});
                      reg2438 <= (((-(reg2433 + (8'hb8))) ^ (8'hb1)) >>> (~^$unsigned({wire2396})));
                      reg2439 <= $signed(reg2442);
                    end
                end
            end
          for (forvar2440 = (1'h0); (forvar2440 < (2'h3)); forvar2440 = (forvar2440 + (1'h1)))
            begin
              if ((!wire2395[(4'he):(4'hd)]))
                begin
                  if ({forvar2437})
                    begin
                      reg2441 <= reg2415;
                      reg2442 <= (+$signed(($signed((8'h9d)) ?
                          reg2430 : $signed(forvar2443))));
                      reg2443 <= forvar2399;
                    end
                  else
                    begin
                      reg2441 <= forvar2440[(3'h4):(3'h4)];
                      reg2442 <= forvar2411;
                      reg2443 <= ((((reg2400 ?
                                  forvar2437 : reg2442) >> $signed(wire2394)) ?
                              (+{forvar2406}) : ((reg2438 ?
                                      forvar2413 : forvar2439) ?
                                  $signed((8'hab)) : $signed((8'hb7)))) ?
                          ($unsigned(reg2431[(4'ha):(2'h3)]) ?
                              (!$signed((8'ha9))) : $signed((+reg2415))) : forvar2406);
                    end
                  for (forvar2444 = (1'h0); (forvar2444 < (1'h0)); forvar2444 = (forvar2444 + (1'h1)))
                    begin
                      reg2445 <= ($unsigned(forvar2443[(3'h6):(2'h2)]) ?
                          (~$unsigned((~&forvar2434))) : $unsigned($unsigned(forvar2419)));
                    end
                end
              else
                begin
                  for (forvar2441 = (1'h0); (forvar2441 < (1'h1)); forvar2441 = (forvar2441 + (1'h1)))
                    begin
                      reg2442 <= $unsigned($unsigned(reg2436[(3'h4):(2'h3)]));
                      reg2443 <= reg2436[(2'h3):(2'h3)];
                    end
                end
              reg2446 <= $signed(reg2414);
              for (forvar2447 = (1'h0); (forvar2447 < (1'h1)); forvar2447 = (forvar2447 + (1'h1)))
                begin
                  if ((!(~|$signed((|reg2424)))))
                    begin
                      reg2448 <= $unsigned((reg2404 ^ (reg2432[(3'h7):(3'h6)] ?
                          (8'had) : $unsigned(forvar2447))));
                      reg2449 <= $unsigned((((+forvar2430) ?
                          reg2405 : {reg2427}) <= {(reg2438 ?
                              forvar2411 : (8'ha8))}));
                    end
                  else
                    begin
                      reg2448 <= ($signed(forvar2399[(4'hc):(4'hb)]) == $signed(((reg2415 ?
                              reg2407 : reg2449) ?
                          (forvar2424 ?
                              forvar2413 : wire2398) : $unsigned(reg2400))));
                      reg2449 <= $unsigned(($unsigned(reg2427[(4'hd):(3'h6)]) ?
                          reg2436 : forvar2402));
                      reg2450 <= ((&$signed($signed(wire2394))) <= forvar2411);
                    end
                  for (forvar2451 = (1'h0); (forvar2451 < (2'h2)); forvar2451 = (forvar2451 + (1'h1)))
                    begin
                      reg2452 <= forvar2424;
                      reg2453 <= reg2421[(2'h3):(1'h1)];
                    end
                  for (forvar2454 = (1'h0); (forvar2454 < (2'h2)); forvar2454 = (forvar2454 + (1'h1)))
                    begin
                      reg2455 <= $signed(((reg2438 | (reg2430 ?
                              (8'hb6) : reg2403)) ?
                          forvar2426[(1'h1):(1'h1)] : {{(8'ha3)}}));
                      reg2456 <= {reg2421};
                    end
                  for (forvar2457 = (1'h0); (forvar2457 < (2'h2)); forvar2457 = (forvar2457 + (1'h1)))
                    begin
                      reg2458 <= (($unsigned((reg2420 ? reg2446 : reg2410)) ?
                              reg2421[(4'hc):(3'h5)] : forvar2421[(4'h9):(3'h6)]) ?
                          (8'haa) : ($unsigned((+reg2421)) ?
                              reg2406[(2'h2):(1'h0)] : forvar2426));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2459 = (1'h0); (forvar2459 < (1'h1)); forvar2459 = (forvar2459 + (1'h1)))
        begin
          for (forvar2460 = (1'h0); (forvar2460 < (2'h2)); forvar2460 = (forvar2460 + (1'h1)))
            begin
              for (forvar2461 = (1'h0); (forvar2461 < (1'h0)); forvar2461 = (forvar2461 + (1'h1)))
                begin
                  for (forvar2462 = (1'h0); (forvar2462 < (1'h0)); forvar2462 = (forvar2462 + (1'h1)))
                    begin
                      reg2463 <= $unsigned(({$signed(reg2441)} | {reg2429[(1'h0):(1'h0)]}));
                      reg2464 <= (~&reg2408[(1'h0):(1'h0)]);
                      reg2465 <= ((~|{(wire2397 ?
                              reg2406 : reg2446)}) + (^reg2414[(1'h0):(1'h0)]));
                    end
                end
            end
          for (forvar2466 = (1'h0); (forvar2466 < (1'h1)); forvar2466 = (forvar2466 + (1'h1)))
            begin
              reg2467 <= $unsigned(($signed((reg2434 ?
                  (8'hb8) : (8'hb3))) <= reg2428[(3'h5):(3'h4)]));
              for (forvar2468 = (1'h0); (forvar2468 < (1'h1)); forvar2468 = (forvar2468 + (1'h1)))
                begin
                  for (forvar2469 = (1'h0); (forvar2469 < (1'h1)); forvar2469 = (forvar2469 + (1'h1)))
                    begin
                      reg2470 <= ({$unsigned(reg2465)} - $signed(((+reg2403) >> $unsigned(reg2446))));
                      reg2471 <= $unsigned((~((8'ha5) != reg2418[(1'h0):(1'h0)])));
                      reg2472 <= ($signed((reg2417 <<< $signed(wire2397))) && reg2403[(2'h3):(1'h0)]);
                      reg2473 <= (+((((8'hb9) ?
                          reg2445 : reg2421) <= reg2436) >= $signed(reg2424)));
                    end
                  for (forvar2474 = (1'h0); (forvar2474 < (2'h2)); forvar2474 = (forvar2474 + (1'h1)))
                    begin
                      reg2475 <= reg2473[(4'ha):(1'h1)];
                      reg2476 <= $unsigned($unsigned($signed((reg2441 ^ reg2405))));
                    end
                end
              if ((forvar2460 ?
                  ($signed(((8'hab) || reg2473)) == (reg2440 ?
                      $unsigned((8'haa)) : (reg2464 == reg2409))) : (-(^$signed(reg2415)))))
                begin
                  for (forvar2477 = (1'h0); (forvar2477 < (2'h2)); forvar2477 = (forvar2477 + (1'h1)))
                    begin
                      reg2478 <= ((-(~^reg2452)) >> $unsigned((8'hb8)));
                      reg2479 <= reg2410[(4'ha):(3'h6)];
                      reg2480 <= {$signed($signed(reg2414[(1'h1):(1'h1)]))};
                      reg2481 <= {wire2397};
                    end
                  if ($signed(($unsigned($signed(reg2403)) ?
                      {reg2439[(1'h0):(1'h0)]} : reg2406)))
                    begin
                      reg2482 <= $unsigned(forvar2461[(4'hf):(4'h8)]);
                      reg2483 <= {reg2417};
                      reg2484 <= (((^~$signed(forvar2466)) ?
                              (reg2449[(3'h4):(3'h4)] >>> (^reg2478)) : $unsigned({forvar2468})) ?
                          (~^reg2415) : reg2444[(3'h5):(1'h0)]);
                      reg2485 <= $unsigned($unsigned((8'hb1)));
                    end
                  else
                    begin
                      reg2482 <= {(^$unsigned(reg2445))};
                      reg2483 <= (8'ha3);
                      reg2484 <= reg2403[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  reg2477 <= (8'hb9);
                  for (forvar2478 = (1'h0); (forvar2478 < (1'h0)); forvar2478 = (forvar2478 + (1'h1)))
                    begin
                      reg2479 <= {(|((reg2476 ?
                              reg2478 : reg2445) && forvar2478))};
                    end
                  if ({forvar2477[(3'h4):(3'h4)]})
                    begin
                      reg2480 <= reg2448;
                    end
                  else
                    begin
                      reg2480 <= reg2456;
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2486 = (1'h0); (forvar2486 < (1'h0)); forvar2486 = (forvar2486 + (1'h1)))
        begin
          if (reg2428)
            begin
              if ({$unsigned(((forvar2486 ? reg2432 : (8'ha4)) ?
                      $unsigned(reg2429) : reg2427[(4'h9):(1'h0)]))})
                begin
                  for (forvar2487 = (1'h0); (forvar2487 < (2'h2)); forvar2487 = (forvar2487 + (1'h1)))
                    begin
                      reg2488 <= reg2428;
                      reg2489 <= reg2411;
                      reg2490 <= (~$signed($unsigned(reg2419)));
                      reg2491 <= (8'hb3);
                    end
                end
              else
                begin
                  if ($unsigned({($signed(reg2429) > $signed(reg2475))}))
                    begin
                      reg2487 <= reg2403[(1'h0):(1'h0)];
                      reg2488 <= reg2481[(2'h2):(2'h2)];
                      reg2489 <= $unsigned(reg2446);
                    end
                  else
                    begin
                      reg2487 <= reg2418[(1'h0):(1'h0)];
                    end
                  if ($signed((({(8'haf)} ?
                      (reg2404 && (8'hae)) : {reg2482}) >>> (^~reg2420))))
                    begin
                      reg2490 <= $signed($signed(reg2477));
                      reg2491 <= (~&$signed((reg2409 ~^ reg2444[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg2490 <= reg2470[(2'h3):(1'h1)];
                      reg2491 <= (reg2405[(3'h5):(2'h2)] << (wire2394[(3'h6):(3'h5)] ?
                          reg2482[(4'ha):(3'h5)] : (((8'ha3) ?
                                  reg2456 : forvar2487) ?
                              (&reg2443) : $signed(reg2414))));
                      reg2492 <= $unsigned(({(^~reg2427)} ^~ $unsigned($unsigned(reg2450))));
                    end
                  reg2493 <= reg2479;
                end
            end
          else
            begin
              reg2487 <= ((^(~|reg2442)) ^~ ($signed(reg2476) ?
                  (reg2433[(4'hc):(3'h4)] ?
                      (-(8'hb8)) : $unsigned(reg2487)) : wire2397[(3'h5):(3'h5)]));
              for (forvar2488 = (1'h0); (forvar2488 < (2'h3)); forvar2488 = (forvar2488 + (1'h1)))
                begin
                  reg2489 <= ((((8'had) ?
                      $unsigned((8'hb3)) : reg2481) < reg2417) & {((reg2458 ?
                          (8'h9f) : reg2487) + reg2446[(3'h6):(1'h1)])});
                end
              for (forvar2490 = (1'h0); (forvar2490 < (2'h2)); forvar2490 = (forvar2490 + (1'h1)))
                begin
                  if ((8'ha6))
                    begin
                      reg2491 <= reg2419[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2491 <= reg2405[(1'h1):(1'h0)];
                    end
                  for (forvar2492 = (1'h0); (forvar2492 < (2'h3)); forvar2492 = (forvar2492 + (1'h1)))
                    begin
                      reg2493 <= (!reg2482[(4'hc):(2'h3)]);
                      reg2494 <= ((reg2419 ?
                          $unsigned(reg2433) : (8'hac)) <<< (reg2481[(4'h9):(3'h5)] | $signed(reg2458)));
                    end
                end
              reg2495 <= ((-$unsigned($signed(reg2488))) ?
                  reg2490[(4'hb):(3'h5)] : reg2439);
            end
        end
    end
  assign wire2496 = $signed($signed(wire2395[(4'hd):(4'hb)]));
  assign wire2497 = ((({(8'hae)} ~^ reg2415) * (((8'had) >>> reg2410) == reg2473[(3'h5):(1'h0)])) + {reg2484});
  assign wire2498 = $unsigned(((8'hb9) <= reg2405[(4'ha):(1'h0)]));
  assign wire2499 = {reg2449[(1'h0):(1'h0)]};
  assign wire2500 = ({((reg2430 ? (8'hb9) : reg2484) ?
                                (&reg2472) : (reg2407 <= reg2452))} ?
                        reg2484 : (reg2409[(2'h3):(2'h3)] ^~ reg2479));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3056  (y, clk, wire3060, wire3059, wire3058, wire3057);
  output wire [(32'hd67):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire3060;
  input wire signed [(3'h7):(1'h0)] wire3059;
  input wire signed [(4'hc):(1'h0)] wire3058;
  input wire [(3'h7):(1'h0)] wire3057;
  wire [(3'h7):(1'h0)] wire3271;
  wire signed [(4'hd):(1'h0)] wire3270;
  wire signed [(4'hc):(1'h0)] wire3269;
  wire [(4'he):(1'h0)] wire3268;
  wire [(3'h7):(1'h0)] wire3267;
  wire signed [(4'h8):(1'h0)] wire3177;
  wire [(4'hc):(1'h0)] wire3176;
  wire signed [(4'hf):(1'h0)] wire3175;
  wire [(4'he):(1'h0)] wire3174;
  wire [(4'ha):(1'h0)] wire3173;
  wire [(5'h10):(1'h0)] wire3064;
  wire signed [(3'h5):(1'h0)] wire3063;
  wire [(3'h5):(1'h0)] wire3062;
  wire signed [(4'ha):(1'h0)] wire3061;
  reg [(4'ha):(1'h0)] reg3384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3383 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3382 = (1'h0);
  reg [(4'hb):(1'h0)] reg3381 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3379 = (1'h0);
  reg [(4'ha):(1'h0)] reg3378 = (1'h0);
  reg [(4'hd):(1'h0)] reg3377 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3375 = (1'h0);
  reg [(3'h6):(1'h0)] reg3374 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3373 = (1'h0);
  reg [(4'ha):(1'h0)] reg3372 = (1'h0);
  reg [(4'hb):(1'h0)] reg3371 = (1'h0);
  reg [(4'hf):(1'h0)] reg3370 = (1'h0);
  reg [(3'h6):(1'h0)] reg3369 = (1'h0);
  reg [(4'hf):(1'h0)] reg3368 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3366 = (1'h0);
  reg [(4'h9):(1'h0)] reg3365 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3364 = (1'h0);
  reg [(4'hc):(1'h0)] reg3362 = (1'h0);
  reg [(2'h3):(1'h0)] reg3352 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3359 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3356 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3355 = (1'h0);
  reg [(3'h4):(1'h0)] reg3354 = (1'h0);
  reg [(2'h2):(1'h0)] reg3353 = (1'h0);
  reg [(4'hc):(1'h0)] reg3351 = (1'h0);
  reg [(2'h3):(1'h0)] reg3350 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3349 = (1'h0);
  reg [(3'h7):(1'h0)] reg3348 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3346 = (1'h0);
  reg [(4'hf):(1'h0)] reg3345 = (1'h0);
  reg [(4'he):(1'h0)] reg3340 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3344 = (1'h0);
  reg [(3'h6):(1'h0)] reg3343 = (1'h0);
  reg [(4'hc):(1'h0)] reg3342 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3341 = (1'h0);
  reg [(4'hd):(1'h0)] reg3323 = (1'h0);
  reg [(4'hd):(1'h0)] reg3339 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3334 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3338 = (1'h0);
  reg [(4'h9):(1'h0)] reg3337 = (1'h0);
  reg [(4'h8):(1'h0)] reg3336 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3335 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3333 = (1'h0);
  reg [(3'h4):(1'h0)] reg3332 = (1'h0);
  reg [(4'h9):(1'h0)] reg3331 = (1'h0);
  reg [(4'ha):(1'h0)] reg3329 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3328 = (1'h0);
  reg [(4'hc):(1'h0)] reg3327 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3326 = (1'h0);
  reg [(4'ha):(1'h0)] reg3325 = (1'h0);
  reg [(5'h10):(1'h0)] reg3324 = (1'h0);
  reg [(4'he):(1'h0)] reg3322 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3321 = (1'h0);
  reg [(3'h6):(1'h0)] reg3320 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3319 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3318 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3317 = (1'h0);
  reg [(2'h3):(1'h0)] reg3316 = (1'h0);
  reg [(4'h9):(1'h0)] reg3315 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3313 = (1'h0);
  reg [(5'h10):(1'h0)] reg3311 = (1'h0);
  reg [(3'h6):(1'h0)] reg3310 = (1'h0);
  reg [(4'hf):(1'h0)] reg3309 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3308 = (1'h0);
  reg [(2'h2):(1'h0)] reg3307 = (1'h0);
  reg [(3'h4):(1'h0)] reg3306 = (1'h0);
  reg [(4'hc):(1'h0)] reg3305 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3304 = (1'h0);
  reg [(4'hc):(1'h0)] reg3302 = (1'h0);
  reg [(3'h4):(1'h0)] reg3301 = (1'h0);
  reg [(3'h6):(1'h0)] reg3300 = (1'h0);
  reg [(4'h9):(1'h0)] reg3299 = (1'h0);
  reg [(4'h8):(1'h0)] reg3298 = (1'h0);
  reg [(4'h8):(1'h0)] reg3297 = (1'h0);
  reg [(4'hf):(1'h0)] reg3296 = (1'h0);
  reg [(4'ha):(1'h0)] reg3295 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3294 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3290 = (1'h0);
  reg [(4'hd):(1'h0)] reg3289 = (1'h0);
  reg [(4'hb):(1'h0)] reg3288 = (1'h0);
  reg [(4'hb):(1'h0)] reg3287 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3284 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3280 = (1'h0);
  reg [(3'h6):(1'h0)] reg3275 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3274 = (1'h0);
  reg [(4'hd):(1'h0)] reg3286 = (1'h0);
  reg [(4'h9):(1'h0)] reg3285 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3283 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3282 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3281 = (1'h0);
  reg [(3'h4):(1'h0)] reg3279 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3278 = (1'h0);
  reg [(4'hc):(1'h0)] reg3277 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3276 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3273 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3272 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3266 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3263 = (1'h0);
  reg [(4'hf):(1'h0)] reg3255 = (1'h0);
  reg [(4'he):(1'h0)] reg3262 = (1'h0);
  reg [(3'h5):(1'h0)] reg3260 = (1'h0);
  reg [(3'h7):(1'h0)] reg3261 = (1'h0);
  reg [(2'h3):(1'h0)] reg3259 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3258 = (1'h0);
  reg [(4'he):(1'h0)] reg3257 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3256 = (1'h0);
  reg [(4'h8):(1'h0)] reg3254 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3253 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3250 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3249 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3243 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3248 = (1'h0);
  reg [(3'h6):(1'h0)] reg3247 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3246 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3245 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3244 = (1'h0);
  reg [(4'hf):(1'h0)] reg3242 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3233 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3232 = (1'h0);
  reg [(2'h2):(1'h0)] reg3227 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3225 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3241 = (1'h0);
  reg [(4'hc):(1'h0)] reg3240 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3239 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3238 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3237 = (1'h0);
  reg [(2'h3):(1'h0)] reg3235 = (1'h0);
  reg [(4'hf):(1'h0)] reg3234 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3231 = (1'h0);
  reg [(5'h10):(1'h0)] reg3230 = (1'h0);
  reg [(4'hf):(1'h0)] reg3229 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3228 = (1'h0);
  reg [(4'h9):(1'h0)] reg3226 = (1'h0);
  reg [(4'hc):(1'h0)] reg3224 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3221 = (1'h0);
  reg [(3'h6):(1'h0)] reg3220 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3219 = (1'h0);
  reg [(2'h2):(1'h0)] reg3218 = (1'h0);
  reg [(2'h3):(1'h0)] reg3217 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3216 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3215 = (1'h0);
  reg [(2'h2):(1'h0)] reg3209 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3214 = (1'h0);
  reg [(4'ha):(1'h0)] reg3213 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3212 = (1'h0);
  reg [(4'hb):(1'h0)] reg3211 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3210 = (1'h0);
  reg [(4'hc):(1'h0)] reg3208 = (1'h0);
  reg [(4'hf):(1'h0)] reg3207 = (1'h0);
  reg [(3'h4):(1'h0)] reg3206 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3204 = (1'h0);
  reg [(2'h2):(1'h0)] reg3203 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3202 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3201 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3200 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3199 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3198 = (1'h0);
  reg [(3'h5):(1'h0)] reg3197 = (1'h0);
  reg [(4'he):(1'h0)] reg3196 = (1'h0);
  reg [(4'he):(1'h0)] reg3195 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3194 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3193 = (1'h0);
  reg [(5'h10):(1'h0)] reg3191 = (1'h0);
  reg [(4'ha):(1'h0)] reg3190 = (1'h0);
  reg [(4'hc):(1'h0)] reg3189 = (1'h0);
  reg [(3'h4):(1'h0)] reg3187 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3186 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3185 = (1'h0);
  reg [(3'h6):(1'h0)] reg3184 = (1'h0);
  reg [(4'hf):(1'h0)] reg3183 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3182 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3181 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3172 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3171 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3170 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3169 = (1'h0);
  reg [(2'h2):(1'h0)] reg3168 = (1'h0);
  reg [(4'he):(1'h0)] reg3166 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3165 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3163 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3161 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3160 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3159 = (1'h0);
  reg [(3'h6):(1'h0)] reg3158 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3157 = (1'h0);
  reg [(4'hf):(1'h0)] reg3155 = (1'h0);
  reg [(4'hc):(1'h0)] reg3154 = (1'h0);
  reg [(4'ha):(1'h0)] reg3153 = (1'h0);
  reg [(5'h10):(1'h0)] reg3152 = (1'h0);
  reg [(3'h4):(1'h0)] reg3150 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3149 = (1'h0);
  reg [(4'h8):(1'h0)] reg3148 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3147 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3145 = (1'h0);
  reg [(4'hb):(1'h0)] reg3144 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3143 = (1'h0);
  reg [(4'he):(1'h0)] reg3142 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3141 = (1'h0);
  reg [(3'h6):(1'h0)] reg3138 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3137 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3135 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3134 = (1'h0);
  reg [(2'h2):(1'h0)] reg3133 = (1'h0);
  reg [(4'he):(1'h0)] reg3130 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3129 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3127 = (1'h0);
  reg [(4'hd):(1'h0)] reg3125 = (1'h0);
  reg [(4'h8):(1'h0)] reg3124 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3123 = (1'h0);
  reg [(4'h9):(1'h0)] reg3122 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3121 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3120 = (1'h0);
  reg [(4'hd):(1'h0)] reg3118 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3117 = (1'h0);
  reg [(3'h7):(1'h0)] reg3116 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3115 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3114 = (1'h0);
  reg [(3'h7):(1'h0)] reg3113 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3112 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3111 = (1'h0);
  reg [(3'h6):(1'h0)] reg3110 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3090 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3086 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3084 = (1'h0);
  reg [(4'hd):(1'h0)] reg3083 = (1'h0);
  reg [(2'h3):(1'h0)] reg3109 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3108 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3107 = (1'h0);
  reg [(3'h7):(1'h0)] reg3106 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3105 = (1'h0);
  reg [(4'he):(1'h0)] reg3104 = (1'h0);
  reg [(4'hd):(1'h0)] reg3093 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3103 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3102 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3101 = (1'h0);
  reg [(5'h10):(1'h0)] reg3100 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3099 = (1'h0);
  reg [(2'h3):(1'h0)] reg3098 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3097 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3096 = (1'h0);
  reg [(4'ha):(1'h0)] reg3095 = (1'h0);
  reg [(4'h8):(1'h0)] reg3094 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3092 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3091 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3089 = (1'h0);
  reg [(4'h8):(1'h0)] reg3088 = (1'h0);
  reg [(4'hb):(1'h0)] reg3087 = (1'h0);
  reg [(3'h6):(1'h0)] reg3085 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3082 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3081 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3080 = (1'h0);
  reg [(3'h6):(1'h0)] reg3079 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3078 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3076 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3075 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3074 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3073 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3071 = (1'h0);
  reg [(4'hc):(1'h0)] reg3070 = (1'h0);
  reg [(2'h3):(1'h0)] reg3069 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3065 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3380 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3376 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3367 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3363 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3361 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3360 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3358 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3357 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3352 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3348 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3347 = (1'h0);
  reg [(4'he):(1'h0)] forvar3344 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3340 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3326 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3321 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3318 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3334 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3330 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3323 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3314 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3312 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3303 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3293 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3292 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3291 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3278 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3276 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3286 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3283 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3277 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3273 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3272 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3284 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3280 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3275 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3274 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3265 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3264 = (1'h0);
  reg [(4'he):(1'h0)] forvar3258 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3256 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3257 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3260 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3255 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3252 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3251 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3242 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3243 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3231 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3228 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3224 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3236 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3233 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3232 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3227 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3225 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3223 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3222 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3213 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3208 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3209 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3205 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3192 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3188 = (1'h0);
  reg [(4'he):(1'h0)] forvar3180 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3179 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3178 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3167 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3164 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3162 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3156 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3151 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3146 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3140 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3139 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3136 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3132 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3131 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3128 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3126 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3119 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3108 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3107 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3106 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3096 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3094 = (1'h0);
  reg [(4'he):(1'h0)] forvar3087 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3098 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3097 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3089 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3100 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3103 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3099 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3093 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3090 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3086 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3084 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3083 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3077 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3072 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3068 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3067 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3066 = (1'h0);
  assign y = {wire3271,
                 wire3270,
                 wire3269,
                 wire3268,
                 wire3267,
                 wire3177,
                 wire3176,
                 wire3175,
                 wire3174,
                 wire3173,
                 wire3064,
                 wire3063,
                 wire3062,
                 wire3061,
                 reg3384,
                 reg3383,
                 reg3382,
                 reg3381,
                 reg3379,
                 reg3378,
                 reg3377,
                 reg3375,
                 reg3374,
                 reg3373,
                 reg3372,
                 reg3371,
                 reg3370,
                 reg3369,
                 reg3368,
                 reg3366,
                 reg3365,
                 reg3364,
                 reg3362,
                 reg3352,
                 reg3359,
                 reg3356,
                 reg3355,
                 reg3354,
                 reg3353,
                 reg3351,
                 reg3350,
                 reg3349,
                 reg3348,
                 reg3346,
                 reg3345,
                 reg3340,
                 reg3344,
                 reg3343,
                 reg3342,
                 reg3341,
                 reg3323,
                 reg3339,
                 reg3334,
                 reg3338,
                 reg3337,
                 reg3336,
                 reg3335,
                 reg3333,
                 reg3332,
                 reg3331,
                 reg3329,
                 reg3328,
                 reg3327,
                 reg3326,
                 reg3325,
                 reg3324,
                 reg3322,
                 reg3321,
                 reg3320,
                 reg3319,
                 reg3318,
                 reg3317,
                 reg3316,
                 reg3315,
                 reg3313,
                 reg3311,
                 reg3310,
                 reg3309,
                 reg3308,
                 reg3307,
                 reg3306,
                 reg3305,
                 reg3304,
                 reg3302,
                 reg3301,
                 reg3300,
                 reg3299,
                 reg3298,
                 reg3297,
                 reg3296,
                 reg3295,
                 reg3294,
                 reg3290,
                 reg3289,
                 reg3288,
                 reg3287,
                 reg3284,
                 reg3280,
                 reg3275,
                 reg3274,
                 reg3286,
                 reg3285,
                 reg3283,
                 reg3282,
                 reg3281,
                 reg3279,
                 reg3278,
                 reg3277,
                 reg3276,
                 reg3273,
                 reg3272,
                 reg3266,
                 reg3263,
                 reg3255,
                 reg3262,
                 reg3260,
                 reg3261,
                 reg3259,
                 reg3258,
                 reg3257,
                 reg3256,
                 reg3254,
                 reg3253,
                 reg3250,
                 reg3249,
                 reg3243,
                 reg3248,
                 reg3247,
                 reg3246,
                 reg3245,
                 reg3244,
                 reg3242,
                 reg3233,
                 reg3232,
                 reg3227,
                 reg3225,
                 reg3241,
                 reg3240,
                 reg3239,
                 reg3238,
                 reg3237,
                 reg3235,
                 reg3234,
                 reg3231,
                 reg3230,
                 reg3229,
                 reg3228,
                 reg3226,
                 reg3224,
                 reg3221,
                 reg3220,
                 reg3219,
                 reg3218,
                 reg3217,
                 reg3216,
                 reg3215,
                 reg3209,
                 reg3214,
                 reg3213,
                 reg3212,
                 reg3211,
                 reg3210,
                 reg3208,
                 reg3207,
                 reg3206,
                 reg3204,
                 reg3203,
                 reg3202,
                 reg3201,
                 reg3200,
                 reg3199,
                 reg3198,
                 reg3197,
                 reg3196,
                 reg3195,
                 reg3194,
                 reg3193,
                 reg3191,
                 reg3190,
                 reg3189,
                 reg3187,
                 reg3186,
                 reg3185,
                 reg3184,
                 reg3183,
                 reg3182,
                 reg3181,
                 reg3172,
                 reg3171,
                 reg3170,
                 reg3169,
                 reg3168,
                 reg3166,
                 reg3165,
                 reg3163,
                 reg3161,
                 reg3160,
                 reg3159,
                 reg3158,
                 reg3157,
                 reg3155,
                 reg3154,
                 reg3153,
                 reg3152,
                 reg3150,
                 reg3149,
                 reg3148,
                 reg3147,
                 reg3145,
                 reg3144,
                 reg3143,
                 reg3142,
                 reg3141,
                 reg3138,
                 reg3137,
                 reg3135,
                 reg3134,
                 reg3133,
                 reg3130,
                 reg3129,
                 reg3127,
                 reg3125,
                 reg3124,
                 reg3123,
                 reg3122,
                 reg3121,
                 reg3120,
                 reg3118,
                 reg3117,
                 reg3116,
                 reg3115,
                 reg3114,
                 reg3113,
                 reg3112,
                 reg3111,
                 reg3110,
                 reg3090,
                 reg3086,
                 reg3084,
                 reg3083,
                 reg3109,
                 reg3108,
                 reg3107,
                 reg3106,
                 reg3105,
                 reg3104,
                 reg3093,
                 reg3103,
                 reg3102,
                 reg3101,
                 reg3100,
                 reg3099,
                 reg3098,
                 reg3097,
                 reg3096,
                 reg3095,
                 reg3094,
                 reg3092,
                 reg3091,
                 reg3089,
                 reg3088,
                 reg3087,
                 reg3085,
                 reg3082,
                 reg3081,
                 reg3080,
                 reg3079,
                 reg3078,
                 reg3076,
                 reg3075,
                 reg3074,
                 reg3073,
                 reg3071,
                 reg3070,
                 reg3069,
                 reg3065,
                 forvar3380,
                 forvar3376,
                 forvar3367,
                 forvar3363,
                 forvar3361,
                 forvar3360,
                 forvar3358,
                 forvar3357,
                 forvar3352,
                 forvar3348,
                 forvar3347,
                 forvar3344,
                 forvar3340,
                 forvar3326,
                 forvar3321,
                 forvar3318,
                 forvar3334,
                 forvar3330,
                 forvar3323,
                 forvar3314,
                 forvar3312,
                 forvar3303,
                 forvar3293,
                 forvar3292,
                 forvar3291,
                 forvar3278,
                 forvar3276,
                 forvar3286,
                 forvar3283,
                 forvar3277,
                 forvar3273,
                 forvar3272,
                 forvar3284,
                 forvar3280,
                 forvar3275,
                 forvar3274,
                 forvar3265,
                 forvar3264,
                 forvar3258,
                 forvar3256,
                 forvar3257,
                 forvar3260,
                 forvar3255,
                 forvar3252,
                 forvar3251,
                 forvar3242,
                 forvar3243,
                 forvar3231,
                 forvar3228,
                 forvar3224,
                 forvar3236,
                 forvar3233,
                 forvar3232,
                 forvar3227,
                 forvar3225,
                 forvar3223,
                 forvar3222,
                 forvar3213,
                 forvar3208,
                 forvar3209,
                 forvar3205,
                 forvar3192,
                 forvar3188,
                 forvar3180,
                 forvar3179,
                 forvar3178,
                 forvar3167,
                 forvar3164,
                 forvar3162,
                 forvar3156,
                 forvar3151,
                 forvar3146,
                 forvar3140,
                 forvar3139,
                 forvar3136,
                 forvar3132,
                 forvar3131,
                 forvar3128,
                 forvar3126,
                 forvar3119,
                 forvar3108,
                 forvar3107,
                 forvar3106,
                 forvar3096,
                 forvar3094,
                 forvar3087,
                 forvar3098,
                 forvar3097,
                 forvar3089,
                 forvar3100,
                 forvar3103,
                 forvar3099,
                 forvar3093,
                 forvar3090,
                 forvar3086,
                 forvar3084,
                 forvar3083,
                 forvar3077,
                 forvar3072,
                 forvar3068,
                 forvar3067,
                 forvar3066,
                 (1'h0)};
  assign wire3061 = wire3058;
  assign wire3062 = $signed($unsigned((wire3057 ^ (wire3061 ?
                        wire3059 : (8'h9c)))));
  assign wire3063 = (wire3059[(3'h6):(3'h5)] != (8'ha8));
  assign wire3064 = (~&{$signed((&(8'ha2)))});
  always
    @(posedge clk) begin
      reg3065 <= $unsigned(((wire3057[(2'h2):(2'h2)] ?
              {(8'hb7)} : (wire3059 | (8'ha3))) ?
          wire3064 : $signed((wire3061 > wire3059))));
      for (forvar3066 = (1'h0); (forvar3066 < (2'h3)); forvar3066 = (forvar3066 + (1'h1)))
        begin
          for (forvar3067 = (1'h0); (forvar3067 < (1'h0)); forvar3067 = (forvar3067 + (1'h1)))
            begin
              for (forvar3068 = (1'h0); (forvar3068 < (1'h0)); forvar3068 = (forvar3068 + (1'h1)))
                begin
                  if ((~^{$signed($signed(wire3061))}))
                    begin
                      reg3069 <= $signed(reg3065[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg3069 <= (-$signed(((wire3058 ? forvar3067 : wire3058) ?
                          (reg3069 && forvar3068) : forvar3067[(3'h5):(2'h3)])));
                      reg3070 <= wire3059[(2'h3):(2'h3)];
                      reg3071 <= forvar3066;
                    end
                end
              if (wire3061[(3'h5):(1'h0)])
                begin
                  for (forvar3072 = (1'h0); (forvar3072 < (2'h3)); forvar3072 = (forvar3072 + (1'h1)))
                    begin
                      reg3073 <= {(~&$unsigned({wire3061}))};
                      reg3074 <= wire3063[(3'h4):(2'h3)];
                      reg3075 <= reg3070[(4'ha):(1'h0)];
                      reg3076 <= $signed(reg3073);
                    end
                  for (forvar3077 = (1'h0); (forvar3077 < (2'h2)); forvar3077 = (forvar3077 + (1'h1)))
                    begin
                      reg3078 <= (8'hba);
                      reg3079 <= $signed((((forvar3077 ?
                              reg3075 : (8'ha1)) < (wire3058 ?
                              wire3063 : reg3071)) ?
                          reg3078[(4'hb):(2'h2)] : forvar3067[(1'h0):(1'h0)]));
                      reg3080 <= ((8'ha4) ? reg3075 : (~&reg3076));
                    end
                end
              else
                begin
                  for (forvar3072 = (1'h0); (forvar3072 < (1'h0)); forvar3072 = (forvar3072 + (1'h1)))
                    begin
                      reg3073 <= reg3070[(3'h4):(3'h4)];
                      reg3074 <= ({$signed($signed(wire3057))} ?
                          ($unsigned($signed(wire3064)) ?
                              reg3076[(3'h5):(2'h3)] : $signed({forvar3067})) : ($unsigned(wire3059) ?
                              ($unsigned(wire3057) | (!reg3071)) : ({wire3059} ?
                                  $unsigned((8'ha3)) : (~^wire3060))));
                      reg3075 <= $unsigned(reg3065[(2'h2):(1'h0)]);
                      reg3076 <= reg3079[(3'h6):(1'h1)];
                    end
                  for (forvar3077 = (1'h0); (forvar3077 < (1'h1)); forvar3077 = (forvar3077 + (1'h1)))
                    begin
                      reg3078 <= $unsigned($unsigned($unsigned((!reg3070))));
                      reg3079 <= (^{$signed($signed(reg3078))});
                      reg3080 <= (~^wire3062[(2'h3):(2'h2)]);
                      reg3081 <= wire3061;
                    end
                end
            end
          reg3082 <= (8'ha6);
        end
      if (($unsigned((^~wire3061)) ?
          $unsigned(reg3078) : ($unsigned($signed(wire3062)) <<< (forvar3067[(2'h3):(1'h0)] ?
              $signed((8'hb2)) : (~&reg3065)))))
        begin
          for (forvar3083 = (1'h0); (forvar3083 < (1'h0)); forvar3083 = (forvar3083 + (1'h1)))
            begin
              for (forvar3084 = (1'h0); (forvar3084 < (2'h2)); forvar3084 = (forvar3084 + (1'h1)))
                begin
                  reg3085 <= (^~(((^reg3071) & wire3058) ?
                      (~&reg3070[(1'h1):(1'h0)]) : reg3073));
                  for (forvar3086 = (1'h0); (forvar3086 < (1'h0)); forvar3086 = (forvar3086 + (1'h1)))
                    begin
                      reg3087 <= (({$unsigned((8'ha5))} < wire3063[(1'h1):(1'h0)]) ?
                          ({$signed(forvar3084)} || (forvar3067[(4'he):(4'ha)] & $signed(reg3069))) : $unsigned((reg3074 >> $signed(reg3079))));
                      reg3088 <= (|(!reg3081[(4'hb):(2'h2)]));
                      reg3089 <= {$signed((8'ha6))};
                    end
                  for (forvar3090 = (1'h0); (forvar3090 < (1'h0)); forvar3090 = (forvar3090 + (1'h1)))
                    begin
                      reg3091 <= ((+(((8'h9e) << (8'ha4)) ?
                              {wire3062} : forvar3066)) ?
                          wire3063[(3'h5):(3'h4)] : ((^(reg3074 ~^ reg3073)) | ($unsigned((8'hb7)) != wire3057[(3'h7):(3'h6)])));
                      reg3092 <= forvar3083[(1'h0):(1'h0)];
                    end
                end
            end
          if ($signed($signed((~^(^~forvar3086)))))
            begin
              for (forvar3093 = (1'h0); (forvar3093 < (1'h1)); forvar3093 = (forvar3093 + (1'h1)))
                begin
                  if ($signed(reg3065[(3'h6):(3'h4)]))
                    begin
                      reg3094 <= $unsigned((~^reg3069[(1'h0):(1'h0)]));
                      reg3095 <= forvar3083;
                      reg3096 <= (wire3063 ^~ forvar3084[(2'h2):(1'h1)]);
                      reg3097 <= reg3079[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg3094 <= {$unsigned(((reg3095 && reg3080) <= reg3065))};
                      reg3095 <= $unsigned((+($signed(reg3080) ?
                          forvar3084[(2'h2):(2'h2)] : (~|forvar3072))));
                      reg3096 <= reg3076[(1'h1):(1'h0)];
                      reg3097 <= $unsigned($signed({(^(8'hb2))}));
                    end
                  reg3098 <= reg3096[(2'h3):(2'h3)];
                  if ((({reg3076[(3'h5):(3'h5)]} * reg3065) ?
                      $unsigned({(reg3074 ?
                              wire3062 : reg3070)}) : $unsigned(forvar3090)))
                    begin
                      reg3099 <= ((($signed(forvar3067) + $signed((8'hb4))) || $unsigned((!forvar3067))) && (~&reg3082));
                      reg3100 <= ($signed($signed($unsigned(reg3073))) ~^ reg3094);
                      reg3101 <= wire3058[(4'hb):(2'h2)];
                      reg3102 <= ($unsigned((~(forvar3066 ?
                          reg3094 : reg3073))) < $unsigned((^(~wire3058))));
                    end
                  else
                    begin
                      reg3099 <= (reg3073 ?
                          (reg3095 != reg3070[(4'hb):(4'h9)]) : (reg3085[(2'h3):(2'h2)] >= reg3078));
                    end
                end
              reg3103 <= {(8'h9c)};
            end
          else
            begin
              reg3093 <= $unsigned($signed($signed($signed(reg3076))));
              reg3094 <= (^~(&(^~reg3103)));
              reg3095 <= $unsigned((&$signed(((8'hac) ?
                  reg3093 : forvar3084))));
              if (reg3070[(3'h7):(2'h2)])
                begin
                  if ($signed((reg3082 & $unsigned($signed(wire3059)))))
                    begin
                      reg3096 <= ($unsigned($signed((forvar3067 ?
                          reg3088 : reg3095))) < ($signed((&forvar3093)) ?
                          ({wire3060} ?
                              {wire3057} : $unsigned(reg3088)) : reg3079));
                    end
                  else
                    begin
                      reg3096 <= reg3085;
                      reg3097 <= wire3059[(3'h6):(1'h0)];
                      reg3098 <= {(reg3079[(3'h4):(1'h1)] ?
                              $unsigned({(8'hb5)}) : forvar3068[(2'h2):(1'h0)])};
                    end
                  for (forvar3099 = (1'h0); (forvar3099 < (2'h3)); forvar3099 = (forvar3099 + (1'h1)))
                    begin
                      reg3100 <= ((|forvar3077) ?
                          $unsigned(reg3076[(3'h5):(3'h5)]) : $unsigned(reg3081[(4'hb):(3'h4)]));
                      reg3101 <= $signed(((forvar3068[(2'h3):(2'h2)] * (~^reg3080)) ?
                          $signed(reg3079) : $unsigned(reg3102[(1'h1):(1'h0)])));
                      reg3102 <= $signed($signed($unsigned(((8'hb4) ?
                          reg3069 : forvar3093))));
                    end
                  for (forvar3103 = (1'h0); (forvar3103 < (2'h2)); forvar3103 = (forvar3103 + (1'h1)))
                    begin
                      reg3104 <= reg3065;
                      reg3105 <= (8'hb0);
                    end
                  if ($unsigned(reg3085))
                    begin
                      reg3106 <= (^reg3101);
                      reg3107 <= $signed((wire3057[(3'h7):(3'h4)] ?
                          ($signed(reg3093) ?
                              reg3105 : $signed(wire3059)) : ((~&reg3074) ?
                              $unsigned(forvar3067) : {forvar3099})));
                      reg3108 <= ($unsigned({$unsigned(reg3076)}) ?
                          reg3091[(2'h3):(2'h2)] : (~$unsigned($unsigned(reg3088))));
                      reg3109 <= reg3082;
                    end
                  else
                    begin
                      reg3106 <= (~^reg3092[(4'h8):(3'h6)]);
                    end
                end
              else
                begin
                  if (((+($signed((8'hba)) ?
                      {(8'had)} : (forvar3086 ?
                          forvar3084 : reg3100))) < reg3078[(3'h7):(3'h6)]))
                    begin
                      reg3096 <= $unsigned(((!$signed(reg3091)) >= (((8'ha0) >= reg3104) ?
                          $unsigned(reg3106) : (|(8'ha3)))));
                      reg3097 <= wire3057[(3'h5):(3'h5)];
                      reg3098 <= $signed(({(forvar3090 ? (8'hb1) : reg3089)} ?
                          ($signed(reg3098) ?
                              forvar3066[(1'h0):(1'h0)] : $unsigned(wire3062)) : forvar3072[(3'h6):(2'h2)]));
                      reg3099 <= (($signed({reg3098}) ?
                          forvar3066[(2'h2):(1'h0)] : (~|reg3082)) | {(-forvar3093)});
                    end
                  else
                    begin
                      reg3096 <= {reg3102};
                    end
                  for (forvar3100 = (1'h0); (forvar3100 < (2'h2)); forvar3100 = (forvar3100 + (1'h1)))
                    begin
                      reg3101 <= (!forvar3084[(3'h7):(3'h4)]);
                      reg3102 <= (|($signed(reg3087[(3'h6):(2'h3)]) ?
                          wire3059[(3'h4):(3'h4)] : (+forvar3084)));
                      reg3103 <= (!$unsigned((8'hb8)));
                      reg3104 <= reg3078[(1'h0):(1'h0)];
                    end
                  if ((reg3065 ? forvar3086 : $unsigned((8'ha0))))
                    begin
                      reg3105 <= reg3093;
                    end
                  else
                    begin
                      reg3105 <= reg3085[(3'h5):(1'h1)];
                      reg3106 <= ((forvar3090[(1'h0):(1'h0)] ?
                          $unsigned((reg3094 || wire3063)) : ((8'hac) ?
                              (forvar3083 ?
                                  forvar3100 : reg3099) : (forvar3084 ?
                                  wire3058 : wire3058))) + $unsigned(reg3107[(2'h2):(1'h1)]));
                      reg3107 <= ((&(8'hba)) >= {$signed($signed(reg3079))});
                      reg3108 <= (reg3087[(3'h4):(2'h3)] | ((&$signed(reg3081)) ?
                          (!(forvar3067 && reg3094)) : (~^forvar3077[(2'h2):(1'h0)])));
                    end
                end
            end
        end
      else
        begin
          if ($signed((~|(~reg3082[(2'h3):(2'h2)]))))
            begin
              if (reg3104[(4'he):(3'h4)])
                begin
                  if (($signed($unsigned($signed(wire3062))) ?
                      ((8'ha4) ?
                          reg3100[(3'h6):(2'h3)] : reg3092[(4'he):(1'h1)]) : reg3101[(3'h5):(2'h3)]))
                    begin
                      reg3083 <= {reg3095};
                    end
                  else
                    begin
                      reg3083 <= $signed((-forvar3067));
                      reg3084 <= ((^($unsigned(reg3065) ?
                          {reg3106} : (&reg3089))) >> reg3091);
                      reg3085 <= ($signed(reg3102[(1'h0):(1'h0)]) ?
                          reg3092[(3'h5):(1'h1)] : reg3096[(3'h5):(3'h4)]);
                      reg3086 <= (8'h9f);
                    end
                  if (((reg3095 ?
                      forvar3066 : forvar3067[(4'hb):(3'h6)]) < reg3107))
                    begin
                      reg3087 <= (^{reg3086});
                    end
                  else
                    begin
                      reg3087 <= (|((~(~^reg3094)) ?
                          $signed($signed(forvar3068)) : ($unsigned((8'ha4)) ?
                              $unsigned(reg3108) : (wire3062 ?
                                  forvar3084 : reg3087))));
                      reg3088 <= forvar3083;
                    end
                  for (forvar3089 = (1'h0); (forvar3089 < (2'h3)); forvar3089 = (forvar3089 + (1'h1)))
                    begin
                      reg3090 <= reg3074[(2'h3):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar3083 = (1'h0); (forvar3083 < (2'h3)); forvar3083 = (forvar3083 + (1'h1)))
                    begin
                      reg3084 <= (^(-(((8'hb0) >> (8'hb0)) ?
                          reg3108[(1'h1):(1'h0)] : $signed((8'ha6)))));
                      reg3085 <= forvar3083[(1'h1):(1'h0)];
                      reg3086 <= reg3096;
                    end
                  if (reg3074[(1'h0):(1'h0)])
                    begin
                      reg3087 <= $signed(({reg3094} + (((8'haf) <<< reg3091) == ((8'hb6) ?
                          forvar3100 : reg3065))));
                      reg3088 <= (~reg3098);
                      reg3089 <= ($signed($unsigned({forvar3077})) ?
                          ($signed({reg3096}) ^~ ({(8'ha2)} ?
                              {wire3058} : {reg3092})) : (reg3083[(3'h5):(2'h2)] < reg3095[(3'h6):(1'h1)]));
                      reg3090 <= reg3079[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3087 <= $signed(reg3080[(4'ha):(3'h7)]);
                      reg3088 <= (reg3089 ?
                          {$unsigned($signed(wire3057))} : $unsigned(forvar3077[(2'h2):(2'h2)]));
                      reg3089 <= (forvar3103[(4'h8):(4'h8)] <<< $unsigned((~&(wire3061 - wire3061))));
                    end
                  if ($signed((({wire3064} - forvar3099[(1'h1):(1'h0)]) & $signed(reg3087[(2'h2):(1'h1)]))))
                    begin
                      reg3091 <= $signed(reg3082);
                    end
                  else
                    begin
                      reg3091 <= wire3061;
                      reg3092 <= (((8'ha1) | $unsigned((^~reg3101))) == reg3087);
                      reg3093 <= (8'hb5);
                      reg3094 <= wire3064;
                    end
                  if ((&$signed((~{reg3102}))))
                    begin
                      reg3095 <= (+(^reg3086));
                    end
                  else
                    begin
                      reg3095 <= {reg3093[(3'h4):(3'h4)]};
                      reg3096 <= {$signed((|(reg3069 != reg3101)))};
                    end
                end
              for (forvar3097 = (1'h0); (forvar3097 < (2'h2)); forvar3097 = (forvar3097 + (1'h1)))
                begin
                  for (forvar3098 = (1'h0); (forvar3098 < (1'h0)); forvar3098 = (forvar3098 + (1'h1)))
                    begin
                      reg3099 <= forvar3086;
                      reg3100 <= $signed(({$signed(reg3076)} * (~|(&reg3076))));
                      reg3101 <= reg3092[(4'hc):(3'h5)];
                      reg3102 <= (reg3106[(2'h3):(1'h0)] * $signed(((~|reg3080) - reg3070[(2'h2):(2'h2)])));
                    end
                  for (forvar3103 = (1'h0); (forvar3103 < (1'h0)); forvar3103 = (forvar3103 + (1'h1)))
                    begin
                      reg3104 <= (forvar3103[(4'h9):(3'h5)] ?
                          (wire3061[(3'h6):(2'h3)] ?
                              (-$unsigned(reg3084)) : $unsigned({reg3092})) : reg3074[(2'h2):(1'h0)]);
                    end
                  reg3105 <= reg3075[(4'h8):(2'h2)];
                end
            end
          else
            begin
              if (reg3080[(2'h2):(2'h2)])
                begin
                  if (($unsigned((~^$unsigned(forvar3083))) && $unsigned((8'hb8))))
                    begin
                      reg3083 <= ($unsigned({(reg3098 - reg3085)}) ?
                          wire3061 : forvar3067);
                    end
                  else
                    begin
                      reg3083 <= $unsigned((((forvar3097 ? (8'ha5) : wire3063) ?
                              (8'hba) : reg3085[(2'h3):(2'h3)]) ?
                          (8'ha2) : reg3082));
                      reg3084 <= $unsigned({((reg3092 ? reg3102 : reg3104) ?
                              $unsigned(wire3060) : ((8'haf) ?
                                  wire3063 : wire3062))});
                      reg3085 <= {(8'ha9)};
                    end
                  for (forvar3086 = (1'h0); (forvar3086 < (1'h1)); forvar3086 = (forvar3086 + (1'h1)))
                    begin
                      reg3087 <= ((8'hae) >= $unsigned(($unsigned(reg3073) ?
                          (&reg3094) : $unsigned(forvar3089))));
                      reg3088 <= reg3089;
                      reg3089 <= $unsigned(reg3105[(4'hc):(1'h1)]);
                    end
                  if (reg3101)
                    begin
                      reg3090 <= ((+($unsigned((8'ha7)) ?
                              ((8'hb8) ~^ reg3104) : (8'ha3))) ?
                          {reg3108[(4'h8):(4'h8)]} : reg3103[(3'h5):(2'h2)]);
                      reg3091 <= $unsigned($unsigned((-(reg3095 ?
                          (8'hb2) : (8'hb7)))));
                    end
                  else
                    begin
                      reg3090 <= ($unsigned(((reg3082 & wire3059) >>> $signed(reg3104))) <= wire3064);
                      reg3091 <= $unsigned((8'hb4));
                      reg3092 <= $unsigned(($signed((~&forvar3084)) > $unsigned(reg3092)));
                      reg3093 <= {reg3094[(1'h1):(1'h1)]};
                    end
                end
              else
                begin
                  if (((forvar3093[(3'h6):(3'h4)] ?
                      ((reg3097 >= (8'hb2)) || reg3076[(3'h6):(1'h1)]) : $unsigned(reg3099[(1'h1):(1'h1)])) << $signed(($unsigned(reg3094) ?
                      (^~reg3108) : reg3071))))
                    begin
                      reg3083 <= forvar3093[(1'h1):(1'h0)];
                      reg3084 <= forvar3086;
                    end
                  else
                    begin
                      reg3083 <= forvar3067;
                      reg3084 <= {($unsigned((+reg3078)) ?
                              reg3095[(3'h5):(3'h5)] : $unsigned(((8'hb4) | forvar3090)))};
                    end
                  reg3085 <= $unsigned($unsigned((reg3109[(2'h3):(2'h3)] ?
                      (|reg3095) : $unsigned(reg3100))));
                  reg3086 <= $unsigned(($unsigned(forvar3084) - $unsigned($unsigned((8'ha4)))));
                  for (forvar3087 = (1'h0); (forvar3087 < (1'h1)); forvar3087 = (forvar3087 + (1'h1)))
                    begin
                      reg3088 <= reg3091;
                      reg3089 <= (((^~reg3069) <= (forvar3087[(4'hb):(2'h2)] ?
                          reg3100 : {forvar3072})) & $unsigned($unsigned(forvar3098[(2'h2):(1'h0)])));
                    end
                end
              for (forvar3094 = (1'h0); (forvar3094 < (1'h0)); forvar3094 = (forvar3094 + (1'h1)))
                begin
                  reg3095 <= (forvar3066[(1'h0):(1'h0)] >>> reg3073[(2'h2):(1'h1)]);
                  for (forvar3096 = (1'h0); (forvar3096 < (2'h3)); forvar3096 = (forvar3096 + (1'h1)))
                    begin
                      reg3097 <= (!$signed($unsigned((^~wire3057))));
                    end
                end
              for (forvar3098 = (1'h0); (forvar3098 < (2'h2)); forvar3098 = (forvar3098 + (1'h1)))
                begin
                  reg3099 <= reg3106;
                end
            end
          for (forvar3106 = (1'h0); (forvar3106 < (1'h1)); forvar3106 = (forvar3106 + (1'h1)))
            begin
              for (forvar3107 = (1'h0); (forvar3107 < (1'h0)); forvar3107 = (forvar3107 + (1'h1)))
                begin
                  for (forvar3108 = (1'h0); (forvar3108 < (2'h3)); forvar3108 = (forvar3108 + (1'h1)))
                    begin
                      reg3109 <= $signed(($unsigned((forvar3106 ?
                          reg3080 : reg3081)) > (reg3070[(3'h7):(3'h4)] * $signed((8'hb6)))));
                      reg3110 <= reg3103[(3'h6):(3'h6)];
                      reg3111 <= ($unsigned(forvar3089) | {reg3085});
                      reg3112 <= ((~|forvar3098) <<< (forvar3067[(2'h3):(1'h1)] && (!$signed(wire3058))));
                    end
                  reg3113 <= (+(8'ha1));
                  if ({reg3070[(3'h7):(3'h5)]})
                    begin
                      reg3114 <= ((((reg3086 >= (8'hba)) ?
                              (forvar3093 & reg3082) : (&forvar3068)) ~^ ((forvar3067 > reg3093) * {reg3078})) ?
                          (wire3059[(1'h0):(1'h0)] << (reg3084[(2'h3):(1'h1)] | (forvar3094 ?
                              forvar3093 : wire3060))) : reg3087[(1'h0):(1'h0)]);
                      reg3115 <= wire3062;
                      reg3116 <= (($unsigned(reg3100) * $unsigned((reg3080 * reg3070))) ?
                          $unsigned(($unsigned((8'hac)) ~^ $unsigned(wire3061))) : {reg3080});
                      reg3117 <= (reg3088[(3'h4):(1'h1)] ?
                          (~|(8'ha6)) : (8'ha0));
                    end
                  else
                    begin
                      reg3114 <= (~^(forvar3077[(2'h2):(1'h0)] < $unsigned(reg3108[(2'h2):(1'h0)])));
                      reg3115 <= $signed((reg3109[(1'h0):(1'h0)] & (reg3096[(2'h3):(2'h2)] & {forvar3087})));
                      reg3116 <= $signed($signed($signed((~&reg3071))));
                    end
                end
              reg3118 <= forvar3066[(2'h2):(2'h2)];
              for (forvar3119 = (1'h0); (forvar3119 < (1'h1)); forvar3119 = (forvar3119 + (1'h1)))
                begin
                  if (forvar3087)
                    begin
                      reg3120 <= (+{reg3073});
                      reg3121 <= ({($unsigned(reg3086) & reg3075[(3'h7):(3'h7)])} - $signed($unsigned((~&forvar3068))));
                    end
                  else
                    begin
                      reg3120 <= reg3106[(2'h3):(2'h2)];
                      reg3121 <= (reg3092[(3'h5):(1'h1)] ~^ $unsigned((8'hab)));
                      reg3122 <= ($signed($signed((reg3096 ?
                              wire3058 : wire3061))) ?
                          $unsigned($signed((^~reg3110))) : {$signed((8'ha8))});
                      reg3123 <= ((&{wire3064}) <= $signed($unsigned($unsigned((8'hb6)))));
                    end
                  reg3124 <= reg3121;
                  reg3125 <= reg3073[(3'h4):(2'h3)];
                  for (forvar3126 = (1'h0); (forvar3126 < (2'h2)); forvar3126 = (forvar3126 + (1'h1)))
                    begin
                      reg3127 <= forvar3126[(1'h1):(1'h0)];
                    end
                end
            end
          for (forvar3128 = (1'h0); (forvar3128 < (2'h2)); forvar3128 = (forvar3128 + (1'h1)))
            begin
              reg3129 <= (+((~|$unsigned(reg3102)) <= ((8'hae) == $signed(reg3112))));
              reg3130 <= ($unsigned((|reg3101)) ?
                  wire3062[(1'h1):(1'h0)] : wire3064[(4'h8):(2'h3)]);
            end
          for (forvar3131 = (1'h0); (forvar3131 < (2'h2)); forvar3131 = (forvar3131 + (1'h1)))
            begin
              for (forvar3132 = (1'h0); (forvar3132 < (2'h3)); forvar3132 = (forvar3132 + (1'h1)))
                begin
                  if ((8'h9c))
                    begin
                      reg3133 <= $signed($unsigned((8'ha9)));
                      reg3134 <= $unsigned((^((reg3105 & forvar3083) ?
                          (reg3075 ? reg3078 : (8'hb3)) : (8'hb2))));
                      reg3135 <= $signed($signed((((8'haa) | reg3065) && $unsigned(reg3082))));
                    end
                  else
                    begin
                      reg3133 <= ((reg3074[(2'h2):(2'h2)] & ((&(8'ha4)) ?
                              ((8'hac) <<< reg3130) : ((8'h9f) ?
                                  reg3133 : reg3065))) ?
                          ($signed((!reg3111)) >> ((8'h9e) ?
                              (8'ha0) : $unsigned((8'ha3)))) : forvar3100[(2'h2):(1'h0)]);
                      reg3134 <= $unsigned({$signed(reg3084)});
                      reg3135 <= $unsigned($unsigned((8'ha0)));
                    end
                  for (forvar3136 = (1'h0); (forvar3136 < (1'h0)); forvar3136 = (forvar3136 + (1'h1)))
                    begin
                      reg3137 <= reg3070[(4'h8):(2'h3)];
                      reg3138 <= (($unsigned((~^wire3060)) ?
                          $unsigned(reg3065) : {(forvar3093 ?
                                  (8'hb9) : wire3061)}) & reg3081);
                    end
                end
              for (forvar3139 = (1'h0); (forvar3139 < (2'h2)); forvar3139 = (forvar3139 + (1'h1)))
                begin
                  for (forvar3140 = (1'h0); (forvar3140 < (2'h2)); forvar3140 = (forvar3140 + (1'h1)))
                    begin
                      reg3141 <= ($signed(($unsigned(wire3058) ?
                          ((8'ha9) == reg3086) : (reg3093 >> reg3103))) ^ ({wire3058} ?
                          {(8'h9e)} : forvar3072[(3'h6):(2'h3)]));
                      reg3142 <= reg3115[(1'h0):(1'h0)];
                      reg3143 <= {reg3137};
                      reg3144 <= (reg3096[(2'h3):(2'h3)] << $unsigned({(reg3110 || reg3088)}));
                    end
                  reg3145 <= $unsigned((forvar3067[(3'h6):(3'h5)] ?
                      wire3059[(1'h1):(1'h1)] : $signed((+forvar3108))));
                  for (forvar3146 = (1'h0); (forvar3146 < (1'h0)); forvar3146 = (forvar3146 + (1'h1)))
                    begin
                      reg3147 <= $unsigned((-$signed((8'hba))));
                      reg3148 <= ((forvar3103 && $unsigned((reg3117 ?
                              reg3100 : reg3133))) ?
                          ($signed((|reg3080)) >>> (~|(~|reg3135))) : reg3109);
                      reg3149 <= $signed({$unsigned(wire3060[(3'h4):(3'h4)])});
                      reg3150 <= reg3100[(3'h5):(3'h5)];
                    end
                  for (forvar3151 = (1'h0); (forvar3151 < (2'h3)); forvar3151 = (forvar3151 + (1'h1)))
                    begin
                      reg3152 <= reg3102;
                      reg3153 <= $signed($unsigned((^(reg3118 ~^ reg3087))));
                      reg3154 <= $unsigned($unsigned((^~$signed(reg3082))));
                      reg3155 <= (-$unsigned(reg3114));
                    end
                end
              for (forvar3156 = (1'h0); (forvar3156 < (2'h3)); forvar3156 = (forvar3156 + (1'h1)))
                begin
                  reg3157 <= (~forvar3131);
                  if (reg3079)
                    begin
                      reg3158 <= forvar3126[(4'h9):(3'h4)];
                      reg3159 <= ($unsigned((!reg3127[(1'h0):(1'h0)])) | reg3137);
                      reg3160 <= (^~reg3116[(3'h4):(1'h0)]);
                      reg3161 <= (8'ha8);
                    end
                  else
                    begin
                      reg3158 <= (|$unsigned($signed($unsigned(reg3149))));
                    end
                end
              for (forvar3162 = (1'h0); (forvar3162 < (1'h1)); forvar3162 = (forvar3162 + (1'h1)))
                begin
                  reg3163 <= ((((!reg3158) ?
                      forvar3139[(2'h3):(2'h2)] : reg3071) <= (~|$unsigned(reg3159))) - $signed((reg3101 ?
                      $unsigned(reg3111) : $unsigned(reg3087))));
                  for (forvar3164 = (1'h0); (forvar3164 < (1'h0)); forvar3164 = (forvar3164 + (1'h1)))
                    begin
                      reg3165 <= (forvar3089[(3'h6):(1'h1)] ?
                          $unsigned(forvar3103[(4'ha):(1'h1)]) : $signed(($signed((8'ha5)) ?
                              {reg3113} : (forvar3066 ?
                                  forvar3156 : reg3113))));
                      reg3166 <= (|forvar3156[(2'h2):(2'h2)]);
                    end
                  for (forvar3167 = (1'h0); (forvar3167 < (1'h0)); forvar3167 = (forvar3167 + (1'h1)))
                    begin
                      reg3168 <= (^~reg3088[(2'h2):(1'h1)]);
                      reg3169 <= ($unsigned((-$unsigned((8'hae)))) - $signed(forvar3099));
                      reg3170 <= reg3076;
                    end
                  if ((+$signed($signed($signed(reg3116)))))
                    begin
                      reg3171 <= $signed((reg3152[(4'hb):(3'h4)] ?
                          $unsigned((^~forvar3107)) : reg3101[(3'h5):(2'h2)]));
                      reg3172 <= reg3120[(3'h6):(1'h0)];
                    end
                  else
                    begin
                      reg3171 <= $signed(forvar3094[(1'h0):(1'h0)]);
                      reg3172 <= (($unsigned(reg3154[(3'h4):(2'h2)]) >>> ((~forvar3139) == forvar3151[(3'h6):(3'h6)])) ?
                          $signed(($signed(reg3093) ?
                              (+reg3082) : ((8'hb4) ^ forvar3066))) : {reg3129[(1'h1):(1'h1)]});
                    end
                end
            end
        end
    end
  assign wire3173 = ((^~reg3134[(4'hd):(4'h8)]) ^ (reg3086 + $unsigned($unsigned(reg3133))));
  assign wire3174 = (($unsigned((|reg3130)) ?
                        $unsigned({(8'ha4)}) : reg3127) > (reg3087 ?
                        (~|(reg3153 ? wire3064 : reg3080)) : (-(!reg3142))));
  assign wire3175 = (reg3108[(3'h4):(3'h4)] ?
                        (((~&reg3166) ?
                            reg3160 : reg3092[(4'he):(1'h1)]) < $signed($unsigned((8'hba)))) : $unsigned(($unsigned(reg3149) ?
                            {reg3117} : $unsigned(wire3058))));
  assign wire3176 = (({reg3137[(3'h4):(2'h2)]} << ({(8'ha0)} <<< $unsigned(reg3144))) ?
                        (-reg3085) : ($signed($signed(reg3086)) ?
                            reg3168 : reg3152[(4'h9):(4'h9)]));
  assign wire3177 = (reg3081[(4'ha):(1'h0)] ?
                        ($unsigned(reg3084[(3'h6):(1'h1)]) - wire3176[(2'h3):(1'h1)]) : $signed($signed((~&reg3070))));
  always
    @(posedge clk) begin
      for (forvar3178 = (1'h0); (forvar3178 < (1'h1)); forvar3178 = (forvar3178 + (1'h1)))
        begin
          for (forvar3179 = (1'h0); (forvar3179 < (1'h1)); forvar3179 = (forvar3179 + (1'h1)))
            begin
              if (($signed($signed(((8'ha3) ? reg3099 : (8'h9d)))) ?
                  $unsigned(reg3130[(2'h2):(1'h0)]) : $unsigned(reg3137)))
                begin
                  for (forvar3180 = (1'h0); (forvar3180 < (2'h2)); forvar3180 = (forvar3180 + (1'h1)))
                    begin
                      reg3181 <= $signed($unsigned((reg3117[(1'h0):(1'h0)] == reg3133)));
                    end
                end
              else
                begin
                  for (forvar3180 = (1'h0); (forvar3180 < (2'h3)); forvar3180 = (forvar3180 + (1'h1)))
                    begin
                      reg3181 <= (reg3094 > $unsigned(((reg3157 ?
                              reg3098 : reg3155) ?
                          $signed((8'h9d)) : wire3176[(4'h8):(3'h7)])));
                      reg3182 <= $unsigned(reg3138);
                      reg3183 <= (reg3084[(3'h7):(3'h6)] | (~|((reg3129 ?
                          wire3058 : (8'hae)) >>> {reg3121})));
                      reg3184 <= reg3073;
                    end
                  if ((reg3172 ?
                      $unsigned((|$unsigned(reg3087))) : $signed($signed($signed((8'hb7))))))
                    begin
                      reg3185 <= ((wire3061[(3'h5):(2'h3)] ?
                              reg3086 : wire3061) ?
                          (((^~(8'ha7)) >= (~wire3174)) ?
                              reg3070[(4'ha):(4'h8)] : (~|(~reg3134))) : $signed($signed($signed(reg3087))));
                    end
                  else
                    begin
                      reg3185 <= reg3092[(3'h5):(1'h1)];
                      reg3186 <= (($signed({reg3138}) ?
                              $signed($signed(reg3088)) : $signed(((8'ha6) | (8'h9e)))) ?
                          $signed(reg3121) : {$signed($signed(reg3099))});
                      reg3187 <= $unsigned((((!reg3099) >> {reg3124}) ?
                          reg3099[(4'hd):(2'h3)] : (reg3170 ?
                              (reg3069 ?
                                  (8'hb9) : wire3060) : reg3069[(1'h0):(1'h0)])));
                    end
                  for (forvar3188 = (1'h0); (forvar3188 < (1'h0)); forvar3188 = (forvar3188 + (1'h1)))
                    begin
                      reg3189 <= reg3161[(4'ha):(3'h5)];
                      reg3190 <= $unsigned($signed($signed((reg3094 ?
                          wire3175 : reg3134))));
                      reg3191 <= (reg3149[(3'h5):(3'h5)] >> $unsigned((reg3065[(4'h8):(3'h6)] <<< $signed(reg3138))));
                    end
                end
              for (forvar3192 = (1'h0); (forvar3192 < (1'h0)); forvar3192 = (forvar3192 + (1'h1)))
                begin
                  if (reg3081)
                    begin
                      reg3193 <= reg3171;
                      reg3194 <= {{($signed((8'h9d)) ?
                                  forvar3192 : reg3102[(3'h4):(3'h4)])}};
                      reg3195 <= (!$unsigned(reg3149));
                      reg3196 <= ((~^((reg3124 ? reg3082 : (8'hb2)) ?
                              {reg3153} : (reg3124 ? wire3059 : wire3173))) ?
                          reg3185[(1'h1):(1'h1)] : $signed({(reg3194 ?
                                  reg3172 : reg3121)}));
                    end
                  else
                    begin
                      reg3193 <= ($signed((reg3144[(4'hb):(4'hb)] ?
                          (~reg3122) : (~^reg3157))) || (forvar3180 ?
                          reg3149 : $signed(((8'hb9) < reg3142))));
                    end
                  if ($unsigned($signed((&$signed(reg3159)))))
                    begin
                      reg3197 <= $unsigned(reg3134[(2'h3):(2'h2)]);
                      reg3198 <= (^~{((~(8'ha3)) != reg3102[(2'h2):(1'h1)])});
                      reg3199 <= reg3081;
                      reg3200 <= ($signed({$unsigned(reg3142)}) ?
                          (~|reg3135[(2'h3):(2'h3)]) : $unsigned(reg3090[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg3197 <= reg3168;
                      reg3198 <= (|reg3096[(2'h3):(1'h0)]);
                      reg3199 <= reg3185[(3'h4):(3'h4)];
                    end
                  if ({(~|$unsigned(wire3063))})
                    begin
                      reg3201 <= (~&(+$unsigned((reg3098 & reg3105))));
                      reg3202 <= reg3075[(1'h0):(1'h0)];
                      reg3203 <= ((((reg3082 & reg3198) ?
                                  (reg3200 ? reg3106 : wire3059) : {(8'hb5)}) ?
                              ((^reg3163) ~^ (reg3084 ?
                                  reg3149 : reg3083)) : {(reg3085 ?
                                      reg3163 : reg3190)}) ?
                          (($unsigned(reg3154) ?
                              ((8'ha5) ?
                                  reg3105 : forvar3178) : reg3147) - (~(reg3081 - reg3100))) : ($signed($signed(reg3201)) >= {$signed((8'had))}));
                      reg3204 <= $signed($signed((reg3097 <<< $unsigned(reg3155))));
                    end
                  else
                    begin
                      reg3201 <= ((~|$signed((reg3142 ? reg3163 : reg3091))) ?
                          wire3173 : (~(8'hb1)));
                      reg3202 <= $signed(reg3184);
                      reg3203 <= reg3130[(2'h3):(2'h3)];
                      reg3204 <= ($signed((reg3141[(1'h1):(1'h0)] <<< (reg3169 - reg3160))) <<< reg3198);
                    end
                  for (forvar3205 = (1'h0); (forvar3205 < (2'h3)); forvar3205 = (forvar3205 + (1'h1)))
                    begin
                      reg3206 <= reg3098[(2'h2):(1'h1)];
                      reg3207 <= (+(8'ha3));
                    end
                end
              if ((reg3118 << reg3135[(3'h6):(3'h5)]))
                begin
                  reg3208 <= (((reg3202[(1'h0):(1'h0)] ?
                          $signed(reg3124) : reg3203[(2'h2):(1'h0)]) ?
                      $signed($unsigned(reg3137)) : reg3097[(1'h1):(1'h0)]) == $unsigned($signed(reg3070[(4'hc):(2'h3)])));
                  for (forvar3209 = (1'h0); (forvar3209 < (2'h3)); forvar3209 = (forvar3209 + (1'h1)))
                    begin
                      reg3210 <= $unsigned($signed($unsigned((reg3165 ?
                          wire3064 : reg3096))));
                      reg3211 <= {reg3198};
                      reg3212 <= reg3106[(3'h4):(2'h2)];
                    end
                  if ((~^{(reg3212 <= reg3210[(2'h3):(2'h2)])}))
                    begin
                      reg3213 <= ((~reg3071[(3'h6):(1'h1)]) <<< $signed($unsigned(reg3111)));
                    end
                  else
                    begin
                      reg3213 <= reg3207[(3'h6):(2'h3)];
                      reg3214 <= (~|reg3148);
                    end
                end
              else
                begin
                  for (forvar3208 = (1'h0); (forvar3208 < (2'h2)); forvar3208 = (forvar3208 + (1'h1)))
                    begin
                      reg3209 <= $unsigned((($signed(reg3150) ?
                          {reg3114} : $signed(reg3101)) > reg3160));
                      reg3210 <= reg3183[(3'h6):(1'h1)];
                      reg3211 <= $unsigned(reg3209[(1'h1):(1'h1)]);
                      reg3212 <= forvar3208[(3'h4):(2'h2)];
                    end
                  for (forvar3213 = (1'h0); (forvar3213 < (1'h0)); forvar3213 = (forvar3213 + (1'h1)))
                    begin
                      reg3214 <= (reg3147 ? (8'ha8) : reg3100[(2'h2):(1'h1)]);
                      reg3215 <= {$signed($signed(reg3191[(1'h0):(1'h0)]))};
                    end
                end
              if ($signed($unsigned({forvar3192})))
                begin
                  reg3216 <= reg3101;
                  reg3217 <= ($signed($unsigned({reg3181})) != (((reg3143 & (8'hb5)) ?
                          $unsigned(reg3096) : $unsigned(reg3078)) ?
                      $signed((reg3208 ?
                          forvar3213 : reg3149)) : ((~&reg3097) << $signed(reg3117))));
                end
              else
                begin
                  reg3216 <= (^~$unsigned(reg3190[(3'h6):(1'h0)]));
                  if (reg3144[(2'h3):(2'h2)])
                    begin
                      reg3217 <= {reg3155[(2'h3):(1'h0)]};
                      reg3218 <= {reg3196};
                    end
                  else
                    begin
                      reg3217 <= reg3213;
                      reg3218 <= $signed(($unsigned((wire3058 ?
                          (8'h9e) : reg3165)) >= $signed({reg3183})));
                      reg3219 <= {reg3118[(1'h1):(1'h1)]};
                    end
                end
            end
          reg3220 <= $unsigned(reg3098);
          reg3221 <= $signed({(reg3189[(4'h8):(1'h1)] ?
                  $signed(reg3110) : reg3183)});
        end
      for (forvar3222 = (1'h0); (forvar3222 < (1'h1)); forvar3222 = (forvar3222 + (1'h1)))
        begin
          if (reg3091[(3'h6):(1'h1)])
            begin
              for (forvar3223 = (1'h0); (forvar3223 < (1'h1)); forvar3223 = (forvar3223 + (1'h1)))
                begin
                  reg3224 <= $signed(($unsigned(reg3182[(3'h5):(2'h2)]) ?
                      ((reg3214 + reg3138) & (reg3121 <<< reg3065)) : reg3219));
                  for (forvar3225 = (1'h0); (forvar3225 < (2'h2)); forvar3225 = (forvar3225 + (1'h1)))
                    begin
                      reg3226 <= reg3185[(2'h3):(1'h1)];
                    end
                  for (forvar3227 = (1'h0); (forvar3227 < (1'h0)); forvar3227 = (forvar3227 + (1'h1)))
                    begin
                      reg3228 <= reg3102[(1'h0):(1'h0)];
                      reg3229 <= ((reg3096[(3'h4):(1'h0)] ?
                              $unsigned((8'hb5)) : {$signed(reg3161)}) ?
                          ((reg3095[(2'h2):(1'h0)] ? {reg3224} : reg3191) ?
                              ($signed(reg3186) >> (+reg3155)) : (&$unsigned(reg3142))) : $unsigned(($unsigned((8'hb4)) ~^ reg3118)));
                      reg3230 <= (~^wire3063[(3'h5):(2'h2)]);
                      reg3231 <= forvar3209;
                    end
                end
              for (forvar3232 = (1'h0); (forvar3232 < (2'h3)); forvar3232 = (forvar3232 + (1'h1)))
                begin
                  for (forvar3233 = (1'h0); (forvar3233 < (2'h3)); forvar3233 = (forvar3233 + (1'h1)))
                    begin
                      reg3234 <= $unsigned((($unsigned(reg3086) && reg3081) + $signed(reg3165[(2'h2):(1'h0)])));
                      reg3235 <= reg3084;
                    end
                  for (forvar3236 = (1'h0); (forvar3236 < (2'h3)); forvar3236 = (forvar3236 + (1'h1)))
                    begin
                      reg3237 <= {($signed({reg3125}) >> $unsigned(reg3163[(1'h1):(1'h0)]))};
                      reg3238 <= $signed((^~(wire3176 ?
                          {forvar3223} : (reg3082 ? reg3109 : (8'hb0)))));
                      reg3239 <= $signed(reg3090[(1'h0):(1'h0)]);
                      reg3240 <= reg3073;
                    end
                end
              reg3241 <= (+(reg3079 > reg3081));
            end
          else
            begin
              for (forvar3223 = (1'h0); (forvar3223 < (2'h2)); forvar3223 = (forvar3223 + (1'h1)))
                begin
                  for (forvar3224 = (1'h0); (forvar3224 < (1'h0)); forvar3224 = (forvar3224 + (1'h1)))
                    begin
                      reg3225 <= (~^$unsigned(($signed(wire3058) || $unsigned((8'ha3)))));
                      reg3226 <= (~|reg3108[(3'h4):(1'h0)]);
                      reg3227 <= (|reg3187[(3'h4):(3'h4)]);
                    end
                  for (forvar3228 = (1'h0); (forvar3228 < (1'h0)); forvar3228 = (forvar3228 + (1'h1)))
                    begin
                      reg3229 <= $signed(((+reg3207[(2'h3):(1'h1)]) ?
                          (~|(forvar3188 & (8'hac))) : reg3105));
                      reg3230 <= reg3148;
                    end
                  for (forvar3231 = (1'h0); (forvar3231 < (1'h1)); forvar3231 = (forvar3231 + (1'h1)))
                    begin
                      reg3232 <= ($unsigned(reg3106[(3'h4):(2'h2)]) << (~reg3133[(1'h1):(1'h1)]));
                      reg3233 <= (((reg3161 >>> (reg3069 << (8'ha4))) ?
                              $signed((wire3062 ?
                                  reg3150 : wire3061)) : ((^~(8'hb9)) ?
                                  reg3198 : (forvar3192 ? reg3084 : (8'hac)))) ?
                          $signed(forvar3224[(4'ha):(1'h1)]) : forvar3209[(2'h2):(2'h2)]);
                    end
                  reg3234 <= (+$unsigned($signed($unsigned(reg3219))));
                end
            end
          if ($unsigned(reg3217))
            begin
              reg3242 <= reg3138;
              for (forvar3243 = (1'h0); (forvar3243 < (2'h3)); forvar3243 = (forvar3243 + (1'h1)))
                begin
                  if (reg3229[(4'hb):(1'h1)])
                    begin
                      reg3244 <= ($signed(reg3219[(1'h1):(1'h0)]) ?
                          reg3089[(4'h8):(3'h4)] : reg3142);
                      reg3245 <= {(8'ha0)};
                      reg3246 <= (reg3232 != reg3113);
                    end
                  else
                    begin
                      reg3244 <= reg3196[(4'he):(3'h5)];
                      reg3245 <= (^$unsigned(((~|reg3189) ?
                          (~|reg3101) : $unsigned(reg3221))));
                      reg3246 <= reg3246[(2'h3):(1'h0)];
                    end
                  reg3247 <= (reg3152[(1'h1):(1'h1)] && $unsigned({$signed(reg3069)}));
                  reg3248 <= ($signed(reg3101[(2'h2):(1'h1)]) ?
                      $signed((-(~|reg3113))) : $signed(($unsigned((8'ha2)) ^~ (^reg3120))));
                end
            end
          else
            begin
              for (forvar3242 = (1'h0); (forvar3242 < (1'h1)); forvar3242 = (forvar3242 + (1'h1)))
                begin
                  reg3243 <= {$signed((-((8'hac) ? reg3163 : reg3110)))};
                  reg3244 <= ((&((reg3080 << (8'ha9)) == (|forvar3243))) ^~ $unsigned($unsigned((forvar3222 & reg3099))));
                  if (({(wire3173 ? reg3189[(3'h6):(3'h5)] : (8'hb2))} ?
                      $signed(reg3083) : reg3219))
                    begin
                      reg3245 <= wire3177[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3245 <= $unsigned(forvar3209);
                      reg3246 <= reg3193;
                    end
                  if (reg3144[(2'h3):(2'h2)])
                    begin
                      reg3247 <= ({(8'ha0)} + (reg3137 ?
                          forvar3223[(2'h3):(2'h2)] : $unsigned({reg3138})));
                      reg3248 <= reg3070;
                    end
                  else
                    begin
                      reg3247 <= reg3206;
                      reg3248 <= ({reg3224[(3'h6):(2'h2)]} ?
                          $signed(($unsigned(forvar3243) ?
                              reg3166[(2'h3):(1'h1)] : reg3225[(3'h5):(2'h2)])) : $unsigned(($signed((8'ha9)) | (!reg3201))));
                      reg3249 <= (8'hb4);
                    end
                end
              reg3250 <= $signed((~&$signed(reg3204[(2'h2):(1'h0)])));
            end
          for (forvar3251 = (1'h0); (forvar3251 < (2'h3)); forvar3251 = (forvar3251 + (1'h1)))
            begin
              for (forvar3252 = (1'h0); (forvar3252 < (1'h1)); forvar3252 = (forvar3252 + (1'h1)))
                begin
                  if ((reg3219 ? $signed(reg3189) : (reg3118 != forvar3178)))
                    begin
                      reg3253 <= reg3203[(1'h1):(1'h0)];
                      reg3254 <= reg3181;
                    end
                  else
                    begin
                      reg3253 <= reg3210;
                      reg3254 <= reg3232;
                    end
                end
            end
          if ($unsigned($unsigned(reg3159[(3'h5):(1'h1)])))
            begin
              if ((^~reg3243[(2'h2):(1'h1)]))
                begin
                  for (forvar3255 = (1'h0); (forvar3255 < (2'h3)); forvar3255 = (forvar3255 + (1'h1)))
                    begin
                      reg3256 <= (~^$signed(reg3166));
                      reg3257 <= $signed($signed($unsigned($unsigned((8'had)))));
                      reg3258 <= ((((~|reg3085) ? {reg3155} : {forvar3213}) ?
                          ($signed(reg3078) ?
                              reg3160 : reg3150) : ((reg3129 >>> reg3074) <<< {(8'hb3)})) + ($signed(((8'hb4) ?
                          (8'hb6) : reg3109)) | {((8'had) ?
                              reg3254 : reg3209)}));
                      reg3259 <= $unsigned((reg3199[(1'h0):(1'h0)] >> (!(reg3191 << reg3153))));
                    end
                  for (forvar3260 = (1'h0); (forvar3260 < (1'h0)); forvar3260 = (forvar3260 + (1'h1)))
                    begin
                      reg3261 <= ($unsigned((~^{reg3204})) ?
                          $signed(wire3177[(2'h3):(1'h0)]) : (reg3137 + (~reg3070)));
                    end
                end
              else
                begin
                  for (forvar3255 = (1'h0); (forvar3255 < (1'h1)); forvar3255 = (forvar3255 + (1'h1)))
                    begin
                      reg3256 <= $unsigned(reg3096);
                    end
                  for (forvar3257 = (1'h0); (forvar3257 < (1'h1)); forvar3257 = (forvar3257 + (1'h1)))
                    begin
                      reg3258 <= $signed(({$signed(reg3235)} ?
                          (~(+forvar3255)) : (~forvar3209[(4'h9):(3'h4)])));
                      reg3259 <= reg3133[(1'h1):(1'h1)];
                      reg3260 <= reg3239[(3'h6):(2'h2)];
                    end
                end
              reg3262 <= (($unsigned((reg3166 ?
                  (8'ha6) : reg3165)) == {$signed(reg3204)}) * ($signed((~&reg3246)) ?
                  $signed(reg3208[(4'hc):(4'ha)]) : $signed(((8'ha9) - reg3259))));
            end
          else
            begin
              reg3255 <= forvar3251;
              if ({(+{(^~reg3207)})})
                begin
                  for (forvar3256 = (1'h0); (forvar3256 < (1'h0)); forvar3256 = (forvar3256 + (1'h1)))
                    begin
                      reg3257 <= (~^(reg3086[(3'h5):(1'h1)] ?
                          reg3071 : forvar3232[(1'h1):(1'h0)]));
                    end
                  for (forvar3258 = (1'h0); (forvar3258 < (1'h0)); forvar3258 = (forvar3258 + (1'h1)))
                    begin
                      reg3259 <= reg3150;
                    end
                end
              else
                begin
                  reg3256 <= ((reg3098 - ($unsigned(reg3125) + $unsigned(reg3215))) ~^ ($unsigned(reg3159[(1'h0):(1'h0)]) | ($unsigned((8'hb5)) >>> ((8'hb1) >= reg3143))));
                  if (((((~reg3081) ?
                          reg3073 : (~|wire3173)) ~^ reg3118[(4'hd):(2'h2)]) ?
                      $unsigned({reg3198}) : $signed(($unsigned(forvar3225) ?
                          ((8'hba) ? reg3182 : reg3249) : (+forvar3257)))))
                    begin
                      reg3257 <= forvar3260[(3'h7):(3'h6)];
                      reg3258 <= (8'ha6);
                      reg3259 <= reg3116;
                    end
                  else
                    begin
                      reg3257 <= $unsigned((8'ha6));
                      reg3258 <= ((|forvar3213[(4'hb):(3'h5)]) ?
                          $signed((-(~forvar3178))) : $unsigned(reg3142));
                      reg3259 <= wire3057[(3'h6):(2'h3)];
                      reg3260 <= $unsigned($unsigned((reg3190 ?
                          (reg3231 ?
                              reg3106 : reg3112) : (reg3160 < reg3201))));
                    end
                  if ((~^$unsigned(reg3154)))
                    begin
                      reg3261 <= {(^(forvar3257[(4'h9):(3'h7)] & $unsigned((8'ha3))))};
                      reg3262 <= reg3112;
                      reg3263 <= $signed(reg3086);
                    end
                  else
                    begin
                      reg3261 <= reg3263[(1'h0):(1'h0)];
                      reg3262 <= reg3166;
                    end
                end
              for (forvar3264 = (1'h0); (forvar3264 < (2'h3)); forvar3264 = (forvar3264 + (1'h1)))
                begin
                  for (forvar3265 = (1'h0); (forvar3265 < (2'h3)); forvar3265 = (forvar3265 + (1'h1)))
                    begin
                      reg3266 <= (forvar3231 ?
                          $unsigned($signed($unsigned((8'ha1)))) : $signed(reg3071[(2'h2):(1'h1)]));
                    end
                end
            end
        end
    end
  assign wire3267 = reg3108;
  assign wire3268 = (reg3133 ?
                        (&reg3203[(1'h1):(1'h0)]) : $unsigned($unsigned((reg3231 && reg3102))));
  assign wire3269 = reg3118[(3'h4):(1'h0)];
  assign wire3270 = $unsigned($signed(((reg3204 < reg3203) - (reg3143 <= reg3226))));
  assign wire3271 = reg3141;
  always
    @(posedge clk) begin
      if (($signed(reg3189) ~^ {reg3245}))
        begin
          reg3272 <= $signed($signed(reg3183));
          reg3273 <= (wire3060[(1'h0):(1'h0)] ? wire3267 : reg3209);
          for (forvar3274 = (1'h0); (forvar3274 < (1'h0)); forvar3274 = (forvar3274 + (1'h1)))
            begin
              for (forvar3275 = (1'h0); (forvar3275 < (2'h3)); forvar3275 = (forvar3275 + (1'h1)))
                begin
                  if ($unsigned(reg3105[(4'ha):(4'h9)]))
                    begin
                      reg3276 <= $unsigned($signed({{reg3107}}));
                      reg3277 <= ($unsigned(($unsigned((8'ha6)) != {reg3212})) >>> wire3267[(2'h3):(1'h0)]);
                      reg3278 <= wire3175;
                      reg3279 <= (~^(reg3259[(2'h3):(2'h3)] <<< reg3150[(2'h3):(2'h2)]));
                    end
                  else
                    begin
                      reg3276 <= $signed(reg3183);
                    end
                  for (forvar3280 = (1'h0); (forvar3280 < (2'h3)); forvar3280 = (forvar3280 + (1'h1)))
                    begin
                      reg3281 <= $unsigned((-$signed(reg3150)));
                      reg3282 <= ({($signed(reg3263) ~^ ((8'ha4) ?
                              reg3123 : reg3279))} + reg3266);
                    end
                  reg3283 <= (~|reg3145);
                  for (forvar3284 = (1'h0); (forvar3284 < (2'h3)); forvar3284 = (forvar3284 + (1'h1)))
                    begin
                      reg3285 <= reg3230[(4'hc):(3'h4)];
                      reg3286 <= (reg3221[(2'h2):(1'h0)] ?
                          {(~|$unsigned(reg3197))} : wire3267);
                    end
                end
            end
        end
      else
        begin
          for (forvar3272 = (1'h0); (forvar3272 < (1'h0)); forvar3272 = (forvar3272 + (1'h1)))
            begin
              for (forvar3273 = (1'h0); (forvar3273 < (1'h1)); forvar3273 = (forvar3273 + (1'h1)))
                begin
                  if ({reg3277[(4'h9):(2'h3)]})
                    begin
                      reg3274 <= {(~&{(reg3160 ? (8'hb2) : wire3060)})};
                      reg3275 <= (((reg3212[(3'h5):(1'h0)] ?
                          $signed(reg3147) : $signed(reg3203)) <= $unsigned($signed(reg3104))) ~^ (-reg3242));
                    end
                  else
                    begin
                      reg3274 <= $unsigned(({$signed((8'hb9))} != reg3208));
                      reg3275 <= reg3117[(4'hb):(2'h3)];
                    end
                end
            end
          if ($unsigned($signed(wire3064)))
            begin
              reg3276 <= (|reg3253);
              for (forvar3277 = (1'h0); (forvar3277 < (2'h3)); forvar3277 = (forvar3277 + (1'h1)))
                begin
                  reg3278 <= reg3237[(4'ha):(1'h1)];
                  if ((~|reg3168))
                    begin
                      reg3279 <= $signed($signed($unsigned((reg3238 ?
                          reg3216 : (8'ha3)))));
                    end
                  else
                    begin
                      reg3279 <= (reg3183[(3'h6):(3'h5)] ?
                          (8'hb2) : (~$unsigned({reg3283})));
                      reg3280 <= (~^reg3283);
                      reg3281 <= (((+(reg3123 >= wire3058)) > ((|reg3263) ?
                              {reg3106} : $signed(reg3212))) ?
                          $unsigned(((reg3231 ? (8'hae) : reg3143) ?
                              (~(8'h9e)) : (wire3060 != wire3060))) : reg3285);
                      reg3282 <= (reg3257[(2'h2):(2'h2)] ?
                          (~^(|$signed(reg3112))) : reg3258[(3'h7):(3'h5)]);
                    end
                end
              if ($unsigned((reg3134[(4'hc):(3'h5)] ?
                  ($unsigned(forvar3272) ?
                      (reg3260 ?
                          reg3183 : reg3248) : reg3195) : ($signed(reg3075) ?
                      (reg3199 ? reg3217 : reg3172) : (reg3076 ?
                          reg3233 : (8'haf))))))
                begin
                  for (forvar3283 = (1'h0); (forvar3283 < (1'h0)); forvar3283 = (forvar3283 + (1'h1)))
                    begin
                      reg3284 <= {reg3244[(2'h3):(1'h0)]};
                    end
                  if ($signed(forvar3280))
                    begin
                      reg3285 <= (|(reg3127 ?
                          {$unsigned((8'ha2))} : $unsigned((~&reg3283))));
                    end
                  else
                    begin
                      reg3285 <= $signed({$unsigned($signed(reg3254))});
                    end
                  for (forvar3286 = (1'h0); (forvar3286 < (2'h2)); forvar3286 = (forvar3286 + (1'h1)))
                    begin
                      reg3287 <= (+reg3159);
                      reg3288 <= $unsigned(reg3198);
                      reg3289 <= $unsigned(reg3207[(4'hd):(4'hd)]);
                      reg3290 <= (&(~((reg3075 ? reg3250 : wire3267) ?
                          (|wire3064) : $signed((8'hb6)))));
                    end
                end
              else
                begin
                  for (forvar3283 = (1'h0); (forvar3283 < (2'h2)); forvar3283 = (forvar3283 + (1'h1)))
                    begin
                      reg3284 <= reg3097;
                      reg3285 <= $unsigned({reg3099});
                    end
                end
            end
          else
            begin
              if (((8'h9f) ?
                  (forvar3277 << (((8'had) ?
                      reg3123 : reg3134) - $signed(reg3257))) : (reg3200[(4'hb):(3'h4)] & wire3060)))
                begin
                  for (forvar3276 = (1'h0); (forvar3276 < (1'h1)); forvar3276 = (forvar3276 + (1'h1)))
                    begin
                      reg3277 <= ((reg3104 ?
                          (-reg3235) : $unsigned((reg3185 > (8'hae)))) <<< $unsigned(reg3200[(2'h2):(2'h2)]));
                      reg3278 <= $signed(wire3057[(3'h6):(3'h5)]);
                      reg3279 <= $unsigned((wire3271 ?
                          reg3083 : (reg3262[(4'ha):(3'h5)] ?
                              $signed(reg3215) : (reg3082 * (8'ha0)))));
                    end
                  for (forvar3280 = (1'h0); (forvar3280 < (1'h1)); forvar3280 = (forvar3280 + (1'h1)))
                    begin
                      reg3281 <= reg3084[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar3276 = (1'h0); (forvar3276 < (2'h3)); forvar3276 = (forvar3276 + (1'h1)))
                    begin
                      reg3277 <= ((-($unsigned(reg3159) == (reg3196 == reg3249))) ?
                          $signed($unsigned(reg3215[(1'h0):(1'h0)])) : $unsigned($unsigned((^reg3083))));
                    end
                  for (forvar3278 = (1'h0); (forvar3278 < (1'h0)); forvar3278 = (forvar3278 + (1'h1)))
                    begin
                      reg3279 <= $unsigned(((reg3110 ?
                              wire3058 : ((8'hba) ? reg3142 : reg3198)) ?
                          $signed(reg3079[(3'h5):(2'h2)]) : $unsigned((reg3100 || (8'ha1)))));
                      reg3280 <= ((wire3176 || $signed(((8'ha6) ?
                              (8'h9d) : reg3212))) ?
                          reg3088[(2'h3):(1'h1)] : $unsigned($unsigned(wire3267)));
                      reg3281 <= $signed($unsigned((~^((8'haa) || reg3254))));
                    end
                  reg3282 <= (~&{(~&reg3198[(1'h1):(1'h1)])});
                  if ((!reg3086))
                    begin
                      reg3283 <= $signed(reg3097[(1'h0):(1'h0)]);
                      reg3284 <= $unsigned($unsigned((~^(^wire3267))));
                      reg3285 <= ((~|(reg3125 ?
                          reg3103[(4'h8):(3'h6)] : {(8'h9e)})) != {forvar3286[(4'h9):(1'h1)]});
                      reg3286 <= $unsigned((reg3283 >> (&$unsigned(reg3275))));
                    end
                  else
                    begin
                      reg3283 <= (~^$signed(reg3114));
                      reg3284 <= (reg3233 != {(&$unsigned(reg3172))});
                      reg3285 <= ((|{$signed(reg3191)}) ?
                          reg3157[(3'h6):(1'h1)] : $unsigned($signed(wire3059)));
                      reg3286 <= $signed((($unsigned(reg3184) ?
                              (reg3073 * reg3246) : (reg3200 > reg3195)) ?
                          {(reg3141 * (8'ha4))} : {$unsigned(reg3190)}));
                    end
                end
            end
          for (forvar3291 = (1'h0); (forvar3291 < (1'h1)); forvar3291 = (forvar3291 + (1'h1)))
            begin
              for (forvar3292 = (1'h0); (forvar3292 < (1'h0)); forvar3292 = (forvar3292 + (1'h1)))
                begin
                  for (forvar3293 = (1'h0); (forvar3293 < (2'h3)); forvar3293 = (forvar3293 + (1'h1)))
                    begin
                      reg3294 <= $unsigned(reg3254);
                    end
                  if (reg3074)
                    begin
                      reg3295 <= (^~(($unsigned(reg3240) >= (-reg3221)) ?
                          reg3266[(3'h6):(3'h4)] : $unsigned((8'hb9))));
                    end
                  else
                    begin
                      reg3295 <= $unsigned($unsigned($unsigned((reg3225 ?
                          reg3098 : reg3133))));
                      reg3296 <= ({reg3207} <= ((~|(reg3217 * (8'haf))) ?
                          (forvar3293 ?
                              reg3245[(1'h1):(1'h0)] : reg3195[(4'he):(4'hd)]) : $signed((reg3254 - reg3274))));
                      reg3297 <= $signed($signed(reg3281[(4'ha):(4'h8)]));
                      reg3298 <= {(~($unsigned(wire3174) || (~reg3208)))};
                    end
                  reg3299 <= reg3285;
                  if ((8'hb7))
                    begin
                      reg3300 <= (^~wire3176[(3'h7):(1'h1)]);
                      reg3301 <= (+(~^$signed(reg3102)));
                    end
                  else
                    begin
                      reg3300 <= (((8'h9c) ?
                              (&(reg3233 < (8'h9c))) : {$signed((8'ha5))}) ?
                          $signed($unsigned((reg3280 ?
                              reg3195 : forvar3275))) : (!$unsigned((+(8'hb5)))));
                      reg3301 <= wire3268;
                      reg3302 <= reg3155[(4'h9):(2'h2)];
                    end
                end
              for (forvar3303 = (1'h0); (forvar3303 < (2'h2)); forvar3303 = (forvar3303 + (1'h1)))
                begin
                  if ($unsigned(reg3200))
                    begin
                      reg3304 <= ($signed(reg3108[(1'h0):(1'h0)]) ?
                          $signed((^(reg3097 ?
                              reg3263 : reg3073))) : (((reg3169 ?
                                  reg3152 : reg3285) >> (~^reg3200)) ?
                              ($unsigned(reg3255) ?
                                  reg3115 : {reg3204}) : $signed((8'hba))));
                      reg3305 <= ($unsigned(reg3169[(4'h8):(3'h6)]) ?
                          $signed(((reg3075 & reg3246) + ((8'hae) ?
                              reg3240 : reg3086))) : (reg3092[(4'hf):(2'h3)] <<< $unsigned(reg3138)));
                      reg3306 <= $unsigned((reg3096 ?
                          $signed($signed(reg3109)) : (~(~&reg3213))));
                      reg3307 <= (($unsigned((reg3098 >= wire3174)) ?
                          (|reg3111) : $unsigned(wire3060[(1'h1):(1'h1)])) == {$unsigned($unsigned(reg3278))});
                    end
                  else
                    begin
                      reg3304 <= $unsigned($unsigned({{(8'hb7)}}));
                    end
                  if ($unsigned((-reg3085)))
                    begin
                      reg3308 <= (($signed($signed(reg3071)) >= reg3083[(3'h5):(1'h0)]) ?
                          (~|reg3170) : $unsigned(reg3154[(3'h6):(2'h2)]));
                      reg3309 <= $signed((~&reg3285));
                    end
                  else
                    begin
                      reg3308 <= reg3089;
                      reg3309 <= $unsigned(reg3285[(3'h5):(2'h3)]);
                      reg3310 <= {$unsigned(((reg3168 ? reg3272 : (8'hb6)) ?
                              (^~reg3266) : reg3106[(3'h7):(3'h6)]))};
                      reg3311 <= (8'hb1);
                    end
                  for (forvar3312 = (1'h0); (forvar3312 < (1'h0)); forvar3312 = (forvar3312 + (1'h1)))
                    begin
                      reg3313 <= reg3181;
                    end
                end
            end
        end
      for (forvar3314 = (1'h0); (forvar3314 < (1'h1)); forvar3314 = (forvar3314 + (1'h1)))
        begin
          if ($signed(reg3259[(2'h3):(1'h0)]))
            begin
              if ((8'ha6))
                begin
                  if (($unsigned(reg3070[(4'h8):(2'h3)]) ?
                      (8'ha3) : (^((^forvar3303) != (~|(8'hb4))))))
                    begin
                      reg3315 <= (((reg3296 ?
                          reg3105[(4'he):(3'h5)] : (reg3094 && reg3281)) && $signed((reg3101 && reg3184))) > reg3289);
                      reg3316 <= $signed(reg3275);
                      reg3317 <= reg3091;
                    end
                  else
                    begin
                      reg3315 <= ((wire3177[(2'h2):(1'h1)] ?
                              ((8'h9c) ?
                                  $unsigned(reg3242) : $unsigned(reg3246)) : {((8'haa) << (8'haf))}) ?
                          (8'hab) : $unsigned(({(8'ha6)} * (reg3134 ?
                              reg3089 : reg3305))));
                      reg3316 <= $signed({reg3280[(4'hb):(4'ha)]});
                      reg3317 <= (!(reg3311 ?
                          (reg3075[(1'h0):(1'h0)] ?
                              $signed(reg3092) : $unsigned((8'ha2))) : ((~^reg3226) < {reg3099})));
                      reg3318 <= reg3258;
                    end
                  if ((&$signed((reg3207[(3'h7):(3'h5)] + (8'hba)))))
                    begin
                      reg3319 <= {reg3313[(1'h1):(1'h0)]};
                      reg3320 <= (((~&(reg3117 ~^ reg3311)) != reg3246) || (-(~{(8'ha7)})));
                      reg3321 <= reg3318;
                      reg3322 <= reg3299;
                    end
                  else
                    begin
                      reg3319 <= reg3196;
                    end
                  for (forvar3323 = (1'h0); (forvar3323 < (2'h3)); forvar3323 = (forvar3323 + (1'h1)))
                    begin
                      reg3324 <= $signed(forvar3280[(2'h3):(1'h1)]);
                      reg3325 <= ($unsigned($unsigned((+wire3177))) ?
                          $signed($unsigned((wire3059 - reg3218))) : reg3218);
                      reg3326 <= $unsigned($unsigned($signed(wire3057[(3'h6):(1'h0)])));
                    end
                  if ($unsigned($signed(((reg3165 + reg3191) ?
                      (wire3064 * reg3320) : $signed(wire3058)))))
                    begin
                      reg3327 <= reg3304;
                      reg3328 <= (8'h9f);
                    end
                  else
                    begin
                      reg3327 <= wire3177;
                      reg3328 <= $signed((&$signed({reg3313})));
                      reg3329 <= reg3213;
                    end
                end
              else
                begin
                  if ($signed(((|$unsigned(wire3270)) ?
                      ($unsigned(reg3089) ?
                          (reg3170 ?
                              (8'ha1) : (8'h9e)) : reg3260) : reg3249[(4'h9):(3'h4)])))
                    begin
                      reg3315 <= forvar3314[(4'ha):(2'h3)];
                    end
                  else
                    begin
                      reg3315 <= $signed(reg3079[(3'h4):(3'h4)]);
                    end
                end
              if ($signed({((reg3212 <<< wire3267) * (~^reg3289))}))
                begin
                  for (forvar3330 = (1'h0); (forvar3330 < (2'h2)); forvar3330 = (forvar3330 + (1'h1)))
                    begin
                      reg3331 <= $signed(forvar3280[(2'h2):(1'h0)]);
                      reg3332 <= (~&reg3084);
                      reg3333 <= {((reg3288[(2'h3):(2'h3)] ?
                              $unsigned(reg3170) : (reg3294 ^~ (8'haa))) - $signed(reg3299[(4'h8):(2'h3)]))};
                    end
                  for (forvar3334 = (1'h0); (forvar3334 < (2'h3)); forvar3334 = (forvar3334 + (1'h1)))
                    begin
                      reg3335 <= $unsigned(wire3059);
                      reg3336 <= reg3144[(3'h7):(1'h0)];
                      reg3337 <= ((+(!$unsigned(reg3092))) ?
                          wire3176 : reg3249);
                      reg3338 <= {$signed({$signed(reg3272)})};
                    end
                end
              else
                begin
                  for (forvar3330 = (1'h0); (forvar3330 < (2'h2)); forvar3330 = (forvar3330 + (1'h1)))
                    begin
                      reg3331 <= (reg3079 || reg3113[(3'h7):(2'h3)]);
                      reg3332 <= {$unsigned(((~|reg3217) << (~^reg3243)))};
                      reg3333 <= (8'haa);
                      reg3334 <= ((reg3181 ?
                              reg3318[(1'h1):(1'h1)] : (forvar3292 && $unsigned(reg3137))) ?
                          reg3118 : ($unsigned((|reg3233)) ?
                              $signed((8'ha9)) : (|(reg3088 ?
                                  reg3187 : reg3115))));
                    end
                end
              reg3339 <= reg3207;
            end
          else
            begin
              if ((^(((^reg3284) ? {reg3083} : (reg3124 - reg3118)) ?
                  $unsigned(reg3281[(4'h9):(2'h2)]) : $signed(reg3336[(3'h5):(1'h0)]))))
                begin
                  if ((~&reg3279[(2'h3):(2'h3)]))
                    begin
                      reg3315 <= reg3166[(4'h8):(3'h7)];
                      reg3316 <= ((reg3086[(2'h2):(2'h2)] - (^~(~^reg3197))) ^ reg3297[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg3315 <= reg3276[(2'h3):(2'h2)];
                      reg3316 <= reg3282[(2'h3):(1'h1)];
                      reg3317 <= {(reg3332 ?
                              (reg3083 ^~ (reg3091 == (8'hb2))) : (&reg3313[(3'h6):(3'h5)]))};
                    end
                  for (forvar3318 = (1'h0); (forvar3318 < (1'h1)); forvar3318 = (forvar3318 + (1'h1)))
                    begin
                      reg3319 <= ((~reg3225[(3'h4):(2'h2)]) != {$signed({(8'ha3)})});
                      reg3320 <= $unsigned(reg3301[(2'h3):(1'h1)]);
                    end
                  for (forvar3321 = (1'h0); (forvar3321 < (1'h1)); forvar3321 = (forvar3321 + (1'h1)))
                    begin
                      reg3322 <= ({$unsigned($unsigned(reg3117))} ?
                          $signed($unsigned({reg3154})) : $signed(reg3087));
                      reg3323 <= $unsigned(reg3111);
                      reg3324 <= (+(!((reg3213 ? reg3112 : reg3302) ?
                          $unsigned(reg3228) : reg3260)));
                    end
                end
              else
                begin
                  reg3315 <= $signed($signed(((reg3263 < reg3153) ?
                      $unsigned(reg3263) : (forvar3272 ^~ (8'hb9)))));
                  if (forvar3277[(3'h6):(2'h3)])
                    begin
                      reg3316 <= reg3274;
                      reg3317 <= reg3295[(4'ha):(3'h6)];
                    end
                  else
                    begin
                      reg3316 <= reg3085[(1'h1):(1'h0)];
                      reg3317 <= ($signed($unsigned($unsigned((8'ha9)))) ?
                          (($unsigned(reg3193) ?
                                  (~|forvar3293) : (reg3306 != reg3254)) ?
                              forvar3293 : $unsigned($unsigned(reg3233))) : (reg3194 ^~ reg3170));
                      reg3318 <= ($signed($signed(reg3231)) ?
                          $unsigned($signed($unsigned((8'hae)))) : $unsigned($signed(reg3324[(3'h7):(3'h4)])));
                      reg3319 <= (~(~^$signed(reg3329[(3'h5):(3'h4)])));
                    end
                end
              reg3325 <= $unsigned((8'ha0));
              for (forvar3326 = (1'h0); (forvar3326 < (1'h1)); forvar3326 = (forvar3326 + (1'h1)))
                begin
                  if ((~|forvar3274[(3'h5):(2'h3)]))
                    begin
                      reg3327 <= reg3212[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg3327 <= forvar3278;
                    end
                end
            end
          if ($signed($unsigned(reg3094[(4'h8):(3'h6)])))
            begin
              if ($signed(forvar3303[(1'h0):(1'h0)]))
                begin
                  for (forvar3340 = (1'h0); (forvar3340 < (1'h1)); forvar3340 = (forvar3340 + (1'h1)))
                    begin
                      reg3341 <= ($signed($unsigned(reg3290)) + (+reg3172));
                      reg3342 <= $unsigned(($signed((!reg3339)) ?
                          ((&reg3322) >= $unsigned(reg3121)) : (forvar3321[(4'ha):(3'h6)] ?
                              $unsigned((8'haf)) : (reg3194 != (8'ha2)))));
                      reg3343 <= reg3111;
                      reg3344 <= reg3084[(2'h2):(1'h1)];
                    end
                end
              else
                begin
                  if (reg3321[(3'h6):(3'h6)])
                    begin
                      reg3340 <= ((reg3248 ?
                              ((-forvar3291) ^~ ((8'hb6) ?
                                  reg3153 : reg3313)) : reg3181[(3'h4):(3'h4)]) ?
                          ((((8'hac) >> reg3332) <<< (reg3342 & reg3090)) ?
                              forvar3291[(2'h2):(2'h2)] : $signed((reg3073 ?
                                  reg3168 : forvar3278))) : (^~$signed($signed(reg3220))));
                      reg3341 <= (reg3198 >= reg3202[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg3340 <= (8'ha2);
                      reg3341 <= reg3278[(4'h8):(4'h8)];
                      reg3342 <= reg3331;
                      reg3343 <= (~&$unsigned(($signed(reg3266) | wire3060)));
                    end
                  for (forvar3344 = (1'h0); (forvar3344 < (1'h1)); forvar3344 = (forvar3344 + (1'h1)))
                    begin
                      reg3345 <= $unsigned(reg3254[(1'h0):(1'h0)]);
                    end
                  if (reg3197[(1'h1):(1'h1)])
                    begin
                      reg3346 <= reg3328[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg3346 <= reg3260;
                    end
                end
            end
          else
            begin
              reg3340 <= reg3199;
            end
        end
      for (forvar3347 = (1'h0); (forvar3347 < (2'h2)); forvar3347 = (forvar3347 + (1'h1)))
        begin
          if (((|($signed(reg3315) >= $signed(reg3294))) ^~ ($signed(reg3297[(3'h6):(3'h6)]) ?
              reg3235[(2'h2):(1'h1)] : reg3182[(3'h6):(1'h0)])))
            begin
              if ($signed(reg3152[(4'hb):(3'h7)]))
                begin
                  reg3348 <= {reg3316};
                  reg3349 <= ($signed($signed($unsigned((8'ha7)))) + ((~$signed((8'hb1))) && {((8'ha3) ?
                          reg3111 : reg3150)}));
                  reg3350 <= $signed(reg3207[(4'hb):(4'h8)]);
                end
              else
                begin
                  for (forvar3348 = (1'h0); (forvar3348 < (1'h1)); forvar3348 = (forvar3348 + (1'h1)))
                    begin
                      reg3349 <= reg3237[(3'h6):(3'h5)];
                      reg3350 <= (-reg3286[(4'h9):(2'h2)]);
                      reg3351 <= (8'hb9);
                    end
                  for (forvar3352 = (1'h0); (forvar3352 < (2'h3)); forvar3352 = (forvar3352 + (1'h1)))
                    begin
                      reg3353 <= ((reg3300[(2'h2):(1'h1)] > $signed((^(8'hb3)))) ?
                          ($unsigned((reg3296 ?
                              reg3204 : wire3063)) == ((reg3345 && reg3263) == $unsigned(reg3193))) : {wire3063});
                      reg3354 <= $unsigned(reg3217[(1'h0):(1'h0)]);
                      reg3355 <= reg3235;
                      reg3356 <= $unsigned($unsigned((|reg3308)));
                    end
                end
              for (forvar3357 = (1'h0); (forvar3357 < (2'h2)); forvar3357 = (forvar3357 + (1'h1)))
                begin
                  for (forvar3358 = (1'h0); (forvar3358 < (1'h0)); forvar3358 = (forvar3358 + (1'h1)))
                    begin
                      reg3359 <= $unsigned(reg3228[(1'h1):(1'h0)]);
                    end
                end
            end
          else
            begin
              for (forvar3348 = (1'h0); (forvar3348 < (1'h1)); forvar3348 = (forvar3348 + (1'h1)))
                begin
                  if (reg3243)
                    begin
                      reg3349 <= reg3127;
                      reg3350 <= reg3100;
                      reg3351 <= reg3235[(1'h1):(1'h0)];
                      reg3352 <= $signed($signed((~&reg3245)));
                    end
                  else
                    begin
                      reg3349 <= (8'hab);
                    end
                end
            end
          for (forvar3360 = (1'h0); (forvar3360 < (1'h0)); forvar3360 = (forvar3360 + (1'h1)))
            begin
              for (forvar3361 = (1'h0); (forvar3361 < (1'h0)); forvar3361 = (forvar3361 + (1'h1)))
                begin
                  reg3362 <= reg3114[(2'h3):(2'h2)];
                end
              for (forvar3363 = (1'h0); (forvar3363 < (2'h2)); forvar3363 = (forvar3363 + (1'h1)))
                begin
                  if (reg3229[(4'ha):(3'h6)])
                    begin
                      reg3364 <= $signed($unsigned($signed($signed(forvar3334))));
                      reg3365 <= (reg3318[(3'h5):(1'h0)] || reg3227);
                      reg3366 <= (reg3260 ?
                          (~{(reg3186 ? reg3148 : reg3184)}) : (reg3364 ?
                              $unsigned($unsigned(reg3169)) : (&reg3161)));
                    end
                  else
                    begin
                      reg3364 <= $signed(($signed(((8'ha2) < reg3170)) != {$unsigned(reg3349)}));
                      reg3365 <= reg3253;
                      reg3366 <= reg3070;
                    end
                  for (forvar3367 = (1'h0); (forvar3367 < (1'h0)); forvar3367 = (forvar3367 + (1'h1)))
                    begin
                      reg3368 <= forvar3361[(4'hd):(2'h3)];
                      reg3369 <= (|{((reg3155 ?
                              reg3153 : forvar3273) - ((8'ha3) >= reg3153))});
                      reg3370 <= $signed($unsigned($unsigned(reg3237[(3'h6):(1'h0)])));
                      reg3371 <= ($unsigned(forvar3363) ?
                          ($unsigned($signed(reg3310)) ?
                              (~&reg3090[(1'h1):(1'h0)]) : reg3368[(3'h7):(2'h2)]) : reg3099);
                    end
                  if (reg3203)
                    begin
                      reg3372 <= $signed(((-$signed(forvar3284)) ?
                          (!$signed(reg3289)) : reg3114[(1'h1):(1'h0)]));
                      reg3373 <= (($signed($signed(forvar3321)) ?
                          ((reg3097 ? reg3195 : reg3199) ?
                              {(8'ha5)} : forvar3283) : ($signed(reg3229) ?
                              (reg3154 ?
                                  wire3062 : reg3201) : (-reg3096))) >= (!$signed($unsigned(reg3234))));
                    end
                  else
                    begin
                      reg3372 <= ((8'haf) >= {(~|$unsigned((8'hb6)))});
                      reg3373 <= $unsigned(reg3311);
                      reg3374 <= reg3350[(1'h1):(1'h1)];
                    end
                end
              reg3375 <= ((+reg3127) ? reg3348 : reg3345[(3'h5):(1'h0)]);
              if (($signed({{(8'ha3)}}) ?
                  $signed({((8'ha4) ?
                          reg3110 : reg3078)}) : reg3262[(4'ha):(1'h0)]))
                begin
                  for (forvar3376 = (1'h0); (forvar3376 < (2'h3)); forvar3376 = (forvar3376 + (1'h1)))
                    begin
                      reg3377 <= reg3232;
                      reg3378 <= {(reg3362[(3'h5):(3'h4)] ?
                              (~^(-forvar3357)) : (((8'hae) ?
                                      (8'hab) : reg3327) ?
                                  reg3280[(4'h9):(1'h0)] : $signed(reg3272)))};
                    end
                end
              else
                begin
                  for (forvar3376 = (1'h0); (forvar3376 < (2'h3)); forvar3376 = (forvar3376 + (1'h1)))
                    begin
                      reg3377 <= (^~(~&$signed((reg3237 ~^ (8'hb1)))));
                      reg3378 <= reg3231[(2'h2):(2'h2)];
                      reg3379 <= $unsigned((!$signed({wire3061})));
                    end
                  for (forvar3380 = (1'h0); (forvar3380 < (1'h0)); forvar3380 = (forvar3380 + (1'h1)))
                    begin
                      reg3381 <= $signed($unsigned($signed((reg3109 >>> reg3204))));
                      reg3382 <= (forvar3360 ?
                          {($signed(forvar3352) ?
                                  (reg3081 ? reg3202 : reg3100) : (reg3297 ?
                                      reg3142 : (8'hb9)))} : (reg3260 ?
                              (reg3224 ^~ {wire3059}) : $signed((!reg3198))));
                      reg3383 <= {((reg3228 << $signed((8'hba))) ?
                              reg3110 : $unsigned($unsigned(reg3220)))};
                    end
                  reg3384 <= reg3070[(3'h6):(3'h6)];
                end
            end
        end
    end
endmodule